module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [28:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [1:0]  io_r_resp_data_0__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [38:0] io_r_resp_data_0_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [2:0]  io_r_resp_data_0_brIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [28:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [1:0]  io_w_req_bits_data__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [38:0] io_w_req_bits_data_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [2:0]  io_w_req_bits_data_brIdx // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_0_R0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_R0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_W0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_W0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_0_clock;
  wire  line_0_reset;
  wire  line_0_valid;
  reg  line_0_valid_reg;
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  line_1_clock;
  wire  line_1_reset;
  wire  line_1_valid;
  reg  line_1_valid_reg;
  wire  _GEN_8 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire  realRen = io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
  wire [73:0] _wdataword_T = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,
    io_w_req_bits_data_brIdx,1'h1}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  wire  line_2_clock;
  wire  line_2_reset;
  wire  line_2_valid;
  reg  line_2_valid_reg;
  wire  line_3_clock;
  wire  line_3_reset;
  wire  line_3_valid;
  reg  line_3_valid_reg;
  reg  rdata_REG; // @[src/main/scala/utils/Hold.scala 28:106]
  reg [73:0] rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_4_clock;
  wire  line_4_reset;
  wire  line_4_valid;
  reg  line_4_valid_reg;
  wire [73:0] _GEN_20 = rdata_REG ? array_0_R0_data : rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  array_0 array_0 ( // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    .R0_addr(array_0_R0_addr),
    .R0_en(array_0_R0_en),
    .R0_clk(array_0_R0_clk),
    .R0_data(array_0_R0_data),
    .W0_addr(array_0_W0_addr),
    .W0_en(array_0_W0_en),
    .W0_clk(array_0_W0_clk),
    .W0_data(array_0_W0_data)
  );
  GEN_w1_line #(.COVER_INDEX(0)) line_0 (
    .clock(line_0_clock),
    .reset(line_0_reset),
    .valid(line_0_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1)) line_1 (
    .clock(line_1_clock),
    .reset(line_1_reset),
    .valid(line_1_valid)
  );
  GEN_w1_line #(.COVER_INDEX(2)) line_2 (
    .clock(line_2_clock),
    .reset(line_2_reset),
    .valid(line_2_valid)
  );
  GEN_w1_line #(.COVER_INDEX(3)) line_3 (
    .clock(line_3_clock),
    .reset(line_3_reset),
    .valid(line_3_valid)
  );
  GEN_w1_line #(.COVER_INDEX(4)) line_4 (
    .clock(line_4_clock),
    .reset(line_4_reset),
    .valid(line_4_valid)
  );
  assign line_0_clock = clock;
  assign line_0_reset = reset;
  assign line_0_valid = resetState ^ line_0_valid_reg;
  assign line_1_clock = clock;
  assign line_1_reset = reset;
  assign line_1_valid = resetFinish ^ line_1_valid_reg;
  assign line_2_clock = clock;
  assign line_2_reset = reset;
  assign line_2_valid = wen ^ line_2_valid_reg;
  assign line_3_clock = clock;
  assign line_3_reset = reset;
  assign line_3_valid = realRen ^ line_3_valid_reg;
  assign line_4_clock = clock;
  assign line_4_reset = reset;
  assign line_4_valid = rdata_REG ^ line_4_valid_reg;
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _GEN_20[73:45]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0__type = _GEN_20[44:43]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_target = _GEN_20[42:4]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_brIdx = _GEN_20[3:1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _GEN_20[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign array_0_R0_addr = io_r_req_bits_setIdx; // @[src/main/scala/utils/Hold.scala 28:87]
  assign array_0_R0_en = io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
  assign array_0_R0_clk = clock; // @[src/main/scala/utils/Hold.scala 28:{87,87}]
  assign array_0_W0_addr = resetState ? resetSet : io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 91:19]
  assign array_0_W0_en = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  assign array_0_W0_clk = clock; // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
  assign array_0_W0_data = resetState ? 74'h0 : _wdataword_T; // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
  always @(posedge clock) begin
    resetState <= reset | _GEN_8; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    line_0_valid_reg <= resetState;
    line_1_valid_reg <= resetFinish;
    line_2_valid_reg <= wen;
    line_3_valid_reg <= realRen;
    rdata_REG <= io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= 74'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (rdata_REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= array_0_R0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_4_valid_reg <= rdata_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  line_0_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_2_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_3_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rdata_REG = _RAND_6[0:0];
  _RAND_7 = {3{`RANDOM}};
  rdata_r_0 = _RAND_7[73:0];
  _RAND_8 = {1{`RANDOM}};
  line_4_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (resetState) begin
      cover(1'h1);
    end
    //
    if (resetFinish) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (realRen) begin
      cover(1'h1);
    end
    //
    if (rdata_REG) begin
      cover(1'h1);
    end
  end
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input  [38:0] io_in_pc_bits, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [38:0] io_out_target, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [2:0]  io_brIdx, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_crosslineJump, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushICache,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_reset; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  reg [1:0] pht [0:511]; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire  pht_phtTaken_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [8:0] pht_phtTaken_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [1:0] pht_phtTaken_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire  pht_cnt_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [8:0] pht_cnt_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [1:0] pht_cnt_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [1:0] pht_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire [8:0] pht_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire  pht_MPORT_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  wire  pht_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  reg [38:0] ras [0:15]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_rasTarget_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_rasTarget_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_MPORT_1_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  reg  flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_5_clock;
  wire  line_5_reset;
  wire  line_5_valid;
  reg  line_5_valid_reg;
  wire  _GEN_11 = io_in_pc_valid ? 1'h0 : flush; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_6_clock;
  wire  line_6_reset;
  wire  line_6_valid;
  reg  line_6_valid_reg;
  wire  _GEN_12 = io_flush | _GEN_11; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire  line_7_clock;
  wire  line_7_reset;
  wire  line_7_valid;
  reg  line_7_valid_reg;
  wire [28:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  _btbHit_T_7 = btb_io_r_req_ready & btb_io_r_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:10] & ~flush & btbHit_REG & ~(pcLatch[1] & btbRead_brIdx[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  wire [1:0] _T_9 = io_out_valid ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 332:94]
  wire  line_8_clock;
  wire  line_8_reset;
  wire  line_8_valid;
  reg  line_8_valid_reg;
  reg [3:0] sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [38:0] rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire  line_9_clock;
  wire  line_9_reset;
  wire  line_9_valid;
  reg  line_9_valid_reg;
  wire  _T_19 = ~bpuUpdateReq_pc[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 353:150]
  wire  _btbWrite_brIdx_T_3 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/BPU.scala 367:46]
  wire [1:0] btbWrite_brIdx_hi = {_btbWrite_brIdx_T_3,bpuUpdateReq_pc[1]}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  reg [1:0] cnt; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
  reg  reqLatch_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg [38:0] reqLatch_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg  reqLatch_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  reg [6:0] reqLatch_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 390:25]
  wire  _T_22 = ~reqLatch_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  _T_23 = reqLatch_valid & _T_22; // @[src/main/scala/nutcore/frontend/BPU.scala 391:24]
  wire  line_10_clock;
  wire  line_10_reset;
  wire  line_10_valid;
  reg  line_10_valid_reg;
  wire [1:0] _newCnt_T_1 = cnt + 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 393:33]
  wire [1:0] _newCnt_T_3 = cnt - 2'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 393:44]
  wire  wen = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 394:44]
  wire  line_11_clock;
  wire  line_11_reset;
  wire  line_11_valid;
  reg  line_11_valid_reg;
  wire  line_12_clock;
  wire  line_12_reset;
  wire  line_12_valid;
  reg  line_12_valid_reg;
  wire  _T_27 = bpuUpdateReq_fuOpType == 7'h5c; // @[src/main/scala/nutcore/frontend/BPU.scala 403:24]
  wire  line_13_clock;
  wire  line_13_reset;
  wire  line_13_valid;
  reg  line_13_valid_reg;
  wire [3:0] _T_29 = sp_value + 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 404:26]
  wire [38:0] _T_31 = bpuUpdateReq_pc + 39'h2; // @[src/main/scala/nutcore/frontend/BPU.scala 404:55]
  wire [38:0] _T_33 = bpuUpdateReq_pc + 39'h4; // @[src/main/scala/nutcore/frontend/BPU.scala 404:69]
  wire  line_14_clock;
  wire  line_14_reset;
  wire  line_14_valid;
  reg  line_14_valid_reg;
  wire  _T_35 = bpuUpdateReq_fuOpType == 7'h5e; // @[src/main/scala/nutcore/frontend/BPU.scala 408:29]
  wire  line_15_clock;
  wire  line_15_reset;
  wire  line_15_valid;
  reg  line_15_valid_reg;
  wire  _T_36 = sp_value == 4'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 409:21]
  wire [3:0] _value_T_4 = sp_value - 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 412:53]
  wire [3:0] _value_T_5 = _T_36 ? 4'h0 : _value_T_4; // @[src/main/scala/nutcore/frontend/BPU.scala 412:22]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [3:0] _io_brIdx_T_1 = {1'h1,crosslineJump,_T_9}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:35]
  wire [3:0] _GEN_39 = {{1'd0}, btbRead_brIdx}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  wire [3:0] _io_brIdx_T_2 = _GEN_39 & _io_brIdx_T_1; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  SRAMTemplate btb ( // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  GEN_w1_line #(.COVER_INDEX(5)) line_5 (
    .clock(line_5_clock),
    .reset(line_5_reset),
    .valid(line_5_valid)
  );
  GEN_w1_line #(.COVER_INDEX(6)) line_6 (
    .clock(line_6_clock),
    .reset(line_6_reset),
    .valid(line_6_valid)
  );
  GEN_w1_line #(.COVER_INDEX(7)) line_7 (
    .clock(line_7_clock),
    .reset(line_7_reset),
    .valid(line_7_valid)
  );
  GEN_w1_line #(.COVER_INDEX(8)) line_8 (
    .clock(line_8_clock),
    .reset(line_8_reset),
    .valid(line_8_valid)
  );
  GEN_w1_line #(.COVER_INDEX(9)) line_9 (
    .clock(line_9_clock),
    .reset(line_9_reset),
    .valid(line_9_valid)
  );
  GEN_w1_line #(.COVER_INDEX(10)) line_10 (
    .clock(line_10_clock),
    .reset(line_10_reset),
    .valid(line_10_valid)
  );
  GEN_w1_line #(.COVER_INDEX(11)) line_11 (
    .clock(line_11_clock),
    .reset(line_11_reset),
    .valid(line_11_valid)
  );
  GEN_w1_line #(.COVER_INDEX(12)) line_12 (
    .clock(line_12_clock),
    .reset(line_12_reset),
    .valid(line_12_valid)
  );
  GEN_w1_line #(.COVER_INDEX(13)) line_13 (
    .clock(line_13_clock),
    .reset(line_13_reset),
    .valid(line_13_valid)
  );
  GEN_w1_line #(.COVER_INDEX(14)) line_14 (
    .clock(line_14_clock),
    .reset(line_14_reset),
    .valid(line_14_valid)
  );
  GEN_w1_line #(.COVER_INDEX(15)) line_15 (
    .clock(line_15_clock),
    .reset(line_15_reset),
    .valid(line_15_valid)
  );
  assign pht_phtTaken_MPORT_en = 1'h1;
  assign pht_phtTaken_MPORT_addr = io_in_pc_bits[9:1];
  assign pht_phtTaken_MPORT_data = pht[pht_phtTaken_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  assign pht_cnt_MPORT_en = 1'h1;
  assign pht_cnt_MPORT_addr = bpuUpdateReq_pc[9:1];
  assign pht_cnt_MPORT_data = pht[pht_cnt_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
  assign pht_MPORT_data = reqLatch_actualTaken ? _newCnt_T_1 : _newCnt_T_3;
  assign pht_MPORT_addr = reqLatch_pc[9:1];
  assign pht_MPORT_mask = 1'h1;
  assign pht_MPORT_en = _T_23 & wen;
  assign ras_rasTarget_MPORT_en = 1'h1;
  assign ras_rasTarget_MPORT_addr = sp_value;
  assign ras_rasTarget_MPORT_data = ras[ras_rasTarget_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  assign ras_MPORT_1_data = bpuUpdateReq_isRVC ? _T_31 : _T_33;
  assign ras_MPORT_1_addr = sp_value + 4'h1;
  assign ras_MPORT_1_mask = 1'h1;
  assign ras_MPORT_1_en = bpuUpdateReq_valid & _T_27;
  assign line_5_clock = clock;
  assign line_5_reset = reset;
  assign line_5_valid = io_in_pc_valid ^ line_5_valid_reg;
  assign line_6_clock = clock;
  assign line_6_reset = reset;
  assign line_6_valid = io_flush ^ line_6_valid_reg;
  assign line_7_clock = clock;
  assign line_7_reset = reset;
  assign line_7_valid = io_in_pc_valid ^ line_7_valid_reg;
  assign line_8_clock = clock;
  assign line_8_reset = reset;
  assign line_8_valid = io_in_pc_valid ^ line_8_valid_reg;
  assign line_9_clock = clock;
  assign line_9_reset = reset;
  assign line_9_valid = io_in_pc_valid ^ line_9_valid_reg;
  assign line_10_clock = clock;
  assign line_10_reset = reset;
  assign line_10_valid = _T_23 ^ line_10_valid_reg;
  assign line_11_clock = clock;
  assign line_11_reset = reset;
  assign line_11_valid = wen ^ line_11_valid_reg;
  assign line_12_clock = clock;
  assign line_12_reset = reset;
  assign line_12_valid = bpuUpdateReq_valid ^ line_12_valid_reg;
  assign line_13_clock = clock;
  assign line_13_reset = reset;
  assign line_13_valid = _T_27 ^ line_13_valid_reg;
  assign line_14_clock = clock;
  assign line_14_reset = reset;
  assign line_14_valid = _T_27 ^ line_14_valid_reg;
  assign line_15_clock = clock;
  assign line_15_reset = reset;
  assign line_15_valid = _T_35 ^ line_15_valid_reg;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[src/main/scala/nutcore/frontend/BPU.scala 416:23]
  assign io_out_valid = 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 420:16]
  assign io_brIdx = _io_brIdx_T_2[2:0]; // @[src/main/scala/nutcore/frontend/BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 375:43]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:10]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_brIdx = {btbWrite_brIdx_hi,_T_19}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  always @(posedge clock) begin
    if (pht_MPORT_en & pht_MPORT_mask) begin
      pht[pht_MPORT_addr] <= pht_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 336:16]
    end
    if (ras_MPORT_1_en & ras_MPORT_1_mask) begin
      ras[ras_MPORT_1_addr] <= ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      flush <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_12;
    end
    line_5_valid_reg <= io_in_pc_valid;
    line_6_valid_reg <= io_flush;
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
      pcLatch <= io_in_pc_bits; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    line_7_valid_reg <= io_in_pc_valid;
    if (reset) begin // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
      btbHit_REG <= 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end else begin
      btbHit_REG <= _btbHit_T_7; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    line_8_valid_reg <= io_in_pc_valid;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      sp_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        sp_value <= _T_29; // @[src/main/scala/nutcore/frontend/BPU.scala 406:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[src/main/scala/nutcore/frontend/BPU.scala 408:48]
        sp_value <= _value_T_5; // @[src/main/scala/nutcore/frontend/BPU.scala 412:16]
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      rasTarget <= ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    line_9_valid_reg <= io_in_pc_valid;
    cnt <= pht_cnt_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 389:20]
    reqLatch_valid <= bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_pc <= bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
    line_10_valid_reg <= _T_23;
    line_11_valid_reg <= wen;
    line_12_valid_reg <= bpuUpdateReq_valid;
    line_13_valid_reg <= _T_27;
    line_14_valid_reg <= _T_27;
    line_15_valid_reg <= _T_35;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_5_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_6_valid_reg = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  pcLatch = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  line_7_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  btbHit_REG = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_8_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sp_value = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  rasTarget = _RAND_10[38:0];
  _RAND_11 = {1{`RANDOM}};
  line_9_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cnt = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  reqLatch_valid = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  reqLatch_pc = _RAND_14[38:0];
  _RAND_15 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  line_10_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_11_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_12_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_13_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_14_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_15_valid_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (io_in_pc_valid) begin
      cover(1'h1);
    end
    //
    if (io_flush) begin
      cover(1'h1);
    end
    //
    if (io_in_pc_valid) begin
      cover(1'h1);
    end
    //
    if (io_in_pc_valid) begin
      cover(1'h1);
    end
    //
    if (io_in_pc_valid) begin
      cover(1'h1);
    end
    //
    if (_T_23) begin
      cover(1'h1);
    end
    //
    if (_T_23 & wen) begin
      cover(1'h1);
    end
    //
    if (bpuUpdateReq_valid) begin
      cover(1'h1);
    end
    //
    if (bpuUpdateReq_valid & _T_27) begin
      cover(1'h1);
    end
    //
    if (bpuUpdateReq_valid & ~_T_27) begin
      cover(1'h1);
    end
    //
    if (bpuUpdateReq_valid & ~_T_27 & _T_35) begin
      cover(1'h1);
    end
  end
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [81:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [81:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input         flushICache,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_reset; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_in_pc_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_in_pc_bits; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_out_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [2:0] bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_crosslineJump; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushICache; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushTLB; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  reg [38:0] pc; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
  wire  _pcUpdate_T = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  pcUpdate = io_redirect_valid | _pcUpdate_T; // @[src/main/scala/nutcore/frontend/IFU.scala 324:36]
  wire [38:0] _snpc_T_2 = pc + 39'h2; // @[src/main/scala/nutcore/frontend/IFU.scala 325:28]
  wire [38:0] _snpc_T_4 = pc + 39'h4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:38]
  wire [38:0] snpc = pc[1] ? _snpc_T_2 : _snpc_T_4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:17]
  reg  crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
  wire  _T = pcUpdate | bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 331:17]
  wire  line_16_clock;
  wire  line_16_reset;
  wire  line_16_valid;
  reg  line_16_valid_reg;
  reg [38:0] crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
  wire  line_17_clock;
  wire  line_17_reset;
  wire  line_17_valid;
  reg  line_17_valid_reg;
  wire [38:0] _npc_T_1 = crosslineJumpLatch ? crosslineJumpTarget : snpc; // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  wire  _npcIsSeq_T_2 = crosslineJumpLatch ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/frontend/IFU.scala 342:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _npcIsSeq_T_2; // @[src/main/scala/nutcore/frontend/IFU.scala 342:21]
  wire [2:0] _brIdx_T = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 350:29]
  wire  line_18_clock;
  wire  line_18_reset;
  wire  line_18_valid;
  reg  line_18_valid_reg;
  wire [42:0] x8_hi = {npcIsSeq,_brIdx_T,npc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  wire  _T_3 = io_imem_resp_ready & io_imem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_19_clock;
  wire  line_19_reset;
  wire  line_19_valid;
  reg  line_19_valid_reg;
  wire  _GEN_8 = io_imem_req_valid | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_20_clock;
  wire  line_20_reset;
  wire  line_20_valid;
  reg  line_20_valid_reg;
  wire  _T_4 = |io_flushVec; // @[src/main/scala/nutcore/frontend/IFU.scala 396:37]
  BPU_inorder bp1 ( // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushICache(bp1_MOUFlushICache),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  GEN_w1_line #(.COVER_INDEX(16)) line_16 (
    .clock(line_16_clock),
    .reset(line_16_reset),
    .valid(line_16_valid)
  );
  GEN_w1_line #(.COVER_INDEX(17)) line_17 (
    .clock(line_17_clock),
    .reset(line_17_reset),
    .valid(line_17_valid)
  );
  GEN_w1_line #(.COVER_INDEX(18)) line_18 (
    .clock(line_18_clock),
    .reset(line_18_reset),
    .valid(line_18_valid)
  );
  GEN_w1_line #(.COVER_INDEX(19)) line_19 (
    .clock(line_19_clock),
    .reset(line_19_reset),
    .valid(line_19_valid)
  );
  GEN_w1_line #(.COVER_INDEX(20)) line_20 (
    .clock(line_20_clock),
    .reset(line_20_reset),
    .valid(line_20_valid)
  );
  assign line_16_clock = clock;
  assign line_16_reset = reset;
  assign line_16_valid = _T ^ line_16_valid_reg;
  assign line_17_clock = clock;
  assign line_17_reset = reset;
  assign line_17_valid = bp1_io_crosslineJump ^ line_17_valid_reg;
  assign line_18_clock = clock;
  assign line_18_reset = reset;
  assign line_18_valid = pcUpdate ^ line_18_valid_reg;
  assign line_19_clock = clock;
  assign line_19_reset = reset;
  assign line_19_valid = io_imem_req_valid ^ line_19_valid_reg;
  assign line_20_clock = clock;
  assign line_20_reset = reset;
  assign line_20_valid = _T_3 ^ line_20_valid_reg;
  assign io_imem_req_valid = io_out_ready; // @[src/main/scala/nutcore/frontend/IFU.scala 373:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[src/main/scala/nutcore/frontend/IFU.scala 371:36]
  assign io_imem_req_bits_user = {x8_hi,pc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 375:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 393:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/IFU.scala 385:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[src/main/scala/nutcore/frontend/IFU.scala 387:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[src/main/scala/nutcore/frontend/IFU.scala 388:26]
  assign io_out_bits_exceptionVec_1 = io_iaf; // @[src/main/scala/nutcore/frontend/IFU.scala 392:46]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[src/main/scala/nutcore/frontend/IFU.scala 389:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 368:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  assign bp1_io_flush = io_redirect_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
  assign bp1_bpuUpdateReq_valid = REG_valid;
  assign bp1_bpuUpdateReq_pc = REG_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = REG_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = REG_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_isRVC;
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
      pc <= 39'h80000000; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end else if (pcUpdate) begin // @[src/main/scala/nutcore/frontend/IFU.scala 361:19]
      if (io_redirect_valid) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= snpc;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
      crosslineJumpLatch <= 1'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 331:34]
      if (bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 332:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    line_16_valid_reg <= _T;
    if (bp1_io_crosslineJump) begin // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
      crosslineJumpTarget <= bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    line_17_valid_reg <= bp1_io_crosslineJump;
    line_18_valid_reg <= pcUpdate;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_3) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_8;
    end
    line_19_valid_reg <= io_imem_req_valid;
    line_20_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_16_valid_reg = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  line_17_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_18_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_19_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_20_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T) begin
      cover(1'h1);
    end
    //
    if (bp1_io_crosslineJump) begin
      cover(1'h1);
    end
    //
    if (pcUpdate) begin
      cover(1'h1);
    end
    //
    if (io_imem_req_valid) begin
      cover(1'h1);
    end
    //
    if (_T_3) begin
      cover(1'h1);
    end
  end
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_0, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_2, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_3, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_4, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_5, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_6, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_7, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_8, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_9, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_10, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_11, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_13, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_14, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_15, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_flush // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
  wire  _instr_T = state == 2'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:23]
  wire  _instr_T_1 = state == 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 44:19]
  reg [15:0] specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
  wire [31:0] _instr_T_4 = {instIn[15:0],specialInstR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:73]
  wire  _pcOffset_T = state == 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:28]
  reg [2:0] pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:21]
  wire  _instr_T_9 = 3'h0 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_13 = _instr_T_9 ? instIn[31:0] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_10 = 3'h2 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_14 = _instr_T_10 ? instIn[47:16] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_17 = _instr_T_13 | _instr_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_11 = 3'h4 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_15 = _instr_T_11 ? instIn[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_18 = _instr_T_17 | _instr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_12 = 3'h6 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_16 = _instr_T_12 ? instIn[79:48] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_19 = _instr_T_18 | _instr_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _instr_T_4 : _instr_T_19; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 34:27]
  wire [7:0] hasException_lo = {io_in_bits_exceptionVec_7,io_in_bits_exceptionVec_6,io_in_bits_exceptionVec_5,
    io_in_bits_exceptionVec_4,io_in_bits_exceptionVec_3,io_in_bits_exceptionVec_2,io_in_bits_exceptionVec_1,
    io_in_bits_exceptionVec_0}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire [15:0] _hasException_T = {io_in_bits_exceptionVec_15,io_in_bits_exceptionVec_14,io_in_bits_exceptionVec_13,
    io_in_bits_exceptionVec_12,io_in_bits_exceptionVec_11,io_in_bits_exceptionVec_10,io_in_bits_exceptionVec_9,
    io_in_bits_exceptionVec_8,hasException_lo}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire  hasException = io_in_valid & |_hasException_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:34]
  wire  _rvcFinish_T = pcOffset == 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:28]
  wire  _rvcFinish_T_1 = ~isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:40]
  wire  _rvcFinish_T_5 = pcOffset == 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:72]
  wire  _rvcFinish_T_11 = pcOffset == 3'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:116]
  wire  _rvcFinish_T_16 = pcOffset == 3'h6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:147]
  wire  _rvcNext_T_13 = _rvcFinish_T_11 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:122]
  wire  _rvcNext_T_15 = ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:135]
  wire  rvcNext = _rvcFinish_T & (isRVC & ~io_in_bits_brIdx[0]) | _rvcFinish_T_5 & (isRVC & ~io_in_bits_brIdx[0]) |
    _rvcFinish_T_11 & _rvcFinish_T_1 & ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:102]
  wire  _rvcSpecial_T_2 = _rvcFinish_T_16 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:37]
  wire  rvcSpecial = _rvcFinish_T_16 & _rvcFinish_T_1 & ~io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:47]
  wire  rvcSpecialJump = _rvcSpecial_T_2 & io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 55:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 56:24]
  wire  _flushIFU_T_2 = _pcOffset_T | state == 2'h1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:36]
  wire  flushIFU = (_pcOffset_T | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:87]
  wire  _T_2 = ~reset; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
  wire  line_21_clock;
  wire  line_21_reset;
  wire  line_21_valid;
  reg  line_21_valid_reg;
  wire  _T_3 = ~(~flushIFU); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
  wire  line_22_clock;
  wire  line_22_reset;
  wire  line_22_valid;
  reg  line_22_valid_reg;
  wire  loadNextInstline = _flushIFU_T_2 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 62:115]
  reg [38:0] specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
  reg [38:0] specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
  reg  specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
  wire  hasCrossBoundaryFault = io_in_bits_exceptionVec_1 | io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 70:73]
  wire  rvcForceLoadNext = _rvcNext_T_13 & io_in_bits_pnpc[2:0] == 3'h4 & _rvcNext_T_15; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 72:86]
  wire  _T_4 = ~io_flush; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:8]
  wire  line_23_clock;
  wire  line_23_reset;
  wire  line_23_valid;
  reg  line_23_valid_reg;
  wire  _T_5 = 2'h0 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire  line_24_clock;
  wire  line_24_reset;
  wire  line_24_valid;
  reg  line_24_valid_reg;
  wire  _canGo_T = rvcFinish | rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:28]
  wire  _canIn_T = rvcFinish | rvcForceLoadNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 104:28]
  wire [38:0] _pnpcOut_T_1 = io_in_bits_pc + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:76]
  wire [38:0] _pnpcOut_T_3 = io_in_bits_pc + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:95]
  wire [38:0] _pnpcOut_T_4 = isRVC ? _pnpcOut_T_1 : _pnpcOut_T_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:55]
  wire [38:0] _pnpcOut_T_5 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:23]
  wire  _T_6 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_7 = _T_6 & rvcFinish; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:26]
  wire  line_25_clock;
  wire  line_25_reset;
  wire  line_25_valid;
  reg  line_25_valid_reg;
  wire [1:0] _GEN_22 = _T_6 & rvcFinish ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:{39,46} 41:22]
  wire  _T_9 = _T_6 & rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:26]
  wire  line_26_clock;
  wire  line_26_reset;
  wire  line_26_valid;
  reg  line_26_valid_reg;
  wire [2:0] _pcOffsetR_T = isRVC ? 3'h2 : 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:38]
  wire [2:0] _pcOffsetR_T_2 = pcOffset + _pcOffsetR_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:33]
  wire [1:0] _GEN_23 = _T_6 & rvcNext ? 2'h1 : _GEN_22; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 109:17]
  wire [2:0] _GEN_24 = _T_6 & rvcNext ? _pcOffsetR_T_2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 110:21 42:26]
  wire  _T_10 = rvcSpecial & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:25]
  wire  line_27_clock;
  wire  line_27_reset;
  wire  line_27_valid;
  reg  line_27_valid_reg;
  wire [1:0] _GEN_25 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_23; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 113:17]
  wire  _T_12 = 2'h1 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire [38:0] _pcOut_T_2 = {io_in_bits_pc[38:3],pcOffsetR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 129:21]
  wire  _T_19 = 2'h2 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire  _T_21 = 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire [38:0] _GEN_49 = 2'h3 == state ? specialPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 164:15 64:23]
  wire [38:0] _GEN_54 = 2'h2 == state ? specialPCR : _GEN_49; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 152:15]
  wire [38:0] _GEN_62 = 2'h1 == state ? _pcOut_T_2 : _GEN_54; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 129:15]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_62; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  wire [38:0] _GEN_26 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 114:22 66:23]
  wire [15:0] _GEN_27 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 115:24 68:25]
  wire  _GEN_28 = rvcSpecial & io_in_valid ? hasCrossBoundaryFault : specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 116:23 69:28]
  wire  _T_11 = rvcSpecialJump & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:29]
  wire  line_28_clock;
  wire  line_28_reset;
  wire  line_28_valid;
  reg  line_28_valid_reg;
  wire [1:0] _GEN_29 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_25; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 119:17]
  wire [38:0] _GEN_30 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_26; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 120:22]
  wire [38:0] _GEN_31 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 121:23 67:24]
  wire [15:0] _GEN_32 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_27; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 122:24]
  wire  _GEN_33 = rvcSpecialJump & io_in_valid ? hasCrossBoundaryFault : _GEN_28; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 123:23]
  wire  line_29_clock;
  wire  line_29_reset;
  wire  line_29_valid;
  reg  line_29_valid_reg;
  wire  line_30_clock;
  wire  line_30_reset;
  wire  line_30_valid;
  reg  line_30_valid_reg;
  wire [38:0] _pnpcOut_T_7 = pcOut + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:68]
  wire [38:0] _pnpcOut_T_9 = pcOut + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:79]
  wire [38:0] _pnpcOut_T_10 = isRVC ? _pnpcOut_T_7 : _pnpcOut_T_9; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:55]
  wire [38:0] _pnpcOut_T_11 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_10; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:23]
  wire  line_31_clock;
  wire  line_31_reset;
  wire  line_31_valid;
  reg  line_31_valid_reg;
  wire  line_32_clock;
  wire  line_32_reset;
  wire  line_32_valid;
  reg  line_32_valid_reg;
  wire  line_33_clock;
  wire  line_33_reset;
  wire  line_33_valid;
  reg  line_33_valid_reg;
  wire  line_34_clock;
  wire  line_34_reset;
  wire  line_34_valid;
  reg  line_34_valid_reg;
  wire  line_35_clock;
  wire  line_35_reset;
  wire  line_35_valid;
  reg  line_35_valid_reg;
  wire  line_36_clock;
  wire  line_36_reset;
  wire  line_36_valid;
  reg  line_36_valid_reg;
  wire [38:0] _pnpcOut_T_13 = specialPCR + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 153:31]
  wire  line_37_clock;
  wire  line_37_reset;
  wire  line_37_valid;
  reg  line_37_valid_reg;
  wire [1:0] _GEN_46 = _T_6 ? 2'h1 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 158:17 41:22]
  wire [2:0] _GEN_47 = _T_6 ? 3'h2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 159:21 42:26]
  wire  line_38_clock;
  wire  line_38_reset;
  wire  line_38_valid;
  reg  line_38_valid_reg;
  wire  line_39_clock;
  wire  line_39_reset;
  wire  line_39_valid;
  reg  line_39_valid_reg;
  wire  line_40_clock;
  wire  line_40_reset;
  wire  line_40_valid;
  reg  line_40_valid_reg;
  wire [1:0] _GEN_48 = _T_6 ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 169:26 170:17 41:22]
  wire [38:0] _GEN_50 = 2'h3 == state ? specialNPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 165:17 65:25]
  wire  _GEN_51 = 2'h3 == state & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 167:15 46:23]
  wire [1:0] _GEN_53 = 2'h3 == state ? _GEN_48 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 41:22]
  wire [38:0] _GEN_55 = 2'h2 == state ? _pnpcOut_T_13 : _GEN_50; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 153:17]
  wire  _GEN_56 = 2'h2 == state ? io_in_valid : _GEN_51; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 155:15]
  wire  _GEN_57 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 156:15]
  wire [1:0] _GEN_58 = 2'h2 == state ? _GEN_46 : _GEN_53; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire [2:0] _GEN_59 = 2'h2 == state ? _GEN_47 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 42:26]
  wire  _GEN_60 = 2'h1 == state ? _canGo_T : _GEN_56; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 127:15]
  wire  _GEN_61 = 2'h1 == state ? _canIn_T : _GEN_57; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 128:15]
  wire [38:0] _GEN_63 = 2'h1 == state ? _pnpcOut_T_11 : _GEN_55; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 130:17]
  wire [1:0] _GEN_64 = 2'h1 == state ? _GEN_29 : _GEN_58; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire  _GEN_70 = 2'h0 == state ? rvcFinish | rvcNext : _GEN_60; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 103:15]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_61; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 104:15]
  wire [38:0] pnpcOut = 2'h0 == state ? _pnpcOut_T_5 : _GEN_63; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  wire  line_41_clock;
  wire  line_41_reset;
  wire  line_41_valid;
  reg  line_41_valid_reg;
  wire  line_42_clock;
  wire  line_42_reset;
  wire  line_42_valid;
  reg  line_42_valid_reg;
  wire  canGo = hasException | _GEN_70; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23 184:11]
  wire  _io_out_bits_brIdx_T_10 = pnpcOut == _pnpcOut_T_9 & _rvcFinish_T_1 | pnpcOut == _pnpcOut_T_7 & isRVC ? 1'h0 : 1'h1
    ; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:27]
  wire  _io_out_bits_exceptionVec_12_T_2 = _instr_T_1 | _instr_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:133]
  GEN_w1_line #(.COVER_INDEX(21)) line_21 (
    .clock(line_21_clock),
    .reset(line_21_reset),
    .valid(line_21_valid)
  );
  GEN_w1_line #(.COVER_INDEX(22)) line_22 (
    .clock(line_22_clock),
    .reset(line_22_reset),
    .valid(line_22_valid)
  );
  GEN_w1_line #(.COVER_INDEX(23)) line_23 (
    .clock(line_23_clock),
    .reset(line_23_reset),
    .valid(line_23_valid)
  );
  GEN_w1_line #(.COVER_INDEX(24)) line_24 (
    .clock(line_24_clock),
    .reset(line_24_reset),
    .valid(line_24_valid)
  );
  GEN_w1_line #(.COVER_INDEX(25)) line_25 (
    .clock(line_25_clock),
    .reset(line_25_reset),
    .valid(line_25_valid)
  );
  GEN_w1_line #(.COVER_INDEX(26)) line_26 (
    .clock(line_26_clock),
    .reset(line_26_reset),
    .valid(line_26_valid)
  );
  GEN_w1_line #(.COVER_INDEX(27)) line_27 (
    .clock(line_27_clock),
    .reset(line_27_reset),
    .valid(line_27_valid)
  );
  GEN_w1_line #(.COVER_INDEX(28)) line_28 (
    .clock(line_28_clock),
    .reset(line_28_reset),
    .valid(line_28_valid)
  );
  GEN_w1_line #(.COVER_INDEX(29)) line_29 (
    .clock(line_29_clock),
    .reset(line_29_reset),
    .valid(line_29_valid)
  );
  GEN_w1_line #(.COVER_INDEX(30)) line_30 (
    .clock(line_30_clock),
    .reset(line_30_reset),
    .valid(line_30_valid)
  );
  GEN_w1_line #(.COVER_INDEX(31)) line_31 (
    .clock(line_31_clock),
    .reset(line_31_reset),
    .valid(line_31_valid)
  );
  GEN_w1_line #(.COVER_INDEX(32)) line_32 (
    .clock(line_32_clock),
    .reset(line_32_reset),
    .valid(line_32_valid)
  );
  GEN_w1_line #(.COVER_INDEX(33)) line_33 (
    .clock(line_33_clock),
    .reset(line_33_reset),
    .valid(line_33_valid)
  );
  GEN_w1_line #(.COVER_INDEX(34)) line_34 (
    .clock(line_34_clock),
    .reset(line_34_reset),
    .valid(line_34_valid)
  );
  GEN_w1_line #(.COVER_INDEX(35)) line_35 (
    .clock(line_35_clock),
    .reset(line_35_reset),
    .valid(line_35_valid)
  );
  GEN_w1_line #(.COVER_INDEX(36)) line_36 (
    .clock(line_36_clock),
    .reset(line_36_reset),
    .valid(line_36_valid)
  );
  GEN_w1_line #(.COVER_INDEX(37)) line_37 (
    .clock(line_37_clock),
    .reset(line_37_reset),
    .valid(line_37_valid)
  );
  GEN_w1_line #(.COVER_INDEX(38)) line_38 (
    .clock(line_38_clock),
    .reset(line_38_reset),
    .valid(line_38_valid)
  );
  GEN_w1_line #(.COVER_INDEX(39)) line_39 (
    .clock(line_39_clock),
    .reset(line_39_reset),
    .valid(line_39_valid)
  );
  GEN_w1_line #(.COVER_INDEX(40)) line_40 (
    .clock(line_40_clock),
    .reset(line_40_reset),
    .valid(line_40_valid)
  );
  GEN_w1_line #(.COVER_INDEX(41)) line_41 (
    .clock(line_41_clock),
    .reset(line_41_reset),
    .valid(line_41_valid)
  );
  GEN_w1_line #(.COVER_INDEX(42)) line_42 (
    .clock(line_42_clock),
    .reset(line_42_reset),
    .valid(line_42_valid)
  );
  assign line_21_clock = clock;
  assign line_21_reset = reset;
  assign line_21_valid = _T_2 ^ line_21_valid_reg;
  assign line_22_clock = clock;
  assign line_22_reset = reset;
  assign line_22_valid = _T_3 ^ line_22_valid_reg;
  assign line_23_clock = clock;
  assign line_23_reset = reset;
  assign line_23_valid = _T_4 ^ line_23_valid_reg;
  assign line_24_clock = clock;
  assign line_24_reset = reset;
  assign line_24_valid = _T_5 ^ line_24_valid_reg;
  assign line_25_clock = clock;
  assign line_25_reset = reset;
  assign line_25_valid = _T_7 ^ line_25_valid_reg;
  assign line_26_clock = clock;
  assign line_26_reset = reset;
  assign line_26_valid = _T_9 ^ line_26_valid_reg;
  assign line_27_clock = clock;
  assign line_27_reset = reset;
  assign line_27_valid = _T_10 ^ line_27_valid_reg;
  assign line_28_clock = clock;
  assign line_28_reset = reset;
  assign line_28_valid = _T_11 ^ line_28_valid_reg;
  assign line_29_clock = clock;
  assign line_29_reset = reset;
  assign line_29_valid = _T_5 ^ line_29_valid_reg;
  assign line_30_clock = clock;
  assign line_30_reset = reset;
  assign line_30_valid = _T_12 ^ line_30_valid_reg;
  assign line_31_clock = clock;
  assign line_31_reset = reset;
  assign line_31_valid = _T_7 ^ line_31_valid_reg;
  assign line_32_clock = clock;
  assign line_32_reset = reset;
  assign line_32_valid = _T_9 ^ line_32_valid_reg;
  assign line_33_clock = clock;
  assign line_33_reset = reset;
  assign line_33_valid = _T_10 ^ line_33_valid_reg;
  assign line_34_clock = clock;
  assign line_34_reset = reset;
  assign line_34_valid = _T_11 ^ line_34_valid_reg;
  assign line_35_clock = clock;
  assign line_35_reset = reset;
  assign line_35_valid = _T_12 ^ line_35_valid_reg;
  assign line_36_clock = clock;
  assign line_36_reset = reset;
  assign line_36_valid = _T_19 ^ line_36_valid_reg;
  assign line_37_clock = clock;
  assign line_37_reset = reset;
  assign line_37_valid = _T_6 ^ line_37_valid_reg;
  assign line_38_clock = clock;
  assign line_38_reset = reset;
  assign line_38_valid = _T_19 ^ line_38_valid_reg;
  assign line_39_clock = clock;
  assign line_39_reset = reset;
  assign line_39_valid = _T_21 ^ line_39_valid_reg;
  assign line_40_clock = clock;
  assign line_40_reset = reset;
  assign line_40_valid = _T_6 ^ line_40_valid_reg;
  assign line_41_clock = clock;
  assign line_41_reset = reset;
  assign line_41_valid = _T_4 ^ line_41_valid_reg;
  assign line_42_clock = clock;
  assign line_42_reset = reset;
  assign line_42_valid = hasException ^ line_42_valid_reg;
  assign io_in_ready = ~io_in_valid | _T_6 & canIn | loadNextInstline; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 196:58]
  assign io_out_valid = io_in_valid & canGo; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 195:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 192:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_62; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  assign io_out_bits_pnpc = 2'h0 == state ? _pnpcOut_T_5 : _GEN_63; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  assign io_out_bits_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 198:28]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_instr_T_1 | _instr_T); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:87]
  assign io_out_bits_brIdx = {{3'd0}, _io_out_bits_brIdx_T_10}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:21]
  assign io_out_bits_crossBoundaryFault = hasCrossBoundaryFault & _io_out_bits_exceptionVec_12_T_2 & ~specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 200:115]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 183:11]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        state <= _GEN_29;
      end else begin
        state <= _GEN_64;
      end
    end else begin
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 175:11]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_32;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_32;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
      pcOffsetR <= 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_24;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_24;
      end else begin
        pcOffsetR <= _GEN_59;
      end
    end
    line_21_valid_reg <= _T_2;
    line_22_valid_reg <= _T_3;
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_30;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_30;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_31;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_31;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
      specialIPFR <= 1'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_33;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_33;
      end
    end
    line_23_valid_reg <= _T_4;
    line_24_valid_reg <= _T_5;
    line_25_valid_reg <= _T_7;
    line_26_valid_reg <= _T_9;
    line_27_valid_reg <= _T_10;
    line_28_valid_reg <= _T_11;
    line_29_valid_reg <= _T_5;
    line_30_valid_reg <= _T_12;
    line_31_valid_reg <= _T_7;
    line_32_valid_reg <= _T_9;
    line_33_valid_reg <= _T_10;
    line_34_valid_reg <= _T_11;
    line_35_valid_reg <= _T_12;
    line_36_valid_reg <= _T_19;
    line_37_valid_reg <= _T_6;
    line_38_valid_reg <= _T_19;
    line_39_valid_reg <= _T_21;
    line_40_valid_reg <= _T_6;
    line_41_valid_reg <= _T_4;
    line_42_valid_reg <= hasException;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~flushIFU)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:61 assert(!flushIFU)\n"); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  line_21_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_22_valid_reg = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  specialPCR = _RAND_5[38:0];
  _RAND_6 = {2{`RANDOM}};
  specialNPCR = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  specialIPFR = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_23_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_24_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_25_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_26_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_27_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_28_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_29_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_30_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_31_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_32_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_33_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_34_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_35_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_36_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_37_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_38_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_39_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_40_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_41_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_42_valid_reg = _RAND_27[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~flushIFU); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_5) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_5 & _T_7) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_5 & _T_9) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_5 & _T_10) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_5 & _T_11) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & _T_12) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & _T_12 & _T_7) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & _T_12 & _T_9) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & _T_12 & _T_10) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & _T_12 & _T_11) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12 & _T_19) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12 & _T_19 & _T_6) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12 & ~_T_19) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12 & ~_T_19 & _T_21) begin
      cover(1'h1);
    end
    //
    if (_T_4 & ~_T_5 & ~_T_12 & ~_T_19 & _T_21 & _T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_4) begin
      cover(1'h1);
    end
    //
    if (hasException) begin
      cover(1'h1);
    end
  end
endmodule
module RVCExpander(
  input         clock,
  input         reset,
  input  [31:0] io_in, // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
  output [31:0] io_out_bits // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 50:20]
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 51:15]
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 33:18]
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 55:23]
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 32:18]
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 54:22]
  wire [27:0] _io_out_s_T_51 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 53:22]
  wire [26:0] _io_out_s_T_73 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f}; // @[src/main/scala/nutcore/frontend/RVC.scala 60:25]
  wire [27:0] _io_out_s_T_93 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 63:23]
  wire [26:0] _io_out_s_T_115 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 62:22]
  wire [27:0] _io_out_s_T_135 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 61:22]
  wire [6:0] _io_out_s_T_144 = io_in[12] ? 7'h7f : 7'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 40:25]
  wire [11:0] _io_out_s_T_146 = {_io_out_s_T_144,io_in[6:2]}; // @[src/main/scala/nutcore/frontend/RVC.scala 40:20]
  wire [31:0] io_out_s_res_8_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 72:24]
  wire  _io_out_s_opc_T_3 = |io_in[11:7]; // @[src/main/scala/nutcore/frontend/RVC.scala 74:24]
  wire [6:0] io_out_s_opc_1 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 74:20]
  wire [31:0] io_out_s_res_9_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],io_out_s_opc_1}; // @[src/main/scala/nutcore/frontend/RVC.scala 75:15]
  wire [31:0] io_out_s_res_10_bits = {_io_out_s_T_144,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 81:22]
  wire  _io_out_s_opc_T_8 = |_io_out_s_T_146; // @[src/main/scala/nutcore/frontend/RVC.scala 87:29]
  wire [6:0] io_out_s_opc_2 = |_io_out_s_T_146 ? 7'h37 : 7'h3f; // @[src/main/scala/nutcore/frontend/RVC.scala 87:20]
  wire [14:0] _io_out_s_me_T_1 = io_in[12] ? 15'h7fff : 15'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 38:24]
  wire [31:0] _io_out_s_me_T_3 = {_io_out_s_me_T_1,io_in[6:2],12'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 38:19]
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_3[31:12],io_in[11:7],io_out_s_opc_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 88:24]
  wire [6:0] io_out_s_opc_3 = _io_out_s_opc_T_8 ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 83:20]
  wire [2:0] _io_out_s_T_183 = io_in[12] ? 3'h7 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 39:29]
  wire [31:0] io_out_s_res_11_bits = {_io_out_s_T_183,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[
    11:7],io_out_s_opc_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 84:15]
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_11_bits : io_out_s_me_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 89:10]
  wire [25:0] _io_out_s_T_205 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 95:21]
  wire [30:0] _GEN_344 = {{5'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [30:0] _io_out_s_T_214 = _GEN_344 | 31'h40000000; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [31:0] _io_out_s_T_223 = {_io_out_s_T_144,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 97:21]
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]}; // @[src/main/scala/nutcore/frontend/RVC.scala 99:77]
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 100:22]
  wire [6:0] io_out_s_opc_4 = io_in[12] ? 7'h3b : 7'h33; // @[src/main/scala/nutcore/frontend/RVC.scala 101:22]
  wire  line_43_clock;
  wire  line_43_reset;
  wire  line_43_valid;
  reg  line_43_valid_reg;
  wire  line_44_clock;
  wire  line_44_reset;
  wire  line_44_valid;
  reg  line_44_valid_reg;
  wire [2:0] _GEN_173 = 3'h1 == _io_out_s_funct_T_2 ? 3'h4 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_45_clock;
  wire  line_45_reset;
  wire  line_45_valid;
  reg  line_45_valid_reg;
  wire [2:0] _GEN_174 = 3'h2 == _io_out_s_funct_T_2 ? 3'h6 : _GEN_173; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_46_clock;
  wire  line_46_reset;
  wire  line_46_valid;
  reg  line_46_valid_reg;
  wire [2:0] _GEN_175 = 3'h3 == _io_out_s_funct_T_2 ? 3'h7 : _GEN_174; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_47_clock;
  wire  line_47_reset;
  wire  line_47_valid;
  reg  line_47_valid_reg;
  wire [2:0] _GEN_176 = 3'h4 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_175; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_48_clock;
  wire  line_48_reset;
  wire  line_48_valid;
  reg  line_48_valid_reg;
  wire [2:0] _GEN_177 = 3'h5 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_176; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_49_clock;
  wire  line_49_reset;
  wire  line_49_valid;
  reg  line_49_valid_reg;
  wire [2:0] _GEN_178 = 3'h6 == _io_out_s_funct_T_2 ? 3'h2 : _GEN_177; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire  line_50_clock;
  wire  line_50_reset;
  wire  line_50_valid;
  reg  line_50_valid_reg;
  wire [2:0] _GEN_179 = 3'h7 == _io_out_s_funct_T_2 ? 3'h3 : _GEN_178; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [24:0] _io_out_s_T_230 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_GEN_179,2'h1,io_in[9:7],io_out_s_opc_4}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:12]
  wire [30:0] _GEN_345 = {{6'd0}, _io_out_s_T_230}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire [30:0] _io_out_s_T_231 = _GEN_345 | io_out_s_sub; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire  line_51_clock;
  wire  line_51_reset;
  wire  line_51_valid;
  reg  line_51_valid_reg;
  wire [31:0] _io_out_s_WIRE_0 = {{6'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire  line_52_clock;
  wire  line_52_reset;
  wire  line_52_valid;
  reg  line_52_valid_reg;
  wire [31:0] _io_out_s_WIRE_1 = {{1'd0}, _io_out_s_T_214}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] _GEN_181 = 2'h1 == io_in[11:10] ? _io_out_s_WIRE_1 : _io_out_s_WIRE_0; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire  line_53_clock;
  wire  line_53_reset;
  wire  line_53_valid;
  reg  line_53_valid_reg;
  wire [31:0] _GEN_182 = 2'h2 == io_in[11:10] ? _io_out_s_T_223 : _GEN_181; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire  line_54_clock;
  wire  line_54_reset;
  wire  line_54_valid;
  reg  line_54_valid_reg;
  wire [31:0] _io_out_s_WIRE_3 = {{1'd0}, _io_out_s_T_231}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] io_out_s_res_12_bits = 2'h3 == io_in[11:10] ? _io_out_s_WIRE_3 : _GEN_182; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [9:0] _io_out_s_T_241 = io_in[12] ? 10'h3ff : 10'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 41:22]
  wire [20:0] _io_out_s_T_249 = {_io_out_s_T_241,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    }; // @[src/main/scala/nutcore/frontend/RVC.scala 41:17]
  wire [31:0] io_out_s_res_13_bits = {_io_out_s_T_249[20],_io_out_s_T_249[10:1],_io_out_s_T_249[11],_io_out_s_T_249[19:
    12],5'h0,7'h6f}; // @[src/main/scala/nutcore/frontend/RVC.scala 91:21]
  wire [4:0] _io_out_s_T_291 = io_in[12] ? 5'h1f : 5'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 42:22]
  wire [12:0] _io_out_s_T_296 = {_io_out_s_T_291,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 42:17]
  wire [31:0] io_out_s_res_14_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h0,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 92:24]
  wire [31:0] io_out_s_res_15_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h1,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 93:24]
  wire [6:0] io_out_s_load_opc = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 110:23]
  wire [25:0] _io_out_s_T_373 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 111:24]
  wire [28:0] _io_out_s_T_383 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 114:25]
  wire [27:0] _io_out_s_T_392 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 113:24]
  wire [28:0] _io_out_s_T_401 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 112:24]
  wire [19:0] _io_out_s_mv_T_2 = {io_in[6:2],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 127:24]
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[src/main/scala/nutcore/frontend/RVC.scala 128:25]
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[src/main/scala/nutcore/frontend/RVC.scala 129:19]
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f}; // @[src/main/scala/nutcore/frontend/RVC.scala 130:25]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[src/main/scala/nutcore/frontend/RVC.scala 131:33]
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2]; // @[src/main/scala/nutcore/frontend/RVC.scala 132:27]
  wire [31:0] io_out_s_mv_bits = {{12'd0}, _io_out_s_mv_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 132:22]
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[src/main/scala/nutcore/frontend/RVC.scala 133:21]
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73}; // @[src/main/scala/nutcore/frontend/RVC.scala 134:23]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000; // @[src/main/scala/nutcore/frontend/RVC.scala 134:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[src/main/scala/nutcore/frontend/RVC.scala 135:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 136:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 137:10]
  wire [8:0] _io_out_s_T_409 = {io_in[9:7],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 37:20]
  wire [28:0] _io_out_s_T_416 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 121:25]
  wire [7:0] _io_out_s_T_422 = {io_in[8:7],io_in[12:9],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 36:20]
  wire [27:0] _io_out_s_T_429 = {_io_out_s_T_422[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_422[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 120:24]
  wire [28:0] _io_out_s_T_442 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 119:24]
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]}; // @[src/main/scala/nutcore/frontend/RVC.scala 148:10]
  wire  line_55_clock;
  wire  line_55_reset;
  wire  line_55_valid;
  reg  line_55_valid_reg;
  wire [31:0] io_out_s_res_bits = {{2'd0}, _io_out_s_T_7}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire  line_56_clock;
  wire  line_56_reset;
  wire  line_56_valid;
  reg  line_56_valid_reg;
  wire [31:0] io_out_s_res_1_bits = {{4'd0}, _io_out_s_T_20}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_185 = 5'h1 == _io_out_T_2 ? io_out_s_res_1_bits : io_out_s_res_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_57_clock;
  wire  line_57_reset;
  wire  line_57_valid;
  reg  line_57_valid_reg;
  wire [31:0] io_out_s_res_2_bits = {{5'd0}, _io_out_s_T_36}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_186 = 5'h2 == _io_out_T_2 ? io_out_s_res_2_bits : _GEN_185; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_58_clock;
  wire  line_58_reset;
  wire  line_58_valid;
  reg  line_58_valid_reg;
  wire [31:0] io_out_s_res_3_bits = {{4'd0}, _io_out_s_T_51}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_187 = 5'h3 == _io_out_T_2 ? io_out_s_res_3_bits : _GEN_186; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_59_clock;
  wire  line_59_reset;
  wire  line_59_valid;
  reg  line_59_valid_reg;
  wire [31:0] io_out_s_res_4_bits = {{5'd0}, _io_out_s_T_73}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_188 = 5'h4 == _io_out_T_2 ? io_out_s_res_4_bits : _GEN_187; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_60_clock;
  wire  line_60_reset;
  wire  line_60_valid;
  reg  line_60_valid_reg;
  wire [31:0] io_out_s_res_5_bits = {{4'd0}, _io_out_s_T_93}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_189 = 5'h5 == _io_out_T_2 ? io_out_s_res_5_bits : _GEN_188; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_61_clock;
  wire  line_61_reset;
  wire  line_61_valid;
  reg  line_61_valid_reg;
  wire [31:0] io_out_s_res_6_bits = {{5'd0}, _io_out_s_T_115}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_190 = 5'h6 == _io_out_T_2 ? io_out_s_res_6_bits : _GEN_189; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_62_clock;
  wire  line_62_reset;
  wire  line_62_valid;
  reg  line_62_valid_reg;
  wire [31:0] io_out_s_res_7_bits = {{4'd0}, _io_out_s_T_135}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_191 = 5'h7 == _io_out_T_2 ? io_out_s_res_7_bits : _GEN_190; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_63_clock;
  wire  line_63_reset;
  wire  line_63_valid;
  reg  line_63_valid_reg;
  wire [31:0] _GEN_192 = 5'h8 == _io_out_T_2 ? io_out_s_res_8_bits : _GEN_191; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_64_clock;
  wire  line_64_reset;
  wire  line_64_valid;
  reg  line_64_valid_reg;
  wire [31:0] _GEN_193 = 5'h9 == _io_out_T_2 ? io_out_s_res_9_bits : _GEN_192; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_65_clock;
  wire  line_65_reset;
  wire  line_65_valid;
  reg  line_65_valid_reg;
  wire [31:0] _GEN_194 = 5'ha == _io_out_T_2 ? io_out_s_res_10_bits : _GEN_193; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_66_clock;
  wire  line_66_reset;
  wire  line_66_valid;
  reg  line_66_valid_reg;
  wire [31:0] _GEN_195 = 5'hb == _io_out_T_2 ? io_out_s_11_bits : _GEN_194; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_67_clock;
  wire  line_67_reset;
  wire  line_67_valid;
  reg  line_67_valid_reg;
  wire [31:0] _GEN_196 = 5'hc == _io_out_T_2 ? io_out_s_res_12_bits : _GEN_195; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_68_clock;
  wire  line_68_reset;
  wire  line_68_valid;
  reg  line_68_valid_reg;
  wire [31:0] _GEN_197 = 5'hd == _io_out_T_2 ? io_out_s_res_13_bits : _GEN_196; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_69_clock;
  wire  line_69_reset;
  wire  line_69_valid;
  reg  line_69_valid_reg;
  wire [31:0] _GEN_198 = 5'he == _io_out_T_2 ? io_out_s_res_14_bits : _GEN_197; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_70_clock;
  wire  line_70_reset;
  wire  line_70_valid;
  reg  line_70_valid_reg;
  wire [31:0] _GEN_199 = 5'hf == _io_out_T_2 ? io_out_s_res_15_bits : _GEN_198; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_71_clock;
  wire  line_71_reset;
  wire  line_71_valid;
  reg  line_71_valid_reg;
  wire [31:0] io_out_s_res_16_bits = {{6'd0}, _io_out_s_T_373}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_200 = 5'h10 == _io_out_T_2 ? io_out_s_res_16_bits : _GEN_199; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_72_clock;
  wire  line_72_reset;
  wire  line_72_valid;
  reg  line_72_valid_reg;
  wire [31:0] io_out_s_res_17_bits = {{3'd0}, _io_out_s_T_383}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_201 = 5'h11 == _io_out_T_2 ? io_out_s_res_17_bits : _GEN_200; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_73_clock;
  wire  line_73_reset;
  wire  line_73_valid;
  reg  line_73_valid_reg;
  wire [31:0] io_out_s_res_18_bits = {{4'd0}, _io_out_s_T_392}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_202 = 5'h12 == _io_out_T_2 ? io_out_s_res_18_bits : _GEN_201; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_74_clock;
  wire  line_74_reset;
  wire  line_74_valid;
  reg  line_74_valid_reg;
  wire [31:0] io_out_s_res_19_bits = {{3'd0}, _io_out_s_T_401}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_203 = 5'h13 == _io_out_T_2 ? io_out_s_res_19_bits : _GEN_202; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_75_clock;
  wire  line_75_reset;
  wire  line_75_valid;
  reg  line_75_valid_reg;
  wire [31:0] _GEN_204 = 5'h14 == _io_out_T_2 ? io_out_s_20_bits : _GEN_203; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_76_clock;
  wire  line_76_reset;
  wire  line_76_valid;
  reg  line_76_valid_reg;
  wire [31:0] io_out_s_res_20_bits = {{3'd0}, _io_out_s_T_416}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_205 = 5'h15 == _io_out_T_2 ? io_out_s_res_20_bits : _GEN_204; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_77_clock;
  wire  line_77_reset;
  wire  line_77_valid;
  reg  line_77_valid_reg;
  wire [31:0] io_out_s_res_21_bits = {{4'd0}, _io_out_s_T_429}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_206 = 5'h16 == _io_out_T_2 ? io_out_s_res_21_bits : _GEN_205; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_78_clock;
  wire  line_78_reset;
  wire  line_78_valid;
  reg  line_78_valid_reg;
  wire [31:0] io_out_s_res_22_bits = {{3'd0}, _io_out_s_T_442}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_207 = 5'h17 == _io_out_T_2 ? io_out_s_res_22_bits : _GEN_206; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_79_clock;
  wire  line_79_reset;
  wire  line_79_valid;
  reg  line_79_valid_reg;
  wire [31:0] _GEN_208 = 5'h18 == _io_out_T_2 ? io_in : _GEN_207; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_80_clock;
  wire  line_80_reset;
  wire  line_80_valid;
  reg  line_80_valid_reg;
  wire [31:0] _GEN_209 = 5'h19 == _io_out_T_2 ? io_in : _GEN_208; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_81_clock;
  wire  line_81_reset;
  wire  line_81_valid;
  reg  line_81_valid_reg;
  wire [31:0] _GEN_210 = 5'h1a == _io_out_T_2 ? io_in : _GEN_209; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_82_clock;
  wire  line_82_reset;
  wire  line_82_valid;
  reg  line_82_valid_reg;
  wire [31:0] _GEN_211 = 5'h1b == _io_out_T_2 ? io_in : _GEN_210; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_83_clock;
  wire  line_83_reset;
  wire  line_83_valid;
  reg  line_83_valid_reg;
  wire [31:0] _GEN_212 = 5'h1c == _io_out_T_2 ? io_in : _GEN_211; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_84_clock;
  wire  line_84_reset;
  wire  line_84_valid;
  reg  line_84_valid_reg;
  wire [31:0] _GEN_213 = 5'h1d == _io_out_T_2 ? io_in : _GEN_212; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_85_clock;
  wire  line_85_reset;
  wire  line_85_valid;
  reg  line_85_valid_reg;
  wire [31:0] _GEN_214 = 5'h1e == _io_out_T_2 ? io_in : _GEN_213; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire  line_86_clock;
  wire  line_86_reset;
  wire  line_86_valid;
  reg  line_86_valid_reg;
  wire  line_87_clock;
  wire  line_87_reset;
  wire  line_87_valid;
  reg  line_87_valid_reg;
  wire  line_88_clock;
  wire  line_88_reset;
  wire  line_88_valid;
  reg  line_88_valid_reg;
  wire  line_89_clock;
  wire  line_89_reset;
  wire  line_89_valid;
  reg  line_89_valid_reg;
  wire  line_90_clock;
  wire  line_90_reset;
  wire  line_90_valid;
  reg  line_90_valid_reg;
  wire  line_91_clock;
  wire  line_91_reset;
  wire  line_91_valid;
  reg  line_91_valid_reg;
  wire  line_92_clock;
  wire  line_92_reset;
  wire  line_92_valid;
  reg  line_92_valid_reg;
  wire  line_93_clock;
  wire  line_93_reset;
  wire  line_93_valid;
  reg  line_93_valid_reg;
  wire  line_94_clock;
  wire  line_94_reset;
  wire  line_94_valid;
  reg  line_94_valid_reg;
  wire  line_95_clock;
  wire  line_95_reset;
  wire  line_95_valid;
  reg  line_95_valid_reg;
  wire  line_96_clock;
  wire  line_96_reset;
  wire  line_96_valid;
  reg  line_96_valid_reg;
  wire  line_97_clock;
  wire  line_97_reset;
  wire  line_97_valid;
  reg  line_97_valid_reg;
  wire  line_98_clock;
  wire  line_98_reset;
  wire  line_98_valid;
  reg  line_98_valid_reg;
  wire  line_99_clock;
  wire  line_99_reset;
  wire  line_99_valid;
  reg  line_99_valid_reg;
  wire  line_100_clock;
  wire  line_100_reset;
  wire  line_100_valid;
  reg  line_100_valid_reg;
  wire  line_101_clock;
  wire  line_101_reset;
  wire  line_101_valid;
  reg  line_101_valid_reg;
  wire  line_102_clock;
  wire  line_102_reset;
  wire  line_102_valid;
  reg  line_102_valid_reg;
  wire  line_103_clock;
  wire  line_103_reset;
  wire  line_103_valid;
  reg  line_103_valid_reg;
  wire  line_104_clock;
  wire  line_104_reset;
  wire  line_104_valid;
  reg  line_104_valid_reg;
  wire  line_105_clock;
  wire  line_105_reset;
  wire  line_105_valid;
  reg  line_105_valid_reg;
  wire  line_106_clock;
  wire  line_106_reset;
  wire  line_106_valid;
  reg  line_106_valid_reg;
  wire  line_107_clock;
  wire  line_107_reset;
  wire  line_107_valid;
  reg  line_107_valid_reg;
  wire  line_108_clock;
  wire  line_108_reset;
  wire  line_108_valid;
  reg  line_108_valid_reg;
  wire  line_109_clock;
  wire  line_109_reset;
  wire  line_109_valid;
  reg  line_109_valid_reg;
  wire  line_110_clock;
  wire  line_110_reset;
  wire  line_110_valid;
  reg  line_110_valid_reg;
  wire  line_111_clock;
  wire  line_111_reset;
  wire  line_111_valid;
  reg  line_111_valid_reg;
  wire  line_112_clock;
  wire  line_112_reset;
  wire  line_112_valid;
  reg  line_112_valid_reg;
  wire  line_113_clock;
  wire  line_113_reset;
  wire  line_113_valid;
  reg  line_113_valid_reg;
  wire  line_114_clock;
  wire  line_114_reset;
  wire  line_114_valid;
  reg  line_114_valid_reg;
  wire  line_115_clock;
  wire  line_115_reset;
  wire  line_115_valid;
  reg  line_115_valid_reg;
  wire  line_116_clock;
  wire  line_116_reset;
  wire  line_116_valid;
  reg  line_116_valid_reg;
  wire  line_117_clock;
  wire  line_117_reset;
  wire  line_117_valid;
  reg  line_117_valid_reg;
  wire  line_118_clock;
  wire  line_118_reset;
  wire  line_118_valid;
  reg  line_118_valid_reg;
  wire  line_119_clock;
  wire  line_119_reset;
  wire  line_119_valid;
  reg  line_119_valid_reg;
  wire  line_120_clock;
  wire  line_120_reset;
  wire  line_120_valid;
  reg  line_120_valid_reg;
  wire  line_121_clock;
  wire  line_121_reset;
  wire  line_121_valid;
  reg  line_121_valid_reg;
  wire  line_122_clock;
  wire  line_122_reset;
  wire  line_122_valid;
  reg  line_122_valid_reg;
  wire  line_123_clock;
  wire  line_123_reset;
  wire  line_123_valid;
  reg  line_123_valid_reg;
  wire  line_124_clock;
  wire  line_124_reset;
  wire  line_124_valid;
  reg  line_124_valid_reg;
  wire  line_125_clock;
  wire  line_125_reset;
  wire  line_125_valid;
  reg  line_125_valid_reg;
  wire  line_126_clock;
  wire  line_126_reset;
  wire  line_126_valid;
  reg  line_126_valid_reg;
  wire  line_127_clock;
  wire  line_127_reset;
  wire  line_127_valid;
  reg  line_127_valid_reg;
  wire  line_128_clock;
  wire  line_128_reset;
  wire  line_128_valid;
  reg  line_128_valid_reg;
  wire  line_129_clock;
  wire  line_129_reset;
  wire  line_129_valid;
  reg  line_129_valid_reg;
  wire  line_130_clock;
  wire  line_130_reset;
  wire  line_130_valid;
  reg  line_130_valid_reg;
  wire  line_131_clock;
  wire  line_131_reset;
  wire  line_131_valid;
  reg  line_131_valid_reg;
  wire  line_132_clock;
  wire  line_132_reset;
  wire  line_132_valid;
  reg  line_132_valid_reg;
  wire  line_133_clock;
  wire  line_133_reset;
  wire  line_133_valid;
  reg  line_133_valid_reg;
  wire  line_134_clock;
  wire  line_134_reset;
  wire  line_134_valid;
  reg  line_134_valid_reg;
  wire  line_135_clock;
  wire  line_135_reset;
  wire  line_135_valid;
  reg  line_135_valid_reg;
  wire  line_136_clock;
  wire  line_136_reset;
  wire  line_136_valid;
  reg  line_136_valid_reg;
  wire  line_137_clock;
  wire  line_137_reset;
  wire  line_137_valid;
  reg  line_137_valid_reg;
  wire  line_138_clock;
  wire  line_138_reset;
  wire  line_138_valid;
  reg  line_138_valid_reg;
  wire  line_139_clock;
  wire  line_139_reset;
  wire  line_139_valid;
  reg  line_139_valid_reg;
  wire  line_140_clock;
  wire  line_140_reset;
  wire  line_140_valid;
  reg  line_140_valid_reg;
  wire  line_141_clock;
  wire  line_141_reset;
  wire  line_141_valid;
  reg  line_141_valid_reg;
  wire  line_142_clock;
  wire  line_142_reset;
  wire  line_142_valid;
  reg  line_142_valid_reg;
  wire  line_143_clock;
  wire  line_143_reset;
  wire  line_143_valid;
  reg  line_143_valid_reg;
  wire  line_144_clock;
  wire  line_144_reset;
  wire  line_144_valid;
  reg  line_144_valid_reg;
  wire  line_145_clock;
  wire  line_145_reset;
  wire  line_145_valid;
  reg  line_145_valid_reg;
  wire  line_146_clock;
  wire  line_146_reset;
  wire  line_146_valid;
  reg  line_146_valid_reg;
  wire  line_147_clock;
  wire  line_147_reset;
  wire  line_147_valid;
  reg  line_147_valid_reg;
  wire  line_148_clock;
  wire  line_148_reset;
  wire  line_148_valid;
  reg  line_148_valid_reg;
  wire  line_149_clock;
  wire  line_149_reset;
  wire  line_149_valid;
  reg  line_149_valid_reg;
  wire  line_150_clock;
  wire  line_150_reset;
  wire  line_150_valid;
  reg  line_150_valid_reg;
  wire  line_151_clock;
  wire  line_151_reset;
  wire  line_151_valid;
  reg  line_151_valid_reg;
  wire  line_152_clock;
  wire  line_152_reset;
  wire  line_152_valid;
  reg  line_152_valid_reg;
  wire  line_153_clock;
  wire  line_153_reset;
  wire  line_153_valid;
  reg  line_153_valid_reg;
  wire  line_154_clock;
  wire  line_154_reset;
  wire  line_154_valid;
  reg  line_154_valid_reg;
  wire  line_155_clock;
  wire  line_155_reset;
  wire  line_155_valid;
  reg  line_155_valid_reg;
  wire  line_156_clock;
  wire  line_156_reset;
  wire  line_156_valid;
  reg  line_156_valid_reg;
  wire  line_157_clock;
  wire  line_157_reset;
  wire  line_157_valid;
  reg  line_157_valid_reg;
  wire  line_158_clock;
  wire  line_158_reset;
  wire  line_158_valid;
  reg  line_158_valid_reg;
  wire  line_159_clock;
  wire  line_159_reset;
  wire  line_159_valid;
  reg  line_159_valid_reg;
  wire  line_160_clock;
  wire  line_160_reset;
  wire  line_160_valid;
  reg  line_160_valid_reg;
  wire  line_161_clock;
  wire  line_161_reset;
  wire  line_161_valid;
  reg  line_161_valid_reg;
  wire  line_162_clock;
  wire  line_162_reset;
  wire  line_162_valid;
  reg  line_162_valid_reg;
  wire  line_163_clock;
  wire  line_163_reset;
  wire  line_163_valid;
  reg  line_163_valid_reg;
  wire  line_164_clock;
  wire  line_164_reset;
  wire  line_164_valid;
  reg  line_164_valid_reg;
  wire  line_165_clock;
  wire  line_165_reset;
  wire  line_165_valid;
  reg  line_165_valid_reg;
  wire  line_166_clock;
  wire  line_166_reset;
  wire  line_166_valid;
  reg  line_166_valid_reg;
  wire  line_167_clock;
  wire  line_167_reset;
  wire  line_167_valid;
  reg  line_167_valid_reg;
  wire  line_168_clock;
  wire  line_168_reset;
  wire  line_168_valid;
  reg  line_168_valid_reg;
  wire  line_169_clock;
  wire  line_169_reset;
  wire  line_169_valid;
  reg  line_169_valid_reg;
  wire  line_170_clock;
  wire  line_170_reset;
  wire  line_170_valid;
  reg  line_170_valid_reg;
  wire  line_171_clock;
  wire  line_171_reset;
  wire  line_171_valid;
  reg  line_171_valid_reg;
  wire  line_172_clock;
  wire  line_172_reset;
  wire  line_172_valid;
  reg  line_172_valid_reg;
  wire  line_173_clock;
  wire  line_173_reset;
  wire  line_173_valid;
  reg  line_173_valid_reg;
  wire  line_174_clock;
  wire  line_174_reset;
  wire  line_174_valid;
  reg  line_174_valid_reg;
  wire  line_175_clock;
  wire  line_175_reset;
  wire  line_175_valid;
  reg  line_175_valid_reg;
  wire  line_176_clock;
  wire  line_176_reset;
  wire  line_176_valid;
  reg  line_176_valid_reg;
  wire  line_177_clock;
  wire  line_177_reset;
  wire  line_177_valid;
  reg  line_177_valid_reg;
  wire  line_178_clock;
  wire  line_178_reset;
  wire  line_178_valid;
  reg  line_178_valid_reg;
  wire  line_179_clock;
  wire  line_179_reset;
  wire  line_179_valid;
  reg  line_179_valid_reg;
  wire  line_180_clock;
  wire  line_180_reset;
  wire  line_180_valid;
  reg  line_180_valid_reg;
  wire  line_181_clock;
  wire  line_181_reset;
  wire  line_181_valid;
  reg  line_181_valid_reg;
  wire  line_182_clock;
  wire  line_182_reset;
  wire  line_182_valid;
  reg  line_182_valid_reg;
  wire  line_183_clock;
  wire  line_183_reset;
  wire  line_183_valid;
  reg  line_183_valid_reg;
  wire  line_184_clock;
  wire  line_184_reset;
  wire  line_184_valid;
  reg  line_184_valid_reg;
  wire  line_185_clock;
  wire  line_185_reset;
  wire  line_185_valid;
  reg  line_185_valid_reg;
  wire  line_186_clock;
  wire  line_186_reset;
  wire  line_186_valid;
  reg  line_186_valid_reg;
  wire  line_187_clock;
  wire  line_187_reset;
  wire  line_187_valid;
  reg  line_187_valid_reg;
  wire  line_188_clock;
  wire  line_188_reset;
  wire  line_188_valid;
  reg  line_188_valid_reg;
  wire  line_189_clock;
  wire  line_189_reset;
  wire  line_189_valid;
  reg  line_189_valid_reg;
  wire  line_190_clock;
  wire  line_190_reset;
  wire  line_190_valid;
  reg  line_190_valid_reg;
  wire  line_191_clock;
  wire  line_191_reset;
  wire  line_191_valid;
  reg  line_191_valid_reg;
  wire  line_192_clock;
  wire  line_192_reset;
  wire  line_192_valid;
  reg  line_192_valid_reg;
  wire  line_193_clock;
  wire  line_193_reset;
  wire  line_193_valid;
  reg  line_193_valid_reg;
  wire  line_194_clock;
  wire  line_194_reset;
  wire  line_194_valid;
  reg  line_194_valid_reg;
  wire  line_195_clock;
  wire  line_195_reset;
  wire  line_195_valid;
  reg  line_195_valid_reg;
  wire  line_196_clock;
  wire  line_196_reset;
  wire  line_196_valid;
  reg  line_196_valid_reg;
  wire  line_197_clock;
  wire  line_197_reset;
  wire  line_197_valid;
  reg  line_197_valid_reg;
  wire  line_198_clock;
  wire  line_198_reset;
  wire  line_198_valid;
  reg  line_198_valid_reg;
  wire  line_199_clock;
  wire  line_199_reset;
  wire  line_199_valid;
  reg  line_199_valid_reg;
  wire  line_200_clock;
  wire  line_200_reset;
  wire  line_200_valid;
  reg  line_200_valid_reg;
  wire  line_201_clock;
  wire  line_201_reset;
  wire  line_201_valid;
  reg  line_201_valid_reg;
  wire  line_202_clock;
  wire  line_202_reset;
  wire  line_202_valid;
  reg  line_202_valid_reg;
  wire  line_203_clock;
  wire  line_203_reset;
  wire  line_203_valid;
  reg  line_203_valid_reg;
  wire  line_204_clock;
  wire  line_204_reset;
  wire  line_204_valid;
  reg  line_204_valid_reg;
  wire  line_205_clock;
  wire  line_205_reset;
  wire  line_205_valid;
  reg  line_205_valid_reg;
  wire  line_206_clock;
  wire  line_206_reset;
  wire  line_206_valid;
  reg  line_206_valid_reg;
  wire  line_207_clock;
  wire  line_207_reset;
  wire  line_207_valid;
  reg  line_207_valid_reg;
  wire  line_208_clock;
  wire  line_208_reset;
  wire  line_208_valid;
  reg  line_208_valid_reg;
  wire  line_209_clock;
  wire  line_209_reset;
  wire  line_209_valid;
  reg  line_209_valid_reg;
  wire  line_210_clock;
  wire  line_210_reset;
  wire  line_210_valid;
  reg  line_210_valid_reg;
  wire  line_211_clock;
  wire  line_211_reset;
  wire  line_211_valid;
  reg  line_211_valid_reg;
  wire  line_212_clock;
  wire  line_212_reset;
  wire  line_212_valid;
  reg  line_212_valid_reg;
  wire  line_213_clock;
  wire  line_213_reset;
  wire  line_213_valid;
  reg  line_213_valid_reg;
  wire  line_214_clock;
  wire  line_214_reset;
  wire  line_214_valid;
  reg  line_214_valid_reg;
  GEN_w1_line #(.COVER_INDEX(43)) line_43 (
    .clock(line_43_clock),
    .reset(line_43_reset),
    .valid(line_43_valid)
  );
  GEN_w1_line #(.COVER_INDEX(44)) line_44 (
    .clock(line_44_clock),
    .reset(line_44_reset),
    .valid(line_44_valid)
  );
  GEN_w1_line #(.COVER_INDEX(45)) line_45 (
    .clock(line_45_clock),
    .reset(line_45_reset),
    .valid(line_45_valid)
  );
  GEN_w1_line #(.COVER_INDEX(46)) line_46 (
    .clock(line_46_clock),
    .reset(line_46_reset),
    .valid(line_46_valid)
  );
  GEN_w1_line #(.COVER_INDEX(47)) line_47 (
    .clock(line_47_clock),
    .reset(line_47_reset),
    .valid(line_47_valid)
  );
  GEN_w1_line #(.COVER_INDEX(48)) line_48 (
    .clock(line_48_clock),
    .reset(line_48_reset),
    .valid(line_48_valid)
  );
  GEN_w1_line #(.COVER_INDEX(49)) line_49 (
    .clock(line_49_clock),
    .reset(line_49_reset),
    .valid(line_49_valid)
  );
  GEN_w1_line #(.COVER_INDEX(50)) line_50 (
    .clock(line_50_clock),
    .reset(line_50_reset),
    .valid(line_50_valid)
  );
  GEN_w1_line #(.COVER_INDEX(51)) line_51 (
    .clock(line_51_clock),
    .reset(line_51_reset),
    .valid(line_51_valid)
  );
  GEN_w1_line #(.COVER_INDEX(52)) line_52 (
    .clock(line_52_clock),
    .reset(line_52_reset),
    .valid(line_52_valid)
  );
  GEN_w1_line #(.COVER_INDEX(53)) line_53 (
    .clock(line_53_clock),
    .reset(line_53_reset),
    .valid(line_53_valid)
  );
  GEN_w1_line #(.COVER_INDEX(54)) line_54 (
    .clock(line_54_clock),
    .reset(line_54_reset),
    .valid(line_54_valid)
  );
  GEN_w1_line #(.COVER_INDEX(55)) line_55 (
    .clock(line_55_clock),
    .reset(line_55_reset),
    .valid(line_55_valid)
  );
  GEN_w1_line #(.COVER_INDEX(56)) line_56 (
    .clock(line_56_clock),
    .reset(line_56_reset),
    .valid(line_56_valid)
  );
  GEN_w1_line #(.COVER_INDEX(57)) line_57 (
    .clock(line_57_clock),
    .reset(line_57_reset),
    .valid(line_57_valid)
  );
  GEN_w1_line #(.COVER_INDEX(58)) line_58 (
    .clock(line_58_clock),
    .reset(line_58_reset),
    .valid(line_58_valid)
  );
  GEN_w1_line #(.COVER_INDEX(59)) line_59 (
    .clock(line_59_clock),
    .reset(line_59_reset),
    .valid(line_59_valid)
  );
  GEN_w1_line #(.COVER_INDEX(60)) line_60 (
    .clock(line_60_clock),
    .reset(line_60_reset),
    .valid(line_60_valid)
  );
  GEN_w1_line #(.COVER_INDEX(61)) line_61 (
    .clock(line_61_clock),
    .reset(line_61_reset),
    .valid(line_61_valid)
  );
  GEN_w1_line #(.COVER_INDEX(62)) line_62 (
    .clock(line_62_clock),
    .reset(line_62_reset),
    .valid(line_62_valid)
  );
  GEN_w1_line #(.COVER_INDEX(63)) line_63 (
    .clock(line_63_clock),
    .reset(line_63_reset),
    .valid(line_63_valid)
  );
  GEN_w1_line #(.COVER_INDEX(64)) line_64 (
    .clock(line_64_clock),
    .reset(line_64_reset),
    .valid(line_64_valid)
  );
  GEN_w1_line #(.COVER_INDEX(65)) line_65 (
    .clock(line_65_clock),
    .reset(line_65_reset),
    .valid(line_65_valid)
  );
  GEN_w1_line #(.COVER_INDEX(66)) line_66 (
    .clock(line_66_clock),
    .reset(line_66_reset),
    .valid(line_66_valid)
  );
  GEN_w1_line #(.COVER_INDEX(67)) line_67 (
    .clock(line_67_clock),
    .reset(line_67_reset),
    .valid(line_67_valid)
  );
  GEN_w1_line #(.COVER_INDEX(68)) line_68 (
    .clock(line_68_clock),
    .reset(line_68_reset),
    .valid(line_68_valid)
  );
  GEN_w1_line #(.COVER_INDEX(69)) line_69 (
    .clock(line_69_clock),
    .reset(line_69_reset),
    .valid(line_69_valid)
  );
  GEN_w1_line #(.COVER_INDEX(70)) line_70 (
    .clock(line_70_clock),
    .reset(line_70_reset),
    .valid(line_70_valid)
  );
  GEN_w1_line #(.COVER_INDEX(71)) line_71 (
    .clock(line_71_clock),
    .reset(line_71_reset),
    .valid(line_71_valid)
  );
  GEN_w1_line #(.COVER_INDEX(72)) line_72 (
    .clock(line_72_clock),
    .reset(line_72_reset),
    .valid(line_72_valid)
  );
  GEN_w1_line #(.COVER_INDEX(73)) line_73 (
    .clock(line_73_clock),
    .reset(line_73_reset),
    .valid(line_73_valid)
  );
  GEN_w1_line #(.COVER_INDEX(74)) line_74 (
    .clock(line_74_clock),
    .reset(line_74_reset),
    .valid(line_74_valid)
  );
  GEN_w1_line #(.COVER_INDEX(75)) line_75 (
    .clock(line_75_clock),
    .reset(line_75_reset),
    .valid(line_75_valid)
  );
  GEN_w1_line #(.COVER_INDEX(76)) line_76 (
    .clock(line_76_clock),
    .reset(line_76_reset),
    .valid(line_76_valid)
  );
  GEN_w1_line #(.COVER_INDEX(77)) line_77 (
    .clock(line_77_clock),
    .reset(line_77_reset),
    .valid(line_77_valid)
  );
  GEN_w1_line #(.COVER_INDEX(78)) line_78 (
    .clock(line_78_clock),
    .reset(line_78_reset),
    .valid(line_78_valid)
  );
  GEN_w1_line #(.COVER_INDEX(79)) line_79 (
    .clock(line_79_clock),
    .reset(line_79_reset),
    .valid(line_79_valid)
  );
  GEN_w1_line #(.COVER_INDEX(80)) line_80 (
    .clock(line_80_clock),
    .reset(line_80_reset),
    .valid(line_80_valid)
  );
  GEN_w1_line #(.COVER_INDEX(81)) line_81 (
    .clock(line_81_clock),
    .reset(line_81_reset),
    .valid(line_81_valid)
  );
  GEN_w1_line #(.COVER_INDEX(82)) line_82 (
    .clock(line_82_clock),
    .reset(line_82_reset),
    .valid(line_82_valid)
  );
  GEN_w1_line #(.COVER_INDEX(83)) line_83 (
    .clock(line_83_clock),
    .reset(line_83_reset),
    .valid(line_83_valid)
  );
  GEN_w1_line #(.COVER_INDEX(84)) line_84 (
    .clock(line_84_clock),
    .reset(line_84_reset),
    .valid(line_84_valid)
  );
  GEN_w1_line #(.COVER_INDEX(85)) line_85 (
    .clock(line_85_clock),
    .reset(line_85_reset),
    .valid(line_85_valid)
  );
  GEN_w1_line #(.COVER_INDEX(86)) line_86 (
    .clock(line_86_clock),
    .reset(line_86_reset),
    .valid(line_86_valid)
  );
  GEN_w1_line #(.COVER_INDEX(87)) line_87 (
    .clock(line_87_clock),
    .reset(line_87_reset),
    .valid(line_87_valid)
  );
  GEN_w1_line #(.COVER_INDEX(88)) line_88 (
    .clock(line_88_clock),
    .reset(line_88_reset),
    .valid(line_88_valid)
  );
  GEN_w1_line #(.COVER_INDEX(89)) line_89 (
    .clock(line_89_clock),
    .reset(line_89_reset),
    .valid(line_89_valid)
  );
  GEN_w1_line #(.COVER_INDEX(90)) line_90 (
    .clock(line_90_clock),
    .reset(line_90_reset),
    .valid(line_90_valid)
  );
  GEN_w1_line #(.COVER_INDEX(91)) line_91 (
    .clock(line_91_clock),
    .reset(line_91_reset),
    .valid(line_91_valid)
  );
  GEN_w1_line #(.COVER_INDEX(92)) line_92 (
    .clock(line_92_clock),
    .reset(line_92_reset),
    .valid(line_92_valid)
  );
  GEN_w1_line #(.COVER_INDEX(93)) line_93 (
    .clock(line_93_clock),
    .reset(line_93_reset),
    .valid(line_93_valid)
  );
  GEN_w1_line #(.COVER_INDEX(94)) line_94 (
    .clock(line_94_clock),
    .reset(line_94_reset),
    .valid(line_94_valid)
  );
  GEN_w1_line #(.COVER_INDEX(95)) line_95 (
    .clock(line_95_clock),
    .reset(line_95_reset),
    .valid(line_95_valid)
  );
  GEN_w1_line #(.COVER_INDEX(96)) line_96 (
    .clock(line_96_clock),
    .reset(line_96_reset),
    .valid(line_96_valid)
  );
  GEN_w1_line #(.COVER_INDEX(97)) line_97 (
    .clock(line_97_clock),
    .reset(line_97_reset),
    .valid(line_97_valid)
  );
  GEN_w1_line #(.COVER_INDEX(98)) line_98 (
    .clock(line_98_clock),
    .reset(line_98_reset),
    .valid(line_98_valid)
  );
  GEN_w1_line #(.COVER_INDEX(99)) line_99 (
    .clock(line_99_clock),
    .reset(line_99_reset),
    .valid(line_99_valid)
  );
  GEN_w1_line #(.COVER_INDEX(100)) line_100 (
    .clock(line_100_clock),
    .reset(line_100_reset),
    .valid(line_100_valid)
  );
  GEN_w1_line #(.COVER_INDEX(101)) line_101 (
    .clock(line_101_clock),
    .reset(line_101_reset),
    .valid(line_101_valid)
  );
  GEN_w1_line #(.COVER_INDEX(102)) line_102 (
    .clock(line_102_clock),
    .reset(line_102_reset),
    .valid(line_102_valid)
  );
  GEN_w1_line #(.COVER_INDEX(103)) line_103 (
    .clock(line_103_clock),
    .reset(line_103_reset),
    .valid(line_103_valid)
  );
  GEN_w1_line #(.COVER_INDEX(104)) line_104 (
    .clock(line_104_clock),
    .reset(line_104_reset),
    .valid(line_104_valid)
  );
  GEN_w1_line #(.COVER_INDEX(105)) line_105 (
    .clock(line_105_clock),
    .reset(line_105_reset),
    .valid(line_105_valid)
  );
  GEN_w1_line #(.COVER_INDEX(106)) line_106 (
    .clock(line_106_clock),
    .reset(line_106_reset),
    .valid(line_106_valid)
  );
  GEN_w1_line #(.COVER_INDEX(107)) line_107 (
    .clock(line_107_clock),
    .reset(line_107_reset),
    .valid(line_107_valid)
  );
  GEN_w1_line #(.COVER_INDEX(108)) line_108 (
    .clock(line_108_clock),
    .reset(line_108_reset),
    .valid(line_108_valid)
  );
  GEN_w1_line #(.COVER_INDEX(109)) line_109 (
    .clock(line_109_clock),
    .reset(line_109_reset),
    .valid(line_109_valid)
  );
  GEN_w1_line #(.COVER_INDEX(110)) line_110 (
    .clock(line_110_clock),
    .reset(line_110_reset),
    .valid(line_110_valid)
  );
  GEN_w1_line #(.COVER_INDEX(111)) line_111 (
    .clock(line_111_clock),
    .reset(line_111_reset),
    .valid(line_111_valid)
  );
  GEN_w1_line #(.COVER_INDEX(112)) line_112 (
    .clock(line_112_clock),
    .reset(line_112_reset),
    .valid(line_112_valid)
  );
  GEN_w1_line #(.COVER_INDEX(113)) line_113 (
    .clock(line_113_clock),
    .reset(line_113_reset),
    .valid(line_113_valid)
  );
  GEN_w1_line #(.COVER_INDEX(114)) line_114 (
    .clock(line_114_clock),
    .reset(line_114_reset),
    .valid(line_114_valid)
  );
  GEN_w1_line #(.COVER_INDEX(115)) line_115 (
    .clock(line_115_clock),
    .reset(line_115_reset),
    .valid(line_115_valid)
  );
  GEN_w1_line #(.COVER_INDEX(116)) line_116 (
    .clock(line_116_clock),
    .reset(line_116_reset),
    .valid(line_116_valid)
  );
  GEN_w1_line #(.COVER_INDEX(117)) line_117 (
    .clock(line_117_clock),
    .reset(line_117_reset),
    .valid(line_117_valid)
  );
  GEN_w1_line #(.COVER_INDEX(118)) line_118 (
    .clock(line_118_clock),
    .reset(line_118_reset),
    .valid(line_118_valid)
  );
  GEN_w1_line #(.COVER_INDEX(119)) line_119 (
    .clock(line_119_clock),
    .reset(line_119_reset),
    .valid(line_119_valid)
  );
  GEN_w1_line #(.COVER_INDEX(120)) line_120 (
    .clock(line_120_clock),
    .reset(line_120_reset),
    .valid(line_120_valid)
  );
  GEN_w1_line #(.COVER_INDEX(121)) line_121 (
    .clock(line_121_clock),
    .reset(line_121_reset),
    .valid(line_121_valid)
  );
  GEN_w1_line #(.COVER_INDEX(122)) line_122 (
    .clock(line_122_clock),
    .reset(line_122_reset),
    .valid(line_122_valid)
  );
  GEN_w1_line #(.COVER_INDEX(123)) line_123 (
    .clock(line_123_clock),
    .reset(line_123_reset),
    .valid(line_123_valid)
  );
  GEN_w1_line #(.COVER_INDEX(124)) line_124 (
    .clock(line_124_clock),
    .reset(line_124_reset),
    .valid(line_124_valid)
  );
  GEN_w1_line #(.COVER_INDEX(125)) line_125 (
    .clock(line_125_clock),
    .reset(line_125_reset),
    .valid(line_125_valid)
  );
  GEN_w1_line #(.COVER_INDEX(126)) line_126 (
    .clock(line_126_clock),
    .reset(line_126_reset),
    .valid(line_126_valid)
  );
  GEN_w1_line #(.COVER_INDEX(127)) line_127 (
    .clock(line_127_clock),
    .reset(line_127_reset),
    .valid(line_127_valid)
  );
  GEN_w1_line #(.COVER_INDEX(128)) line_128 (
    .clock(line_128_clock),
    .reset(line_128_reset),
    .valid(line_128_valid)
  );
  GEN_w1_line #(.COVER_INDEX(129)) line_129 (
    .clock(line_129_clock),
    .reset(line_129_reset),
    .valid(line_129_valid)
  );
  GEN_w1_line #(.COVER_INDEX(130)) line_130 (
    .clock(line_130_clock),
    .reset(line_130_reset),
    .valid(line_130_valid)
  );
  GEN_w1_line #(.COVER_INDEX(131)) line_131 (
    .clock(line_131_clock),
    .reset(line_131_reset),
    .valid(line_131_valid)
  );
  GEN_w1_line #(.COVER_INDEX(132)) line_132 (
    .clock(line_132_clock),
    .reset(line_132_reset),
    .valid(line_132_valid)
  );
  GEN_w1_line #(.COVER_INDEX(133)) line_133 (
    .clock(line_133_clock),
    .reset(line_133_reset),
    .valid(line_133_valid)
  );
  GEN_w1_line #(.COVER_INDEX(134)) line_134 (
    .clock(line_134_clock),
    .reset(line_134_reset),
    .valid(line_134_valid)
  );
  GEN_w1_line #(.COVER_INDEX(135)) line_135 (
    .clock(line_135_clock),
    .reset(line_135_reset),
    .valid(line_135_valid)
  );
  GEN_w1_line #(.COVER_INDEX(136)) line_136 (
    .clock(line_136_clock),
    .reset(line_136_reset),
    .valid(line_136_valid)
  );
  GEN_w1_line #(.COVER_INDEX(137)) line_137 (
    .clock(line_137_clock),
    .reset(line_137_reset),
    .valid(line_137_valid)
  );
  GEN_w1_line #(.COVER_INDEX(138)) line_138 (
    .clock(line_138_clock),
    .reset(line_138_reset),
    .valid(line_138_valid)
  );
  GEN_w1_line #(.COVER_INDEX(139)) line_139 (
    .clock(line_139_clock),
    .reset(line_139_reset),
    .valid(line_139_valid)
  );
  GEN_w1_line #(.COVER_INDEX(140)) line_140 (
    .clock(line_140_clock),
    .reset(line_140_reset),
    .valid(line_140_valid)
  );
  GEN_w1_line #(.COVER_INDEX(141)) line_141 (
    .clock(line_141_clock),
    .reset(line_141_reset),
    .valid(line_141_valid)
  );
  GEN_w1_line #(.COVER_INDEX(142)) line_142 (
    .clock(line_142_clock),
    .reset(line_142_reset),
    .valid(line_142_valid)
  );
  GEN_w1_line #(.COVER_INDEX(143)) line_143 (
    .clock(line_143_clock),
    .reset(line_143_reset),
    .valid(line_143_valid)
  );
  GEN_w1_line #(.COVER_INDEX(144)) line_144 (
    .clock(line_144_clock),
    .reset(line_144_reset),
    .valid(line_144_valid)
  );
  GEN_w1_line #(.COVER_INDEX(145)) line_145 (
    .clock(line_145_clock),
    .reset(line_145_reset),
    .valid(line_145_valid)
  );
  GEN_w1_line #(.COVER_INDEX(146)) line_146 (
    .clock(line_146_clock),
    .reset(line_146_reset),
    .valid(line_146_valid)
  );
  GEN_w1_line #(.COVER_INDEX(147)) line_147 (
    .clock(line_147_clock),
    .reset(line_147_reset),
    .valid(line_147_valid)
  );
  GEN_w1_line #(.COVER_INDEX(148)) line_148 (
    .clock(line_148_clock),
    .reset(line_148_reset),
    .valid(line_148_valid)
  );
  GEN_w1_line #(.COVER_INDEX(149)) line_149 (
    .clock(line_149_clock),
    .reset(line_149_reset),
    .valid(line_149_valid)
  );
  GEN_w1_line #(.COVER_INDEX(150)) line_150 (
    .clock(line_150_clock),
    .reset(line_150_reset),
    .valid(line_150_valid)
  );
  GEN_w1_line #(.COVER_INDEX(151)) line_151 (
    .clock(line_151_clock),
    .reset(line_151_reset),
    .valid(line_151_valid)
  );
  GEN_w1_line #(.COVER_INDEX(152)) line_152 (
    .clock(line_152_clock),
    .reset(line_152_reset),
    .valid(line_152_valid)
  );
  GEN_w1_line #(.COVER_INDEX(153)) line_153 (
    .clock(line_153_clock),
    .reset(line_153_reset),
    .valid(line_153_valid)
  );
  GEN_w1_line #(.COVER_INDEX(154)) line_154 (
    .clock(line_154_clock),
    .reset(line_154_reset),
    .valid(line_154_valid)
  );
  GEN_w1_line #(.COVER_INDEX(155)) line_155 (
    .clock(line_155_clock),
    .reset(line_155_reset),
    .valid(line_155_valid)
  );
  GEN_w1_line #(.COVER_INDEX(156)) line_156 (
    .clock(line_156_clock),
    .reset(line_156_reset),
    .valid(line_156_valid)
  );
  GEN_w1_line #(.COVER_INDEX(157)) line_157 (
    .clock(line_157_clock),
    .reset(line_157_reset),
    .valid(line_157_valid)
  );
  GEN_w1_line #(.COVER_INDEX(158)) line_158 (
    .clock(line_158_clock),
    .reset(line_158_reset),
    .valid(line_158_valid)
  );
  GEN_w1_line #(.COVER_INDEX(159)) line_159 (
    .clock(line_159_clock),
    .reset(line_159_reset),
    .valid(line_159_valid)
  );
  GEN_w1_line #(.COVER_INDEX(160)) line_160 (
    .clock(line_160_clock),
    .reset(line_160_reset),
    .valid(line_160_valid)
  );
  GEN_w1_line #(.COVER_INDEX(161)) line_161 (
    .clock(line_161_clock),
    .reset(line_161_reset),
    .valid(line_161_valid)
  );
  GEN_w1_line #(.COVER_INDEX(162)) line_162 (
    .clock(line_162_clock),
    .reset(line_162_reset),
    .valid(line_162_valid)
  );
  GEN_w1_line #(.COVER_INDEX(163)) line_163 (
    .clock(line_163_clock),
    .reset(line_163_reset),
    .valid(line_163_valid)
  );
  GEN_w1_line #(.COVER_INDEX(164)) line_164 (
    .clock(line_164_clock),
    .reset(line_164_reset),
    .valid(line_164_valid)
  );
  GEN_w1_line #(.COVER_INDEX(165)) line_165 (
    .clock(line_165_clock),
    .reset(line_165_reset),
    .valid(line_165_valid)
  );
  GEN_w1_line #(.COVER_INDEX(166)) line_166 (
    .clock(line_166_clock),
    .reset(line_166_reset),
    .valid(line_166_valid)
  );
  GEN_w1_line #(.COVER_INDEX(167)) line_167 (
    .clock(line_167_clock),
    .reset(line_167_reset),
    .valid(line_167_valid)
  );
  GEN_w1_line #(.COVER_INDEX(168)) line_168 (
    .clock(line_168_clock),
    .reset(line_168_reset),
    .valid(line_168_valid)
  );
  GEN_w1_line #(.COVER_INDEX(169)) line_169 (
    .clock(line_169_clock),
    .reset(line_169_reset),
    .valid(line_169_valid)
  );
  GEN_w1_line #(.COVER_INDEX(170)) line_170 (
    .clock(line_170_clock),
    .reset(line_170_reset),
    .valid(line_170_valid)
  );
  GEN_w1_line #(.COVER_INDEX(171)) line_171 (
    .clock(line_171_clock),
    .reset(line_171_reset),
    .valid(line_171_valid)
  );
  GEN_w1_line #(.COVER_INDEX(172)) line_172 (
    .clock(line_172_clock),
    .reset(line_172_reset),
    .valid(line_172_valid)
  );
  GEN_w1_line #(.COVER_INDEX(173)) line_173 (
    .clock(line_173_clock),
    .reset(line_173_reset),
    .valid(line_173_valid)
  );
  GEN_w1_line #(.COVER_INDEX(174)) line_174 (
    .clock(line_174_clock),
    .reset(line_174_reset),
    .valid(line_174_valid)
  );
  GEN_w1_line #(.COVER_INDEX(175)) line_175 (
    .clock(line_175_clock),
    .reset(line_175_reset),
    .valid(line_175_valid)
  );
  GEN_w1_line #(.COVER_INDEX(176)) line_176 (
    .clock(line_176_clock),
    .reset(line_176_reset),
    .valid(line_176_valid)
  );
  GEN_w1_line #(.COVER_INDEX(177)) line_177 (
    .clock(line_177_clock),
    .reset(line_177_reset),
    .valid(line_177_valid)
  );
  GEN_w1_line #(.COVER_INDEX(178)) line_178 (
    .clock(line_178_clock),
    .reset(line_178_reset),
    .valid(line_178_valid)
  );
  GEN_w1_line #(.COVER_INDEX(179)) line_179 (
    .clock(line_179_clock),
    .reset(line_179_reset),
    .valid(line_179_valid)
  );
  GEN_w1_line #(.COVER_INDEX(180)) line_180 (
    .clock(line_180_clock),
    .reset(line_180_reset),
    .valid(line_180_valid)
  );
  GEN_w1_line #(.COVER_INDEX(181)) line_181 (
    .clock(line_181_clock),
    .reset(line_181_reset),
    .valid(line_181_valid)
  );
  GEN_w1_line #(.COVER_INDEX(182)) line_182 (
    .clock(line_182_clock),
    .reset(line_182_reset),
    .valid(line_182_valid)
  );
  GEN_w1_line #(.COVER_INDEX(183)) line_183 (
    .clock(line_183_clock),
    .reset(line_183_reset),
    .valid(line_183_valid)
  );
  GEN_w1_line #(.COVER_INDEX(184)) line_184 (
    .clock(line_184_clock),
    .reset(line_184_reset),
    .valid(line_184_valid)
  );
  GEN_w1_line #(.COVER_INDEX(185)) line_185 (
    .clock(line_185_clock),
    .reset(line_185_reset),
    .valid(line_185_valid)
  );
  GEN_w1_line #(.COVER_INDEX(186)) line_186 (
    .clock(line_186_clock),
    .reset(line_186_reset),
    .valid(line_186_valid)
  );
  GEN_w1_line #(.COVER_INDEX(187)) line_187 (
    .clock(line_187_clock),
    .reset(line_187_reset),
    .valid(line_187_valid)
  );
  GEN_w1_line #(.COVER_INDEX(188)) line_188 (
    .clock(line_188_clock),
    .reset(line_188_reset),
    .valid(line_188_valid)
  );
  GEN_w1_line #(.COVER_INDEX(189)) line_189 (
    .clock(line_189_clock),
    .reset(line_189_reset),
    .valid(line_189_valid)
  );
  GEN_w1_line #(.COVER_INDEX(190)) line_190 (
    .clock(line_190_clock),
    .reset(line_190_reset),
    .valid(line_190_valid)
  );
  GEN_w1_line #(.COVER_INDEX(191)) line_191 (
    .clock(line_191_clock),
    .reset(line_191_reset),
    .valid(line_191_valid)
  );
  GEN_w1_line #(.COVER_INDEX(192)) line_192 (
    .clock(line_192_clock),
    .reset(line_192_reset),
    .valid(line_192_valid)
  );
  GEN_w1_line #(.COVER_INDEX(193)) line_193 (
    .clock(line_193_clock),
    .reset(line_193_reset),
    .valid(line_193_valid)
  );
  GEN_w1_line #(.COVER_INDEX(194)) line_194 (
    .clock(line_194_clock),
    .reset(line_194_reset),
    .valid(line_194_valid)
  );
  GEN_w1_line #(.COVER_INDEX(195)) line_195 (
    .clock(line_195_clock),
    .reset(line_195_reset),
    .valid(line_195_valid)
  );
  GEN_w1_line #(.COVER_INDEX(196)) line_196 (
    .clock(line_196_clock),
    .reset(line_196_reset),
    .valid(line_196_valid)
  );
  GEN_w1_line #(.COVER_INDEX(197)) line_197 (
    .clock(line_197_clock),
    .reset(line_197_reset),
    .valid(line_197_valid)
  );
  GEN_w1_line #(.COVER_INDEX(198)) line_198 (
    .clock(line_198_clock),
    .reset(line_198_reset),
    .valid(line_198_valid)
  );
  GEN_w1_line #(.COVER_INDEX(199)) line_199 (
    .clock(line_199_clock),
    .reset(line_199_reset),
    .valid(line_199_valid)
  );
  GEN_w1_line #(.COVER_INDEX(200)) line_200 (
    .clock(line_200_clock),
    .reset(line_200_reset),
    .valid(line_200_valid)
  );
  GEN_w1_line #(.COVER_INDEX(201)) line_201 (
    .clock(line_201_clock),
    .reset(line_201_reset),
    .valid(line_201_valid)
  );
  GEN_w1_line #(.COVER_INDEX(202)) line_202 (
    .clock(line_202_clock),
    .reset(line_202_reset),
    .valid(line_202_valid)
  );
  GEN_w1_line #(.COVER_INDEX(203)) line_203 (
    .clock(line_203_clock),
    .reset(line_203_reset),
    .valid(line_203_valid)
  );
  GEN_w1_line #(.COVER_INDEX(204)) line_204 (
    .clock(line_204_clock),
    .reset(line_204_reset),
    .valid(line_204_valid)
  );
  GEN_w1_line #(.COVER_INDEX(205)) line_205 (
    .clock(line_205_clock),
    .reset(line_205_reset),
    .valid(line_205_valid)
  );
  GEN_w1_line #(.COVER_INDEX(206)) line_206 (
    .clock(line_206_clock),
    .reset(line_206_reset),
    .valid(line_206_valid)
  );
  GEN_w1_line #(.COVER_INDEX(207)) line_207 (
    .clock(line_207_clock),
    .reset(line_207_reset),
    .valid(line_207_valid)
  );
  GEN_w1_line #(.COVER_INDEX(208)) line_208 (
    .clock(line_208_clock),
    .reset(line_208_reset),
    .valid(line_208_valid)
  );
  GEN_w1_line #(.COVER_INDEX(209)) line_209 (
    .clock(line_209_clock),
    .reset(line_209_reset),
    .valid(line_209_valid)
  );
  GEN_w1_line #(.COVER_INDEX(210)) line_210 (
    .clock(line_210_clock),
    .reset(line_210_reset),
    .valid(line_210_valid)
  );
  GEN_w1_line #(.COVER_INDEX(211)) line_211 (
    .clock(line_211_clock),
    .reset(line_211_reset),
    .valid(line_211_valid)
  );
  GEN_w1_line #(.COVER_INDEX(212)) line_212 (
    .clock(line_212_clock),
    .reset(line_212_reset),
    .valid(line_212_valid)
  );
  GEN_w1_line #(.COVER_INDEX(213)) line_213 (
    .clock(line_213_clock),
    .reset(line_213_reset),
    .valid(line_213_valid)
  );
  GEN_w1_line #(.COVER_INDEX(214)) line_214 (
    .clock(line_214_clock),
    .reset(line_214_reset),
    .valid(line_214_valid)
  );
  assign line_43_clock = clock;
  assign line_43_reset = reset;
  assign line_43_valid = 3'h0 == _io_out_s_funct_T_2 ^ line_43_valid_reg;
  assign line_44_clock = clock;
  assign line_44_reset = reset;
  assign line_44_valid = 3'h1 == _io_out_s_funct_T_2 ^ line_44_valid_reg;
  assign line_45_clock = clock;
  assign line_45_reset = reset;
  assign line_45_valid = 3'h2 == _io_out_s_funct_T_2 ^ line_45_valid_reg;
  assign line_46_clock = clock;
  assign line_46_reset = reset;
  assign line_46_valid = 3'h3 == _io_out_s_funct_T_2 ^ line_46_valid_reg;
  assign line_47_clock = clock;
  assign line_47_reset = reset;
  assign line_47_valid = 3'h4 == _io_out_s_funct_T_2 ^ line_47_valid_reg;
  assign line_48_clock = clock;
  assign line_48_reset = reset;
  assign line_48_valid = 3'h5 == _io_out_s_funct_T_2 ^ line_48_valid_reg;
  assign line_49_clock = clock;
  assign line_49_reset = reset;
  assign line_49_valid = 3'h6 == _io_out_s_funct_T_2 ^ line_49_valid_reg;
  assign line_50_clock = clock;
  assign line_50_reset = reset;
  assign line_50_valid = 3'h7 == _io_out_s_funct_T_2 ^ line_50_valid_reg;
  assign line_51_clock = clock;
  assign line_51_reset = reset;
  assign line_51_valid = 2'h0 == io_in[11:10] ^ line_51_valid_reg;
  assign line_52_clock = clock;
  assign line_52_reset = reset;
  assign line_52_valid = 2'h1 == io_in[11:10] ^ line_52_valid_reg;
  assign line_53_clock = clock;
  assign line_53_reset = reset;
  assign line_53_valid = 2'h2 == io_in[11:10] ^ line_53_valid_reg;
  assign line_54_clock = clock;
  assign line_54_reset = reset;
  assign line_54_valid = 2'h3 == io_in[11:10] ^ line_54_valid_reg;
  assign line_55_clock = clock;
  assign line_55_reset = reset;
  assign line_55_valid = 5'h0 == _io_out_T_2 ^ line_55_valid_reg;
  assign line_56_clock = clock;
  assign line_56_reset = reset;
  assign line_56_valid = 5'h1 == _io_out_T_2 ^ line_56_valid_reg;
  assign line_57_clock = clock;
  assign line_57_reset = reset;
  assign line_57_valid = 5'h2 == _io_out_T_2 ^ line_57_valid_reg;
  assign line_58_clock = clock;
  assign line_58_reset = reset;
  assign line_58_valid = 5'h3 == _io_out_T_2 ^ line_58_valid_reg;
  assign line_59_clock = clock;
  assign line_59_reset = reset;
  assign line_59_valid = 5'h4 == _io_out_T_2 ^ line_59_valid_reg;
  assign line_60_clock = clock;
  assign line_60_reset = reset;
  assign line_60_valid = 5'h5 == _io_out_T_2 ^ line_60_valid_reg;
  assign line_61_clock = clock;
  assign line_61_reset = reset;
  assign line_61_valid = 5'h6 == _io_out_T_2 ^ line_61_valid_reg;
  assign line_62_clock = clock;
  assign line_62_reset = reset;
  assign line_62_valid = 5'h7 == _io_out_T_2 ^ line_62_valid_reg;
  assign line_63_clock = clock;
  assign line_63_reset = reset;
  assign line_63_valid = 5'h8 == _io_out_T_2 ^ line_63_valid_reg;
  assign line_64_clock = clock;
  assign line_64_reset = reset;
  assign line_64_valid = 5'h9 == _io_out_T_2 ^ line_64_valid_reg;
  assign line_65_clock = clock;
  assign line_65_reset = reset;
  assign line_65_valid = 5'ha == _io_out_T_2 ^ line_65_valid_reg;
  assign line_66_clock = clock;
  assign line_66_reset = reset;
  assign line_66_valid = 5'hb == _io_out_T_2 ^ line_66_valid_reg;
  assign line_67_clock = clock;
  assign line_67_reset = reset;
  assign line_67_valid = 5'hc == _io_out_T_2 ^ line_67_valid_reg;
  assign line_68_clock = clock;
  assign line_68_reset = reset;
  assign line_68_valid = 5'hd == _io_out_T_2 ^ line_68_valid_reg;
  assign line_69_clock = clock;
  assign line_69_reset = reset;
  assign line_69_valid = 5'he == _io_out_T_2 ^ line_69_valid_reg;
  assign line_70_clock = clock;
  assign line_70_reset = reset;
  assign line_70_valid = 5'hf == _io_out_T_2 ^ line_70_valid_reg;
  assign line_71_clock = clock;
  assign line_71_reset = reset;
  assign line_71_valid = 5'h10 == _io_out_T_2 ^ line_71_valid_reg;
  assign line_72_clock = clock;
  assign line_72_reset = reset;
  assign line_72_valid = 5'h11 == _io_out_T_2 ^ line_72_valid_reg;
  assign line_73_clock = clock;
  assign line_73_reset = reset;
  assign line_73_valid = 5'h12 == _io_out_T_2 ^ line_73_valid_reg;
  assign line_74_clock = clock;
  assign line_74_reset = reset;
  assign line_74_valid = 5'h13 == _io_out_T_2 ^ line_74_valid_reg;
  assign line_75_clock = clock;
  assign line_75_reset = reset;
  assign line_75_valid = 5'h14 == _io_out_T_2 ^ line_75_valid_reg;
  assign line_76_clock = clock;
  assign line_76_reset = reset;
  assign line_76_valid = 5'h15 == _io_out_T_2 ^ line_76_valid_reg;
  assign line_77_clock = clock;
  assign line_77_reset = reset;
  assign line_77_valid = 5'h16 == _io_out_T_2 ^ line_77_valid_reg;
  assign line_78_clock = clock;
  assign line_78_reset = reset;
  assign line_78_valid = 5'h17 == _io_out_T_2 ^ line_78_valid_reg;
  assign line_79_clock = clock;
  assign line_79_reset = reset;
  assign line_79_valid = 5'h18 == _io_out_T_2 ^ line_79_valid_reg;
  assign line_80_clock = clock;
  assign line_80_reset = reset;
  assign line_80_valid = 5'h19 == _io_out_T_2 ^ line_80_valid_reg;
  assign line_81_clock = clock;
  assign line_81_reset = reset;
  assign line_81_valid = 5'h1a == _io_out_T_2 ^ line_81_valid_reg;
  assign line_82_clock = clock;
  assign line_82_reset = reset;
  assign line_82_valid = 5'h1b == _io_out_T_2 ^ line_82_valid_reg;
  assign line_83_clock = clock;
  assign line_83_reset = reset;
  assign line_83_valid = 5'h1c == _io_out_T_2 ^ line_83_valid_reg;
  assign line_84_clock = clock;
  assign line_84_reset = reset;
  assign line_84_valid = 5'h1d == _io_out_T_2 ^ line_84_valid_reg;
  assign line_85_clock = clock;
  assign line_85_reset = reset;
  assign line_85_valid = 5'h1e == _io_out_T_2 ^ line_85_valid_reg;
  assign line_86_clock = clock;
  assign line_86_reset = reset;
  assign line_86_valid = 5'h1f == _io_out_T_2 ^ line_86_valid_reg;
  assign line_87_clock = clock;
  assign line_87_reset = reset;
  assign line_87_valid = 5'h0 == _io_out_T_2 ^ line_87_valid_reg;
  assign line_88_clock = clock;
  assign line_88_reset = reset;
  assign line_88_valid = 5'h1 == _io_out_T_2 ^ line_88_valid_reg;
  assign line_89_clock = clock;
  assign line_89_reset = reset;
  assign line_89_valid = 5'h2 == _io_out_T_2 ^ line_89_valid_reg;
  assign line_90_clock = clock;
  assign line_90_reset = reset;
  assign line_90_valid = 5'h3 == _io_out_T_2 ^ line_90_valid_reg;
  assign line_91_clock = clock;
  assign line_91_reset = reset;
  assign line_91_valid = 5'h4 == _io_out_T_2 ^ line_91_valid_reg;
  assign line_92_clock = clock;
  assign line_92_reset = reset;
  assign line_92_valid = 5'h5 == _io_out_T_2 ^ line_92_valid_reg;
  assign line_93_clock = clock;
  assign line_93_reset = reset;
  assign line_93_valid = 5'h6 == _io_out_T_2 ^ line_93_valid_reg;
  assign line_94_clock = clock;
  assign line_94_reset = reset;
  assign line_94_valid = 5'h7 == _io_out_T_2 ^ line_94_valid_reg;
  assign line_95_clock = clock;
  assign line_95_reset = reset;
  assign line_95_valid = 5'h8 == _io_out_T_2 ^ line_95_valid_reg;
  assign line_96_clock = clock;
  assign line_96_reset = reset;
  assign line_96_valid = 5'h9 == _io_out_T_2 ^ line_96_valid_reg;
  assign line_97_clock = clock;
  assign line_97_reset = reset;
  assign line_97_valid = 5'ha == _io_out_T_2 ^ line_97_valid_reg;
  assign line_98_clock = clock;
  assign line_98_reset = reset;
  assign line_98_valid = 5'hb == _io_out_T_2 ^ line_98_valid_reg;
  assign line_99_clock = clock;
  assign line_99_reset = reset;
  assign line_99_valid = 5'hc == _io_out_T_2 ^ line_99_valid_reg;
  assign line_100_clock = clock;
  assign line_100_reset = reset;
  assign line_100_valid = 5'hd == _io_out_T_2 ^ line_100_valid_reg;
  assign line_101_clock = clock;
  assign line_101_reset = reset;
  assign line_101_valid = 5'he == _io_out_T_2 ^ line_101_valid_reg;
  assign line_102_clock = clock;
  assign line_102_reset = reset;
  assign line_102_valid = 5'hf == _io_out_T_2 ^ line_102_valid_reg;
  assign line_103_clock = clock;
  assign line_103_reset = reset;
  assign line_103_valid = 5'h10 == _io_out_T_2 ^ line_103_valid_reg;
  assign line_104_clock = clock;
  assign line_104_reset = reset;
  assign line_104_valid = 5'h11 == _io_out_T_2 ^ line_104_valid_reg;
  assign line_105_clock = clock;
  assign line_105_reset = reset;
  assign line_105_valid = 5'h12 == _io_out_T_2 ^ line_105_valid_reg;
  assign line_106_clock = clock;
  assign line_106_reset = reset;
  assign line_106_valid = 5'h13 == _io_out_T_2 ^ line_106_valid_reg;
  assign line_107_clock = clock;
  assign line_107_reset = reset;
  assign line_107_valid = 5'h14 == _io_out_T_2 ^ line_107_valid_reg;
  assign line_108_clock = clock;
  assign line_108_reset = reset;
  assign line_108_valid = 5'h15 == _io_out_T_2 ^ line_108_valid_reg;
  assign line_109_clock = clock;
  assign line_109_reset = reset;
  assign line_109_valid = 5'h16 == _io_out_T_2 ^ line_109_valid_reg;
  assign line_110_clock = clock;
  assign line_110_reset = reset;
  assign line_110_valid = 5'h17 == _io_out_T_2 ^ line_110_valid_reg;
  assign line_111_clock = clock;
  assign line_111_reset = reset;
  assign line_111_valid = 5'h18 == _io_out_T_2 ^ line_111_valid_reg;
  assign line_112_clock = clock;
  assign line_112_reset = reset;
  assign line_112_valid = 5'h19 == _io_out_T_2 ^ line_112_valid_reg;
  assign line_113_clock = clock;
  assign line_113_reset = reset;
  assign line_113_valid = 5'h1a == _io_out_T_2 ^ line_113_valid_reg;
  assign line_114_clock = clock;
  assign line_114_reset = reset;
  assign line_114_valid = 5'h1b == _io_out_T_2 ^ line_114_valid_reg;
  assign line_115_clock = clock;
  assign line_115_reset = reset;
  assign line_115_valid = 5'h1c == _io_out_T_2 ^ line_115_valid_reg;
  assign line_116_clock = clock;
  assign line_116_reset = reset;
  assign line_116_valid = 5'h1d == _io_out_T_2 ^ line_116_valid_reg;
  assign line_117_clock = clock;
  assign line_117_reset = reset;
  assign line_117_valid = 5'h1e == _io_out_T_2 ^ line_117_valid_reg;
  assign line_118_clock = clock;
  assign line_118_reset = reset;
  assign line_118_valid = 5'h1f == _io_out_T_2 ^ line_118_valid_reg;
  assign line_119_clock = clock;
  assign line_119_reset = reset;
  assign line_119_valid = 5'h0 == _io_out_T_2 ^ line_119_valid_reg;
  assign line_120_clock = clock;
  assign line_120_reset = reset;
  assign line_120_valid = 5'h1 == _io_out_T_2 ^ line_120_valid_reg;
  assign line_121_clock = clock;
  assign line_121_reset = reset;
  assign line_121_valid = 5'h2 == _io_out_T_2 ^ line_121_valid_reg;
  assign line_122_clock = clock;
  assign line_122_reset = reset;
  assign line_122_valid = 5'h3 == _io_out_T_2 ^ line_122_valid_reg;
  assign line_123_clock = clock;
  assign line_123_reset = reset;
  assign line_123_valid = 5'h4 == _io_out_T_2 ^ line_123_valid_reg;
  assign line_124_clock = clock;
  assign line_124_reset = reset;
  assign line_124_valid = 5'h5 == _io_out_T_2 ^ line_124_valid_reg;
  assign line_125_clock = clock;
  assign line_125_reset = reset;
  assign line_125_valid = 5'h6 == _io_out_T_2 ^ line_125_valid_reg;
  assign line_126_clock = clock;
  assign line_126_reset = reset;
  assign line_126_valid = 5'h7 == _io_out_T_2 ^ line_126_valid_reg;
  assign line_127_clock = clock;
  assign line_127_reset = reset;
  assign line_127_valid = 5'h8 == _io_out_T_2 ^ line_127_valid_reg;
  assign line_128_clock = clock;
  assign line_128_reset = reset;
  assign line_128_valid = 5'h9 == _io_out_T_2 ^ line_128_valid_reg;
  assign line_129_clock = clock;
  assign line_129_reset = reset;
  assign line_129_valid = 5'ha == _io_out_T_2 ^ line_129_valid_reg;
  assign line_130_clock = clock;
  assign line_130_reset = reset;
  assign line_130_valid = 5'hb == _io_out_T_2 ^ line_130_valid_reg;
  assign line_131_clock = clock;
  assign line_131_reset = reset;
  assign line_131_valid = 5'hc == _io_out_T_2 ^ line_131_valid_reg;
  assign line_132_clock = clock;
  assign line_132_reset = reset;
  assign line_132_valid = 5'hd == _io_out_T_2 ^ line_132_valid_reg;
  assign line_133_clock = clock;
  assign line_133_reset = reset;
  assign line_133_valid = 5'he == _io_out_T_2 ^ line_133_valid_reg;
  assign line_134_clock = clock;
  assign line_134_reset = reset;
  assign line_134_valid = 5'hf == _io_out_T_2 ^ line_134_valid_reg;
  assign line_135_clock = clock;
  assign line_135_reset = reset;
  assign line_135_valid = 5'h10 == _io_out_T_2 ^ line_135_valid_reg;
  assign line_136_clock = clock;
  assign line_136_reset = reset;
  assign line_136_valid = 5'h11 == _io_out_T_2 ^ line_136_valid_reg;
  assign line_137_clock = clock;
  assign line_137_reset = reset;
  assign line_137_valid = 5'h12 == _io_out_T_2 ^ line_137_valid_reg;
  assign line_138_clock = clock;
  assign line_138_reset = reset;
  assign line_138_valid = 5'h13 == _io_out_T_2 ^ line_138_valid_reg;
  assign line_139_clock = clock;
  assign line_139_reset = reset;
  assign line_139_valid = 5'h14 == _io_out_T_2 ^ line_139_valid_reg;
  assign line_140_clock = clock;
  assign line_140_reset = reset;
  assign line_140_valid = 5'h15 == _io_out_T_2 ^ line_140_valid_reg;
  assign line_141_clock = clock;
  assign line_141_reset = reset;
  assign line_141_valid = 5'h16 == _io_out_T_2 ^ line_141_valid_reg;
  assign line_142_clock = clock;
  assign line_142_reset = reset;
  assign line_142_valid = 5'h17 == _io_out_T_2 ^ line_142_valid_reg;
  assign line_143_clock = clock;
  assign line_143_reset = reset;
  assign line_143_valid = 5'h18 == _io_out_T_2 ^ line_143_valid_reg;
  assign line_144_clock = clock;
  assign line_144_reset = reset;
  assign line_144_valid = 5'h19 == _io_out_T_2 ^ line_144_valid_reg;
  assign line_145_clock = clock;
  assign line_145_reset = reset;
  assign line_145_valid = 5'h1a == _io_out_T_2 ^ line_145_valid_reg;
  assign line_146_clock = clock;
  assign line_146_reset = reset;
  assign line_146_valid = 5'h1b == _io_out_T_2 ^ line_146_valid_reg;
  assign line_147_clock = clock;
  assign line_147_reset = reset;
  assign line_147_valid = 5'h1c == _io_out_T_2 ^ line_147_valid_reg;
  assign line_148_clock = clock;
  assign line_148_reset = reset;
  assign line_148_valid = 5'h1d == _io_out_T_2 ^ line_148_valid_reg;
  assign line_149_clock = clock;
  assign line_149_reset = reset;
  assign line_149_valid = 5'h1e == _io_out_T_2 ^ line_149_valid_reg;
  assign line_150_clock = clock;
  assign line_150_reset = reset;
  assign line_150_valid = 5'h1f == _io_out_T_2 ^ line_150_valid_reg;
  assign line_151_clock = clock;
  assign line_151_reset = reset;
  assign line_151_valid = 5'h0 == _io_out_T_2 ^ line_151_valid_reg;
  assign line_152_clock = clock;
  assign line_152_reset = reset;
  assign line_152_valid = 5'h1 == _io_out_T_2 ^ line_152_valid_reg;
  assign line_153_clock = clock;
  assign line_153_reset = reset;
  assign line_153_valid = 5'h2 == _io_out_T_2 ^ line_153_valid_reg;
  assign line_154_clock = clock;
  assign line_154_reset = reset;
  assign line_154_valid = 5'h3 == _io_out_T_2 ^ line_154_valid_reg;
  assign line_155_clock = clock;
  assign line_155_reset = reset;
  assign line_155_valid = 5'h4 == _io_out_T_2 ^ line_155_valid_reg;
  assign line_156_clock = clock;
  assign line_156_reset = reset;
  assign line_156_valid = 5'h5 == _io_out_T_2 ^ line_156_valid_reg;
  assign line_157_clock = clock;
  assign line_157_reset = reset;
  assign line_157_valid = 5'h6 == _io_out_T_2 ^ line_157_valid_reg;
  assign line_158_clock = clock;
  assign line_158_reset = reset;
  assign line_158_valid = 5'h7 == _io_out_T_2 ^ line_158_valid_reg;
  assign line_159_clock = clock;
  assign line_159_reset = reset;
  assign line_159_valid = 5'h8 == _io_out_T_2 ^ line_159_valid_reg;
  assign line_160_clock = clock;
  assign line_160_reset = reset;
  assign line_160_valid = 5'h9 == _io_out_T_2 ^ line_160_valid_reg;
  assign line_161_clock = clock;
  assign line_161_reset = reset;
  assign line_161_valid = 5'ha == _io_out_T_2 ^ line_161_valid_reg;
  assign line_162_clock = clock;
  assign line_162_reset = reset;
  assign line_162_valid = 5'hb == _io_out_T_2 ^ line_162_valid_reg;
  assign line_163_clock = clock;
  assign line_163_reset = reset;
  assign line_163_valid = 5'hc == _io_out_T_2 ^ line_163_valid_reg;
  assign line_164_clock = clock;
  assign line_164_reset = reset;
  assign line_164_valid = 5'hd == _io_out_T_2 ^ line_164_valid_reg;
  assign line_165_clock = clock;
  assign line_165_reset = reset;
  assign line_165_valid = 5'he == _io_out_T_2 ^ line_165_valid_reg;
  assign line_166_clock = clock;
  assign line_166_reset = reset;
  assign line_166_valid = 5'hf == _io_out_T_2 ^ line_166_valid_reg;
  assign line_167_clock = clock;
  assign line_167_reset = reset;
  assign line_167_valid = 5'h10 == _io_out_T_2 ^ line_167_valid_reg;
  assign line_168_clock = clock;
  assign line_168_reset = reset;
  assign line_168_valid = 5'h11 == _io_out_T_2 ^ line_168_valid_reg;
  assign line_169_clock = clock;
  assign line_169_reset = reset;
  assign line_169_valid = 5'h12 == _io_out_T_2 ^ line_169_valid_reg;
  assign line_170_clock = clock;
  assign line_170_reset = reset;
  assign line_170_valid = 5'h13 == _io_out_T_2 ^ line_170_valid_reg;
  assign line_171_clock = clock;
  assign line_171_reset = reset;
  assign line_171_valid = 5'h14 == _io_out_T_2 ^ line_171_valid_reg;
  assign line_172_clock = clock;
  assign line_172_reset = reset;
  assign line_172_valid = 5'h15 == _io_out_T_2 ^ line_172_valid_reg;
  assign line_173_clock = clock;
  assign line_173_reset = reset;
  assign line_173_valid = 5'h16 == _io_out_T_2 ^ line_173_valid_reg;
  assign line_174_clock = clock;
  assign line_174_reset = reset;
  assign line_174_valid = 5'h17 == _io_out_T_2 ^ line_174_valid_reg;
  assign line_175_clock = clock;
  assign line_175_reset = reset;
  assign line_175_valid = 5'h18 == _io_out_T_2 ^ line_175_valid_reg;
  assign line_176_clock = clock;
  assign line_176_reset = reset;
  assign line_176_valid = 5'h19 == _io_out_T_2 ^ line_176_valid_reg;
  assign line_177_clock = clock;
  assign line_177_reset = reset;
  assign line_177_valid = 5'h1a == _io_out_T_2 ^ line_177_valid_reg;
  assign line_178_clock = clock;
  assign line_178_reset = reset;
  assign line_178_valid = 5'h1b == _io_out_T_2 ^ line_178_valid_reg;
  assign line_179_clock = clock;
  assign line_179_reset = reset;
  assign line_179_valid = 5'h1c == _io_out_T_2 ^ line_179_valid_reg;
  assign line_180_clock = clock;
  assign line_180_reset = reset;
  assign line_180_valid = 5'h1d == _io_out_T_2 ^ line_180_valid_reg;
  assign line_181_clock = clock;
  assign line_181_reset = reset;
  assign line_181_valid = 5'h1e == _io_out_T_2 ^ line_181_valid_reg;
  assign line_182_clock = clock;
  assign line_182_reset = reset;
  assign line_182_valid = 5'h1f == _io_out_T_2 ^ line_182_valid_reg;
  assign line_183_clock = clock;
  assign line_183_reset = reset;
  assign line_183_valid = 5'h0 == _io_out_T_2 ^ line_183_valid_reg;
  assign line_184_clock = clock;
  assign line_184_reset = reset;
  assign line_184_valid = 5'h1 == _io_out_T_2 ^ line_184_valid_reg;
  assign line_185_clock = clock;
  assign line_185_reset = reset;
  assign line_185_valid = 5'h2 == _io_out_T_2 ^ line_185_valid_reg;
  assign line_186_clock = clock;
  assign line_186_reset = reset;
  assign line_186_valid = 5'h3 == _io_out_T_2 ^ line_186_valid_reg;
  assign line_187_clock = clock;
  assign line_187_reset = reset;
  assign line_187_valid = 5'h4 == _io_out_T_2 ^ line_187_valid_reg;
  assign line_188_clock = clock;
  assign line_188_reset = reset;
  assign line_188_valid = 5'h5 == _io_out_T_2 ^ line_188_valid_reg;
  assign line_189_clock = clock;
  assign line_189_reset = reset;
  assign line_189_valid = 5'h6 == _io_out_T_2 ^ line_189_valid_reg;
  assign line_190_clock = clock;
  assign line_190_reset = reset;
  assign line_190_valid = 5'h7 == _io_out_T_2 ^ line_190_valid_reg;
  assign line_191_clock = clock;
  assign line_191_reset = reset;
  assign line_191_valid = 5'h8 == _io_out_T_2 ^ line_191_valid_reg;
  assign line_192_clock = clock;
  assign line_192_reset = reset;
  assign line_192_valid = 5'h9 == _io_out_T_2 ^ line_192_valid_reg;
  assign line_193_clock = clock;
  assign line_193_reset = reset;
  assign line_193_valid = 5'ha == _io_out_T_2 ^ line_193_valid_reg;
  assign line_194_clock = clock;
  assign line_194_reset = reset;
  assign line_194_valid = 5'hb == _io_out_T_2 ^ line_194_valid_reg;
  assign line_195_clock = clock;
  assign line_195_reset = reset;
  assign line_195_valid = 5'hc == _io_out_T_2 ^ line_195_valid_reg;
  assign line_196_clock = clock;
  assign line_196_reset = reset;
  assign line_196_valid = 5'hd == _io_out_T_2 ^ line_196_valid_reg;
  assign line_197_clock = clock;
  assign line_197_reset = reset;
  assign line_197_valid = 5'he == _io_out_T_2 ^ line_197_valid_reg;
  assign line_198_clock = clock;
  assign line_198_reset = reset;
  assign line_198_valid = 5'hf == _io_out_T_2 ^ line_198_valid_reg;
  assign line_199_clock = clock;
  assign line_199_reset = reset;
  assign line_199_valid = 5'h10 == _io_out_T_2 ^ line_199_valid_reg;
  assign line_200_clock = clock;
  assign line_200_reset = reset;
  assign line_200_valid = 5'h11 == _io_out_T_2 ^ line_200_valid_reg;
  assign line_201_clock = clock;
  assign line_201_reset = reset;
  assign line_201_valid = 5'h12 == _io_out_T_2 ^ line_201_valid_reg;
  assign line_202_clock = clock;
  assign line_202_reset = reset;
  assign line_202_valid = 5'h13 == _io_out_T_2 ^ line_202_valid_reg;
  assign line_203_clock = clock;
  assign line_203_reset = reset;
  assign line_203_valid = 5'h14 == _io_out_T_2 ^ line_203_valid_reg;
  assign line_204_clock = clock;
  assign line_204_reset = reset;
  assign line_204_valid = 5'h15 == _io_out_T_2 ^ line_204_valid_reg;
  assign line_205_clock = clock;
  assign line_205_reset = reset;
  assign line_205_valid = 5'h16 == _io_out_T_2 ^ line_205_valid_reg;
  assign line_206_clock = clock;
  assign line_206_reset = reset;
  assign line_206_valid = 5'h17 == _io_out_T_2 ^ line_206_valid_reg;
  assign line_207_clock = clock;
  assign line_207_reset = reset;
  assign line_207_valid = 5'h18 == _io_out_T_2 ^ line_207_valid_reg;
  assign line_208_clock = clock;
  assign line_208_reset = reset;
  assign line_208_valid = 5'h19 == _io_out_T_2 ^ line_208_valid_reg;
  assign line_209_clock = clock;
  assign line_209_reset = reset;
  assign line_209_valid = 5'h1a == _io_out_T_2 ^ line_209_valid_reg;
  assign line_210_clock = clock;
  assign line_210_reset = reset;
  assign line_210_valid = 5'h1b == _io_out_T_2 ^ line_210_valid_reg;
  assign line_211_clock = clock;
  assign line_211_reset = reset;
  assign line_211_valid = 5'h1c == _io_out_T_2 ^ line_211_valid_reg;
  assign line_212_clock = clock;
  assign line_212_reset = reset;
  assign line_212_valid = 5'h1d == _io_out_T_2 ^ line_212_valid_reg;
  assign line_213_clock = clock;
  assign line_213_reset = reset;
  assign line_213_valid = 5'h1e == _io_out_T_2 ^ line_213_valid_reg;
  assign line_214_clock = clock;
  assign line_214_reset = reset;
  assign line_214_valid = 5'h1f == _io_out_T_2 ^ line_214_valid_reg;
  assign io_out_bits = 5'h1f == _io_out_T_2 ? io_in : _GEN_214; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  always @(posedge clock) begin
    line_43_valid_reg <= 3'h0 == _io_out_s_funct_T_2;
    line_44_valid_reg <= 3'h1 == _io_out_s_funct_T_2;
    line_45_valid_reg <= 3'h2 == _io_out_s_funct_T_2;
    line_46_valid_reg <= 3'h3 == _io_out_s_funct_T_2;
    line_47_valid_reg <= 3'h4 == _io_out_s_funct_T_2;
    line_48_valid_reg <= 3'h5 == _io_out_s_funct_T_2;
    line_49_valid_reg <= 3'h6 == _io_out_s_funct_T_2;
    line_50_valid_reg <= 3'h7 == _io_out_s_funct_T_2;
    line_51_valid_reg <= 2'h0 == io_in[11:10];
    line_52_valid_reg <= 2'h1 == io_in[11:10];
    line_53_valid_reg <= 2'h2 == io_in[11:10];
    line_54_valid_reg <= 2'h3 == io_in[11:10];
    line_55_valid_reg <= 5'h0 == _io_out_T_2;
    line_56_valid_reg <= 5'h1 == _io_out_T_2;
    line_57_valid_reg <= 5'h2 == _io_out_T_2;
    line_58_valid_reg <= 5'h3 == _io_out_T_2;
    line_59_valid_reg <= 5'h4 == _io_out_T_2;
    line_60_valid_reg <= 5'h5 == _io_out_T_2;
    line_61_valid_reg <= 5'h6 == _io_out_T_2;
    line_62_valid_reg <= 5'h7 == _io_out_T_2;
    line_63_valid_reg <= 5'h8 == _io_out_T_2;
    line_64_valid_reg <= 5'h9 == _io_out_T_2;
    line_65_valid_reg <= 5'ha == _io_out_T_2;
    line_66_valid_reg <= 5'hb == _io_out_T_2;
    line_67_valid_reg <= 5'hc == _io_out_T_2;
    line_68_valid_reg <= 5'hd == _io_out_T_2;
    line_69_valid_reg <= 5'he == _io_out_T_2;
    line_70_valid_reg <= 5'hf == _io_out_T_2;
    line_71_valid_reg <= 5'h10 == _io_out_T_2;
    line_72_valid_reg <= 5'h11 == _io_out_T_2;
    line_73_valid_reg <= 5'h12 == _io_out_T_2;
    line_74_valid_reg <= 5'h13 == _io_out_T_2;
    line_75_valid_reg <= 5'h14 == _io_out_T_2;
    line_76_valid_reg <= 5'h15 == _io_out_T_2;
    line_77_valid_reg <= 5'h16 == _io_out_T_2;
    line_78_valid_reg <= 5'h17 == _io_out_T_2;
    line_79_valid_reg <= 5'h18 == _io_out_T_2;
    line_80_valid_reg <= 5'h19 == _io_out_T_2;
    line_81_valid_reg <= 5'h1a == _io_out_T_2;
    line_82_valid_reg <= 5'h1b == _io_out_T_2;
    line_83_valid_reg <= 5'h1c == _io_out_T_2;
    line_84_valid_reg <= 5'h1d == _io_out_T_2;
    line_85_valid_reg <= 5'h1e == _io_out_T_2;
    line_86_valid_reg <= 5'h1f == _io_out_T_2;
    line_87_valid_reg <= 5'h0 == _io_out_T_2;
    line_88_valid_reg <= 5'h1 == _io_out_T_2;
    line_89_valid_reg <= 5'h2 == _io_out_T_2;
    line_90_valid_reg <= 5'h3 == _io_out_T_2;
    line_91_valid_reg <= 5'h4 == _io_out_T_2;
    line_92_valid_reg <= 5'h5 == _io_out_T_2;
    line_93_valid_reg <= 5'h6 == _io_out_T_2;
    line_94_valid_reg <= 5'h7 == _io_out_T_2;
    line_95_valid_reg <= 5'h8 == _io_out_T_2;
    line_96_valid_reg <= 5'h9 == _io_out_T_2;
    line_97_valid_reg <= 5'ha == _io_out_T_2;
    line_98_valid_reg <= 5'hb == _io_out_T_2;
    line_99_valid_reg <= 5'hc == _io_out_T_2;
    line_100_valid_reg <= 5'hd == _io_out_T_2;
    line_101_valid_reg <= 5'he == _io_out_T_2;
    line_102_valid_reg <= 5'hf == _io_out_T_2;
    line_103_valid_reg <= 5'h10 == _io_out_T_2;
    line_104_valid_reg <= 5'h11 == _io_out_T_2;
    line_105_valid_reg <= 5'h12 == _io_out_T_2;
    line_106_valid_reg <= 5'h13 == _io_out_T_2;
    line_107_valid_reg <= 5'h14 == _io_out_T_2;
    line_108_valid_reg <= 5'h15 == _io_out_T_2;
    line_109_valid_reg <= 5'h16 == _io_out_T_2;
    line_110_valid_reg <= 5'h17 == _io_out_T_2;
    line_111_valid_reg <= 5'h18 == _io_out_T_2;
    line_112_valid_reg <= 5'h19 == _io_out_T_2;
    line_113_valid_reg <= 5'h1a == _io_out_T_2;
    line_114_valid_reg <= 5'h1b == _io_out_T_2;
    line_115_valid_reg <= 5'h1c == _io_out_T_2;
    line_116_valid_reg <= 5'h1d == _io_out_T_2;
    line_117_valid_reg <= 5'h1e == _io_out_T_2;
    line_118_valid_reg <= 5'h1f == _io_out_T_2;
    line_119_valid_reg <= 5'h0 == _io_out_T_2;
    line_120_valid_reg <= 5'h1 == _io_out_T_2;
    line_121_valid_reg <= 5'h2 == _io_out_T_2;
    line_122_valid_reg <= 5'h3 == _io_out_T_2;
    line_123_valid_reg <= 5'h4 == _io_out_T_2;
    line_124_valid_reg <= 5'h5 == _io_out_T_2;
    line_125_valid_reg <= 5'h6 == _io_out_T_2;
    line_126_valid_reg <= 5'h7 == _io_out_T_2;
    line_127_valid_reg <= 5'h8 == _io_out_T_2;
    line_128_valid_reg <= 5'h9 == _io_out_T_2;
    line_129_valid_reg <= 5'ha == _io_out_T_2;
    line_130_valid_reg <= 5'hb == _io_out_T_2;
    line_131_valid_reg <= 5'hc == _io_out_T_2;
    line_132_valid_reg <= 5'hd == _io_out_T_2;
    line_133_valid_reg <= 5'he == _io_out_T_2;
    line_134_valid_reg <= 5'hf == _io_out_T_2;
    line_135_valid_reg <= 5'h10 == _io_out_T_2;
    line_136_valid_reg <= 5'h11 == _io_out_T_2;
    line_137_valid_reg <= 5'h12 == _io_out_T_2;
    line_138_valid_reg <= 5'h13 == _io_out_T_2;
    line_139_valid_reg <= 5'h14 == _io_out_T_2;
    line_140_valid_reg <= 5'h15 == _io_out_T_2;
    line_141_valid_reg <= 5'h16 == _io_out_T_2;
    line_142_valid_reg <= 5'h17 == _io_out_T_2;
    line_143_valid_reg <= 5'h18 == _io_out_T_2;
    line_144_valid_reg <= 5'h19 == _io_out_T_2;
    line_145_valid_reg <= 5'h1a == _io_out_T_2;
    line_146_valid_reg <= 5'h1b == _io_out_T_2;
    line_147_valid_reg <= 5'h1c == _io_out_T_2;
    line_148_valid_reg <= 5'h1d == _io_out_T_2;
    line_149_valid_reg <= 5'h1e == _io_out_T_2;
    line_150_valid_reg <= 5'h1f == _io_out_T_2;
    line_151_valid_reg <= 5'h0 == _io_out_T_2;
    line_152_valid_reg <= 5'h1 == _io_out_T_2;
    line_153_valid_reg <= 5'h2 == _io_out_T_2;
    line_154_valid_reg <= 5'h3 == _io_out_T_2;
    line_155_valid_reg <= 5'h4 == _io_out_T_2;
    line_156_valid_reg <= 5'h5 == _io_out_T_2;
    line_157_valid_reg <= 5'h6 == _io_out_T_2;
    line_158_valid_reg <= 5'h7 == _io_out_T_2;
    line_159_valid_reg <= 5'h8 == _io_out_T_2;
    line_160_valid_reg <= 5'h9 == _io_out_T_2;
    line_161_valid_reg <= 5'ha == _io_out_T_2;
    line_162_valid_reg <= 5'hb == _io_out_T_2;
    line_163_valid_reg <= 5'hc == _io_out_T_2;
    line_164_valid_reg <= 5'hd == _io_out_T_2;
    line_165_valid_reg <= 5'he == _io_out_T_2;
    line_166_valid_reg <= 5'hf == _io_out_T_2;
    line_167_valid_reg <= 5'h10 == _io_out_T_2;
    line_168_valid_reg <= 5'h11 == _io_out_T_2;
    line_169_valid_reg <= 5'h12 == _io_out_T_2;
    line_170_valid_reg <= 5'h13 == _io_out_T_2;
    line_171_valid_reg <= 5'h14 == _io_out_T_2;
    line_172_valid_reg <= 5'h15 == _io_out_T_2;
    line_173_valid_reg <= 5'h16 == _io_out_T_2;
    line_174_valid_reg <= 5'h17 == _io_out_T_2;
    line_175_valid_reg <= 5'h18 == _io_out_T_2;
    line_176_valid_reg <= 5'h19 == _io_out_T_2;
    line_177_valid_reg <= 5'h1a == _io_out_T_2;
    line_178_valid_reg <= 5'h1b == _io_out_T_2;
    line_179_valid_reg <= 5'h1c == _io_out_T_2;
    line_180_valid_reg <= 5'h1d == _io_out_T_2;
    line_181_valid_reg <= 5'h1e == _io_out_T_2;
    line_182_valid_reg <= 5'h1f == _io_out_T_2;
    line_183_valid_reg <= 5'h0 == _io_out_T_2;
    line_184_valid_reg <= 5'h1 == _io_out_T_2;
    line_185_valid_reg <= 5'h2 == _io_out_T_2;
    line_186_valid_reg <= 5'h3 == _io_out_T_2;
    line_187_valid_reg <= 5'h4 == _io_out_T_2;
    line_188_valid_reg <= 5'h5 == _io_out_T_2;
    line_189_valid_reg <= 5'h6 == _io_out_T_2;
    line_190_valid_reg <= 5'h7 == _io_out_T_2;
    line_191_valid_reg <= 5'h8 == _io_out_T_2;
    line_192_valid_reg <= 5'h9 == _io_out_T_2;
    line_193_valid_reg <= 5'ha == _io_out_T_2;
    line_194_valid_reg <= 5'hb == _io_out_T_2;
    line_195_valid_reg <= 5'hc == _io_out_T_2;
    line_196_valid_reg <= 5'hd == _io_out_T_2;
    line_197_valid_reg <= 5'he == _io_out_T_2;
    line_198_valid_reg <= 5'hf == _io_out_T_2;
    line_199_valid_reg <= 5'h10 == _io_out_T_2;
    line_200_valid_reg <= 5'h11 == _io_out_T_2;
    line_201_valid_reg <= 5'h12 == _io_out_T_2;
    line_202_valid_reg <= 5'h13 == _io_out_T_2;
    line_203_valid_reg <= 5'h14 == _io_out_T_2;
    line_204_valid_reg <= 5'h15 == _io_out_T_2;
    line_205_valid_reg <= 5'h16 == _io_out_T_2;
    line_206_valid_reg <= 5'h17 == _io_out_T_2;
    line_207_valid_reg <= 5'h18 == _io_out_T_2;
    line_208_valid_reg <= 5'h19 == _io_out_T_2;
    line_209_valid_reg <= 5'h1a == _io_out_T_2;
    line_210_valid_reg <= 5'h1b == _io_out_T_2;
    line_211_valid_reg <= 5'h1c == _io_out_T_2;
    line_212_valid_reg <= 5'h1d == _io_out_T_2;
    line_213_valid_reg <= 5'h1e == _io_out_T_2;
    line_214_valid_reg <= 5'h1f == _io_out_T_2;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_43_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_44_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_45_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_46_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_47_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_48_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_49_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_50_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_51_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_52_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_53_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_54_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_55_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_56_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_57_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_58_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_59_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_60_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_61_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_62_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_63_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_64_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_65_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_66_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_67_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_68_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_69_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_70_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_71_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_72_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_73_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_74_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_75_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_76_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_77_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_78_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_79_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_80_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_81_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_82_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_83_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_84_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_85_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_86_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_87_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_88_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_89_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_90_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_91_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_92_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_93_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_94_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_95_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_96_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_97_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_98_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_99_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_100_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_101_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_102_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_103_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_104_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_105_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_106_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_107_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_108_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_109_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_110_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_111_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_112_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_113_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_114_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_115_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_116_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_117_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_118_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_119_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_120_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_121_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_122_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_123_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_124_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_125_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_126_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_127_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_128_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_129_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_130_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_131_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_132_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_133_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_134_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_135_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_136_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_137_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_138_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_139_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_140_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_141_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_142_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_143_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_144_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_145_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_146_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_147_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_148_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_149_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_150_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_151_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_152_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_153_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_154_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_155_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_156_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_157_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_158_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_159_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_160_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_161_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_162_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_163_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_164_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_165_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_166_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_167_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_168_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_169_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_170_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_171_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_172_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_173_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_174_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_175_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_176_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_177_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_178_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_179_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_180_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_181_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_182_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_183_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_184_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_185_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_186_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_187_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_188_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_189_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_190_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_191_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_192_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_193_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_194_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_195_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_196_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_197_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_198_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_199_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_200_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_201_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_202_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_203_valid_reg = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  line_204_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  line_205_valid_reg = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  line_206_valid_reg = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  line_207_valid_reg = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  line_208_valid_reg = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  line_209_valid_reg = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  line_210_valid_reg = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  line_211_valid_reg = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  line_212_valid_reg = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  line_213_valid_reg = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  line_214_valid_reg = _RAND_171[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (3'h0 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h1 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h2 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h3 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h4 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h5 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h6 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (3'h7 == _io_out_s_funct_T_2) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_in[11:10]) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_in[11:10]) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_in[11:10]) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_in[11:10]) begin
      cover(1'h1);
    end
    //
    if (5'h0 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'ha == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hb == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hc == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hd == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'he == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hf == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h0 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'ha == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hb == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hc == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hd == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'he == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hf == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h0 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'ha == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hb == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hc == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hd == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'he == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hf == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h0 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'ha == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hb == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hc == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hd == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'he == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hf == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h0 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'ha == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hb == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hc == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hd == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'he == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'hf == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == _io_out_T_2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == _io_out_T_2) begin
      cover(1'h1);
    end
  end
endmodule
module Decoder(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_isWFI, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  expander_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire  expander_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] expander_io_in; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] expander_io_out_bits; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] _decodeList_T = expander_io_out_bits & 32'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_1 = 32'h13 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_2 = expander_io_out_bits & 32'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_3 = 32'h1013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_5 = 32'h2013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_7 = 32'h3013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_9 = 32'h4013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_11 = 32'h5013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_13 = 32'h6013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_15 = 32'h7013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_17 = 32'h40005013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_18 = expander_io_out_bits & 32'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_19 = 32'h33 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_21 = 32'h1033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_23 = 32'h2033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_25 = 32'h3033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_27 = 32'h4033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_29 = 32'h5033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_31 = 32'h6033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_33 = 32'h7033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_35 = 32'h40000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_37 = 32'h40005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_38 = expander_io_out_bits & 32'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_39 = 32'h17 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_41 = 32'h37 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_43 = 32'h6f == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_45 = 32'h67 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_47 = 32'h63 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_49 = 32'h1063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_51 = 32'h4063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_53 = 32'h5063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_55 = 32'h6063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_57 = 32'h7063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_59 = 32'h3 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_61 = 32'h1003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_63 = 32'h2003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_65 = 32'h4003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_67 = 32'h5003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_69 = 32'h23 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_71 = 32'h1023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_73 = 32'h2023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_75 = 32'h1b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_77 = 32'h101b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_79 = 32'h501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_81 = 32'h4000501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_83 = 32'h103b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_85 = 32'h503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_87 = 32'h4000503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_89 = 32'h3b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_91 = 32'h4000003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_93 = 32'h6003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_95 = 32'h3003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_97 = 32'h3023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_99 = 32'h6b == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_101 = 32'h2000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_103 = 32'h2001033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_105 = 32'h2002033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_107 = 32'h2003033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_109 = 32'h2004033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_111 = 32'h2005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_113 = 32'h2006033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_115 = 32'h2007033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_117 = 32'h200003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_119 = 32'h200403b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_121 = 32'h200503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_123 = 32'h200603b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_125 = 32'h200703b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_126 = expander_io_out_bits; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_127 = 32'h73 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_129 = 32'h100073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_131 = 32'h30200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_133 = 32'hf == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_135 = 32'h10500073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_137 = 32'h10200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_138 = expander_io_out_bits & 32'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_139 = 32'h12000073 == _decodeList_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_140 = expander_io_out_bits & 32'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_141 = 32'h1000302f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_143 = 32'h1000202f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_144 = expander_io_out_bits & 32'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_145 = 32'h1800302f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_147 = 32'h1800202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_148 = expander_io_out_bits & 32'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_149 = 32'h800202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_151 = 32'h202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_153 = 32'h2000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_155 = 32'h6000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_157 = 32'h4000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_159 = 32'h8000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_161 = 32'ha000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_163 = 32'hc000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_165 = 32'he000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_167 = 32'h1073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_169 = 32'h2073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_171 = 32'h3073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_173 = 32'h5073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_175 = 32'h6073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_177 = 32'h7073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_179 = 32'h100f == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _decodeList_T_181 = _decodeList_T_177 ? 3'h4 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_182 = _decodeList_T_175 ? 3'h4 : _decodeList_T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_183 = _decodeList_T_173 ? 3'h4 : _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_184 = _decodeList_T_171 ? 3'h4 : _decodeList_T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_185 = _decodeList_T_169 ? 3'h4 : _decodeList_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_186 = _decodeList_T_167 ? 3'h4 : _decodeList_T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_187 = _decodeList_T_165 ? 3'h5 : _decodeList_T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_188 = _decodeList_T_163 ? 3'h5 : _decodeList_T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_189 = _decodeList_T_161 ? 3'h5 : _decodeList_T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_190 = _decodeList_T_159 ? 3'h5 : _decodeList_T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_191 = _decodeList_T_157 ? 3'h5 : _decodeList_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_192 = _decodeList_T_155 ? 3'h5 : _decodeList_T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_193 = _decodeList_T_153 ? 3'h5 : _decodeList_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_194 = _decodeList_T_151 ? 3'h5 : _decodeList_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_195 = _decodeList_T_149 ? 3'h5 : _decodeList_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_196 = _decodeList_T_147 ? 4'hf : {{1'd0}, _decodeList_T_195}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_197 = _decodeList_T_145 ? 4'hf : _decodeList_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_198 = _decodeList_T_143 ? 4'h5 : _decodeList_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_199 = _decodeList_T_141 ? 4'h5 : _decodeList_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_200 = _decodeList_T_139 ? 4'h5 : _decodeList_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_201 = _decodeList_T_137 ? 4'h4 : _decodeList_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_202 = _decodeList_T_135 ? 4'h4 : _decodeList_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_203 = _decodeList_T_133 ? 4'h2 : _decodeList_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_204 = _decodeList_T_131 ? 4'h4 : _decodeList_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_205 = _decodeList_T_129 ? 4'h4 : _decodeList_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_206 = _decodeList_T_127 ? 4'h4 : _decodeList_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_207 = _decodeList_T_125 ? 4'h5 : _decodeList_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_208 = _decodeList_T_123 ? 4'h5 : _decodeList_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_209 = _decodeList_T_121 ? 4'h5 : _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_210 = _decodeList_T_119 ? 4'h5 : _decodeList_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_211 = _decodeList_T_117 ? 4'h5 : _decodeList_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_212 = _decodeList_T_115 ? 4'h5 : _decodeList_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_213 = _decodeList_T_113 ? 4'h5 : _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_214 = _decodeList_T_111 ? 4'h5 : _decodeList_T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_215 = _decodeList_T_109 ? 4'h5 : _decodeList_T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_216 = _decodeList_T_107 ? 4'h5 : _decodeList_T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_217 = _decodeList_T_105 ? 4'h5 : _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_218 = _decodeList_T_103 ? 4'h5 : _decodeList_T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_219 = _decodeList_T_101 ? 4'h5 : _decodeList_T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_220 = _decodeList_T_99 ? 4'h4 : _decodeList_T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_221 = _decodeList_T_97 ? 4'h2 : _decodeList_T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_222 = _decodeList_T_95 ? 4'h4 : _decodeList_T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_223 = _decodeList_T_93 ? 4'h4 : _decodeList_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_224 = _decodeList_T_91 ? 4'h5 : _decodeList_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_225 = _decodeList_T_89 ? 4'h5 : _decodeList_T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_226 = _decodeList_T_87 ? 4'h5 : _decodeList_T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_227 = _decodeList_T_85 ? 4'h5 : _decodeList_T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_228 = _decodeList_T_83 ? 4'h5 : _decodeList_T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_229 = _decodeList_T_81 ? 4'h4 : _decodeList_T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_230 = _decodeList_T_79 ? 4'h4 : _decodeList_T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_231 = _decodeList_T_77 ? 4'h4 : _decodeList_T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_232 = _decodeList_T_75 ? 4'h4 : _decodeList_T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_233 = _decodeList_T_73 ? 4'h2 : _decodeList_T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_234 = _decodeList_T_71 ? 4'h2 : _decodeList_T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_235 = _decodeList_T_69 ? 4'h2 : _decodeList_T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_236 = _decodeList_T_67 ? 4'h4 : _decodeList_T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_237 = _decodeList_T_65 ? 4'h4 : _decodeList_T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_238 = _decodeList_T_63 ? 4'h4 : _decodeList_T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_239 = _decodeList_T_61 ? 4'h4 : _decodeList_T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_240 = _decodeList_T_59 ? 4'h4 : _decodeList_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_241 = _decodeList_T_57 ? 4'h1 : _decodeList_T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_242 = _decodeList_T_55 ? 4'h1 : _decodeList_T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_243 = _decodeList_T_53 ? 4'h1 : _decodeList_T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_244 = _decodeList_T_51 ? 4'h1 : _decodeList_T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_245 = _decodeList_T_49 ? 4'h1 : _decodeList_T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_246 = _decodeList_T_47 ? 4'h1 : _decodeList_T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_247 = _decodeList_T_45 ? 4'h4 : _decodeList_T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_248 = _decodeList_T_43 ? 4'h7 : _decodeList_T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_249 = _decodeList_T_41 ? 4'h6 : _decodeList_T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_250 = _decodeList_T_39 ? 4'h6 : _decodeList_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_251 = _decodeList_T_37 ? 4'h5 : _decodeList_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_252 = _decodeList_T_35 ? 4'h5 : _decodeList_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_253 = _decodeList_T_33 ? 4'h5 : _decodeList_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_254 = _decodeList_T_31 ? 4'h5 : _decodeList_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_255 = _decodeList_T_29 ? 4'h5 : _decodeList_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_256 = _decodeList_T_27 ? 4'h5 : _decodeList_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_257 = _decodeList_T_25 ? 4'h5 : _decodeList_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_258 = _decodeList_T_23 ? 4'h5 : _decodeList_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_259 = _decodeList_T_21 ? 4'h5 : _decodeList_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_260 = _decodeList_T_19 ? 4'h5 : _decodeList_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_261 = _decodeList_T_17 ? 4'h4 : _decodeList_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_262 = _decodeList_T_15 ? 4'h4 : _decodeList_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_263 = _decodeList_T_13 ? 4'h4 : _decodeList_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_264 = _decodeList_T_11 ? 4'h4 : _decodeList_T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_265 = _decodeList_T_9 ? 4'h4 : _decodeList_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_266 = _decodeList_T_7 ? 4'h4 : _decodeList_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_267 = _decodeList_T_5 ? 4'h4 : _decodeList_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_268 = _decodeList_T_3 ? 4'h4 : _decodeList_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] decodeList_0 = _decodeList_T_1 ? 4'h4 : _decodeList_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_269 = _decodeList_T_179 ? 3'h4 : 3'h3; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_270 = _decodeList_T_177 ? 3'h3 : _decodeList_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_271 = _decodeList_T_175 ? 3'h3 : _decodeList_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_272 = _decodeList_T_173 ? 3'h3 : _decodeList_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_273 = _decodeList_T_171 ? 3'h3 : _decodeList_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_274 = _decodeList_T_169 ? 3'h3 : _decodeList_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_275 = _decodeList_T_167 ? 3'h3 : _decodeList_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_276 = _decodeList_T_165 ? 3'h1 : _decodeList_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_277 = _decodeList_T_163 ? 3'h1 : _decodeList_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_278 = _decodeList_T_161 ? 3'h1 : _decodeList_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_279 = _decodeList_T_159 ? 3'h1 : _decodeList_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_280 = _decodeList_T_157 ? 3'h1 : _decodeList_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_281 = _decodeList_T_155 ? 3'h1 : _decodeList_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_282 = _decodeList_T_153 ? 3'h1 : _decodeList_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_283 = _decodeList_T_151 ? 3'h1 : _decodeList_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_284 = _decodeList_T_149 ? 3'h1 : _decodeList_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_285 = _decodeList_T_147 ? 3'h1 : _decodeList_T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_286 = _decodeList_T_145 ? 3'h1 : _decodeList_T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_287 = _decodeList_T_143 ? 3'h1 : _decodeList_T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_288 = _decodeList_T_141 ? 3'h1 : _decodeList_T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_289 = _decodeList_T_139 ? 3'h4 : _decodeList_T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_290 = _decodeList_T_137 ? 3'h3 : _decodeList_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_291 = _decodeList_T_135 ? 3'h0 : _decodeList_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_292 = _decodeList_T_133 ? 3'h4 : _decodeList_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_293 = _decodeList_T_131 ? 3'h3 : _decodeList_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_294 = _decodeList_T_129 ? 3'h3 : _decodeList_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_295 = _decodeList_T_127 ? 3'h3 : _decodeList_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_296 = _decodeList_T_125 ? 3'h2 : _decodeList_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_297 = _decodeList_T_123 ? 3'h2 : _decodeList_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_298 = _decodeList_T_121 ? 3'h2 : _decodeList_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_299 = _decodeList_T_119 ? 3'h2 : _decodeList_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_300 = _decodeList_T_117 ? 3'h2 : _decodeList_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_301 = _decodeList_T_115 ? 3'h2 : _decodeList_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_302 = _decodeList_T_113 ? 3'h2 : _decodeList_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_303 = _decodeList_T_111 ? 3'h2 : _decodeList_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_304 = _decodeList_T_109 ? 3'h2 : _decodeList_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_305 = _decodeList_T_107 ? 3'h2 : _decodeList_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_306 = _decodeList_T_105 ? 3'h2 : _decodeList_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_307 = _decodeList_T_103 ? 3'h2 : _decodeList_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_308 = _decodeList_T_101 ? 3'h2 : _decodeList_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_309 = _decodeList_T_99 ? 3'h3 : _decodeList_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_310 = _decodeList_T_97 ? 3'h1 : _decodeList_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_311 = _decodeList_T_95 ? 3'h1 : _decodeList_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_312 = _decodeList_T_93 ? 3'h1 : _decodeList_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_313 = _decodeList_T_91 ? 3'h0 : _decodeList_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_314 = _decodeList_T_89 ? 3'h0 : _decodeList_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_315 = _decodeList_T_87 ? 3'h0 : _decodeList_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_316 = _decodeList_T_85 ? 3'h0 : _decodeList_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_317 = _decodeList_T_83 ? 3'h0 : _decodeList_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_318 = _decodeList_T_81 ? 3'h0 : _decodeList_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_319 = _decodeList_T_79 ? 3'h0 : _decodeList_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_320 = _decodeList_T_77 ? 3'h0 : _decodeList_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_321 = _decodeList_T_75 ? 3'h0 : _decodeList_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_322 = _decodeList_T_73 ? 3'h1 : _decodeList_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_323 = _decodeList_T_71 ? 3'h1 : _decodeList_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_324 = _decodeList_T_69 ? 3'h1 : _decodeList_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_325 = _decodeList_T_67 ? 3'h1 : _decodeList_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_326 = _decodeList_T_65 ? 3'h1 : _decodeList_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_327 = _decodeList_T_63 ? 3'h1 : _decodeList_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_328 = _decodeList_T_61 ? 3'h1 : _decodeList_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_329 = _decodeList_T_59 ? 3'h1 : _decodeList_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_330 = _decodeList_T_57 ? 3'h0 : _decodeList_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_331 = _decodeList_T_55 ? 3'h0 : _decodeList_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_332 = _decodeList_T_53 ? 3'h0 : _decodeList_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_333 = _decodeList_T_51 ? 3'h0 : _decodeList_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_334 = _decodeList_T_49 ? 3'h0 : _decodeList_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_335 = _decodeList_T_47 ? 3'h0 : _decodeList_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_336 = _decodeList_T_45 ? 3'h0 : _decodeList_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_337 = _decodeList_T_43 ? 3'h0 : _decodeList_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_338 = _decodeList_T_41 ? 3'h0 : _decodeList_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_339 = _decodeList_T_39 ? 3'h0 : _decodeList_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_340 = _decodeList_T_37 ? 3'h0 : _decodeList_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_341 = _decodeList_T_35 ? 3'h0 : _decodeList_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_342 = _decodeList_T_33 ? 3'h0 : _decodeList_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_343 = _decodeList_T_31 ? 3'h0 : _decodeList_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_344 = _decodeList_T_29 ? 3'h0 : _decodeList_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_345 = _decodeList_T_27 ? 3'h0 : _decodeList_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_346 = _decodeList_T_25 ? 3'h0 : _decodeList_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_347 = _decodeList_T_23 ? 3'h0 : _decodeList_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_348 = _decodeList_T_21 ? 3'h0 : _decodeList_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_349 = _decodeList_T_19 ? 3'h0 : _decodeList_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_350 = _decodeList_T_17 ? 3'h0 : _decodeList_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_351 = _decodeList_T_15 ? 3'h0 : _decodeList_T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_352 = _decodeList_T_13 ? 3'h0 : _decodeList_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_353 = _decodeList_T_11 ? 3'h0 : _decodeList_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_354 = _decodeList_T_9 ? 3'h0 : _decodeList_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_355 = _decodeList_T_7 ? 3'h0 : _decodeList_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_356 = _decodeList_T_5 ? 3'h0 : _decodeList_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_357 = _decodeList_T_3 ? 3'h0 : _decodeList_T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] decodeList_1 = _decodeList_T_1 ? 3'h0 : _decodeList_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_359 = _decodeList_T_177 ? 3'h7 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_360 = _decodeList_T_175 ? 3'h6 : _decodeList_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_361 = _decodeList_T_173 ? 3'h5 : _decodeList_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_362 = _decodeList_T_171 ? 3'h3 : _decodeList_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_363 = _decodeList_T_169 ? 3'h2 : _decodeList_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_364 = _decodeList_T_167 ? 3'h1 : _decodeList_T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_365 = _decodeList_T_165 ? 6'h32 : {{3'd0}, _decodeList_T_364}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_366 = _decodeList_T_163 ? 6'h31 : _decodeList_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_367 = _decodeList_T_161 ? 6'h30 : _decodeList_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_368 = _decodeList_T_159 ? 6'h37 : _decodeList_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_369 = _decodeList_T_157 ? 6'h26 : _decodeList_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_370 = _decodeList_T_155 ? 6'h25 : _decodeList_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_371 = _decodeList_T_153 ? 6'h24 : _decodeList_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_372 = _decodeList_T_151 ? 7'h63 : {{1'd0}, _decodeList_T_371}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_373 = _decodeList_T_149 ? 7'h22 : _decodeList_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_374 = _decodeList_T_147 ? 7'h21 : _decodeList_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_375 = _decodeList_T_145 ? 7'h21 : _decodeList_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_376 = _decodeList_T_143 ? 7'h20 : _decodeList_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_377 = _decodeList_T_141 ? 7'h20 : _decodeList_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_378 = _decodeList_T_139 ? 7'h2 : _decodeList_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_379 = _decodeList_T_137 ? 7'h0 : _decodeList_T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_380 = _decodeList_T_135 ? 7'h40 : _decodeList_T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_381 = _decodeList_T_133 ? 7'h0 : _decodeList_T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_382 = _decodeList_T_131 ? 7'h0 : _decodeList_T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_383 = _decodeList_T_129 ? 7'h0 : _decodeList_T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_384 = _decodeList_T_127 ? 7'h0 : _decodeList_T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_385 = _decodeList_T_125 ? 7'hf : _decodeList_T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_386 = _decodeList_T_123 ? 7'he : _decodeList_T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_387 = _decodeList_T_121 ? 7'hd : _decodeList_T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_388 = _decodeList_T_119 ? 7'hc : _decodeList_T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_389 = _decodeList_T_117 ? 7'h8 : _decodeList_T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_390 = _decodeList_T_115 ? 7'h7 : _decodeList_T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_391 = _decodeList_T_113 ? 7'h6 : _decodeList_T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_392 = _decodeList_T_111 ? 7'h5 : _decodeList_T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_393 = _decodeList_T_109 ? 7'h4 : _decodeList_T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_394 = _decodeList_T_107 ? 7'h3 : _decodeList_T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_395 = _decodeList_T_105 ? 7'h2 : _decodeList_T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_396 = _decodeList_T_103 ? 7'h1 : _decodeList_T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_397 = _decodeList_T_101 ? 7'h0 : _decodeList_T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_398 = _decodeList_T_99 ? 7'h2 : _decodeList_T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_399 = _decodeList_T_97 ? 7'hb : _decodeList_T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_400 = _decodeList_T_95 ? 7'h3 : _decodeList_T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_401 = _decodeList_T_93 ? 7'h6 : _decodeList_T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_402 = _decodeList_T_91 ? 7'h28 : _decodeList_T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_403 = _decodeList_T_89 ? 7'h60 : _decodeList_T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_404 = _decodeList_T_87 ? 7'h2d : _decodeList_T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_405 = _decodeList_T_85 ? 7'h25 : _decodeList_T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_406 = _decodeList_T_83 ? 7'h21 : _decodeList_T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_407 = _decodeList_T_81 ? 7'h2d : _decodeList_T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_408 = _decodeList_T_79 ? 7'h25 : _decodeList_T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_409 = _decodeList_T_77 ? 7'h21 : _decodeList_T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_410 = _decodeList_T_75 ? 7'h60 : _decodeList_T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_411 = _decodeList_T_73 ? 7'ha : _decodeList_T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_412 = _decodeList_T_71 ? 7'h9 : _decodeList_T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_413 = _decodeList_T_69 ? 7'h8 : _decodeList_T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_414 = _decodeList_T_67 ? 7'h5 : _decodeList_T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_415 = _decodeList_T_65 ? 7'h4 : _decodeList_T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_416 = _decodeList_T_63 ? 7'h2 : _decodeList_T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_417 = _decodeList_T_61 ? 7'h1 : _decodeList_T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_418 = _decodeList_T_59 ? 7'h0 : _decodeList_T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_419 = _decodeList_T_57 ? 7'h17 : _decodeList_T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_420 = _decodeList_T_55 ? 7'h16 : _decodeList_T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_421 = _decodeList_T_53 ? 7'h15 : _decodeList_T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_422 = _decodeList_T_51 ? 7'h14 : _decodeList_T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_423 = _decodeList_T_49 ? 7'h11 : _decodeList_T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_424 = _decodeList_T_47 ? 7'h10 : _decodeList_T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_425 = _decodeList_T_45 ? 7'h5a : _decodeList_T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_426 = _decodeList_T_43 ? 7'h58 : _decodeList_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_427 = _decodeList_T_41 ? 7'h40 : _decodeList_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_428 = _decodeList_T_39 ? 7'h40 : _decodeList_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_429 = _decodeList_T_37 ? 7'hd : _decodeList_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_430 = _decodeList_T_35 ? 7'h8 : _decodeList_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_431 = _decodeList_T_33 ? 7'h7 : _decodeList_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_432 = _decodeList_T_31 ? 7'h6 : _decodeList_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_433 = _decodeList_T_29 ? 7'h5 : _decodeList_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_434 = _decodeList_T_27 ? 7'h4 : _decodeList_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_435 = _decodeList_T_25 ? 7'h3 : _decodeList_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_436 = _decodeList_T_23 ? 7'h2 : _decodeList_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_437 = _decodeList_T_21 ? 7'h1 : _decodeList_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_438 = _decodeList_T_19 ? 7'h40 : _decodeList_T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_439 = _decodeList_T_17 ? 7'hd : _decodeList_T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_440 = _decodeList_T_15 ? 7'h7 : _decodeList_T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_441 = _decodeList_T_13 ? 7'h6 : _decodeList_T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_442 = _decodeList_T_11 ? 7'h5 : _decodeList_T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_443 = _decodeList_T_9 ? 7'h4 : _decodeList_T_442; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_444 = _decodeList_T_7 ? 7'h3 : _decodeList_T_443; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_445 = _decodeList_T_5 ? 7'h2 : _decodeList_T_444; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_446 = _decodeList_T_3 ? 7'h1 : _decodeList_T_445; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] decodeList_2 = _decodeList_T_1 ? 7'h40 : _decodeList_T_446; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  hasIntr = |intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 130:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire  _src1Type_T = 4'h4 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = expander_io_out_bits[19:15]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:28]
  wire [4:0] rt = expander_io_out_bits[24:20]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:43]
  wire [4:0] rd = expander_io_out_bits[11:7]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:58]
  wire  imm_signBit = expander_io_out_bits[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_1 = imm_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_2 = {_imm_T_1,expander_io_out_bits[31:20]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [11:0] _imm_T_5 = {expander_io_out_bits[31:25],rd}; // @[src/main/scala/nutcore/frontend/IDU.scala 82:27]
  wire  imm_signBit_1 = _imm_T_5[11]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_6 = imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_7 = {_imm_T_6,expander_io_out_bits[31:25],rd}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [12:0] _imm_T_17 = {expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 84:27]
  wire  imm_signBit_3 = _imm_T_17[12]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [50:0] _imm_T_18 = imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_19 = {_imm_T_18,expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [31:0] _imm_T_21 = {expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 85:27]
  wire  imm_signBit_4 = _imm_T_21[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _imm_T_22 = imm_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_23 = {_imm_T_22,expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [20:0] _imm_T_28 = {expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 86:27]
  wire  imm_signBit_5 = _imm_T_28[20]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [42:0] _imm_T_29 = imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_30 = {_imm_T_29,expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imm_T_37 = _src1Type_T ? _imm_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_38 = _src1Type_T_2 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_39 = _src1Type_T_3 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_40 = _src1Type_T_4 ? _imm_T_19 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_41 = _src1Type_T_5 ? _imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_42 = _src1Type_T_6 ? _imm_T_30 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_43 = _imm_T_37 | _imm_T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_44 = _imm_T_43 | _imm_T_39; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_45 = _imm_T_44 | _imm_T_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_46 = _imm_T_45 | _imm_T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_6 = fuType == 3'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 90:16]
  wire  line_215_clock;
  wire  line_215_reset;
  wire  line_215_valid;
  reg  line_215_valid_reg;
  wire  _T_9 = rd == 5'h1 | rd == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire  _T_11 = _T_9 & fuOpType == 7'h58; // @[src/main/scala/nutcore/frontend/IDU.scala 92:26]
  wire  line_216_clock;
  wire  line_216_reset;
  wire  line_216_valid;
  reg  line_216_valid_reg;
  wire [6:0] _GEN_5 = _T_9 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 92:{57,85}]
  wire  _T_12 = fuOpType == 7'h5a; // @[src/main/scala/nutcore/frontend/IDU.scala 93:20]
  wire  line_217_clock;
  wire  line_217_reset;
  wire  line_217_valid;
  reg  line_217_valid_reg;
  wire  _T_15 = rs == 5'h1 | rs == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire  line_218_clock;
  wire  line_218_reset;
  wire  line_218_valid;
  reg  line_218_valid_reg;
  wire [6:0] _GEN_6 = _T_15 ? 7'h5e : _GEN_5; // @[src/main/scala/nutcore/frontend/IDU.scala 94:{29,57}]
  wire  line_219_clock;
  wire  line_219_reset;
  wire  line_219_valid;
  reg  line_219_valid_reg;
  wire [6:0] _GEN_7 = _T_9 ? 7'h5c : _GEN_6; // @[src/main/scala/nutcore/frontend/IDU.scala 95:{29,57}]
  wire [6:0] _GEN_8 = fuOpType == 7'h5a ? _GEN_7 : _GEN_5; // @[src/main/scala/nutcore/frontend/IDU.scala 93:40]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  is_sfence_vma = fuType == 3'h4 & fuOpType == 7'h2; // @[src/main/scala/nutcore/frontend/IDU.scala 136:45]
  wire  sfence_vma_illegal = is_sfence_vma & io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 137:42]
  wire  wfi_illegal = io_isWFI & io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 138:30]
  wire  illegal_instr = instrType == 4'h0 | sfence_vma_illegal | wfi_illegal; // @[src/main/scala/nutcore/frontend/IDU.scala 139:82]
  RVCExpander expander ( // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
    .clock(expander_clock),
    .reset(expander_reset),
    .io_in(expander_io_in),
    .io_out_bits(expander_io_out_bits)
  );
  GEN_w1_line #(.COVER_INDEX(215)) line_215 (
    .clock(line_215_clock),
    .reset(line_215_reset),
    .valid(line_215_valid)
  );
  GEN_w1_line #(.COVER_INDEX(216)) line_216 (
    .clock(line_216_clock),
    .reset(line_216_reset),
    .valid(line_216_valid)
  );
  GEN_w1_line #(.COVER_INDEX(217)) line_217 (
    .clock(line_217_clock),
    .reset(line_217_reset),
    .valid(line_217_valid)
  );
  GEN_w1_line #(.COVER_INDEX(218)) line_218 (
    .clock(line_218_clock),
    .reset(line_218_reset),
    .valid(line_218_valid)
  );
  GEN_w1_line #(.COVER_INDEX(219)) line_219 (
    .clock(line_219_clock),
    .reset(line_219_reset),
    .valid(line_219_valid)
  );
  assign line_215_clock = clock;
  assign line_215_reset = reset;
  assign line_215_valid = _T_6 ^ line_215_valid_reg;
  assign line_216_clock = clock;
  assign line_216_reset = reset;
  assign line_216_valid = _T_11 ^ line_216_valid_reg;
  assign line_217_clock = clock;
  assign line_217_reset = reset;
  assign line_217_valid = _T_12 ^ line_217_valid_reg;
  assign line_218_clock = clock;
  assign line_218_reset = reset;
  assign line_218_valid = _T_15 ^ line_218_valid_reg;
  assign line_219_clock = clock;
  assign line_219_reset = reset;
  assign line_219_valid = _T_9 ^ line_219_valid_reg;
  assign io_in_ready = ~io_in_valid | _io_in_ready_T_1; // @[src/main/scala/nutcore/frontend/IDU.scala 120:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 119:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 142:49]
  assign io_out_bits_cf_exceptionVec_2 = illegal_instr & ~hasIntr & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 140:74]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 141:47]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_ctrl_src1Type = expander_io_out_bits[6:0] == 7'h37 ? 1'h0 : src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 99:35]
  assign io_out_bits_ctrl_src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_8 : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 90:32]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rs; // @[src/main/scala/nutcore/frontend/IDU.scala 74:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rt : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 75:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[src/main/scala/nutcore/Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rd : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 77:33]
  assign io_out_bits_ctrl_isNutCoreTrap = _decodeList_T_99 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 144:66]
  assign io_out_bits_data_imm = _imm_T_46 | _imm_T_42; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_isWFI = _decodeList_T_135 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 145:43]
  assign expander_clock = clock;
  assign expander_reset = reset;
  assign expander_io_in = io_in_bits_instr[31:0]; // @[src/main/scala/nutcore/frontend/IDU.scala 36:18]
  always @(posedge clock) begin
    line_215_valid_reg <= _T_6;
    line_216_valid_reg <= _T_11;
    line_217_valid_reg <= _T_12;
    line_218_valid_reg <= _T_15;
    line_219_valid_reg <= _T_9;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_215_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_216_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_217_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_218_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_219_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_6) begin
      cover(1'h1);
    end
    //
    if (_T_6 & _T_11) begin
      cover(1'h1);
    end
    //
    if (_T_6 & _T_12) begin
      cover(1'h1);
    end
    //
    if (_T_6 & _T_12 & _T_15) begin
      cover(1'h1);
    end
    //
    if (_T_6 & _T_12 & _T_9) begin
      cover(1'h1);
    end
  end
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [63:0] io_in_0_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [3:0]  io_in_0_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        isWFI_0,
  input  [11:0] intrVecIDU
);
  wire  decoder_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [2:0] decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [6:0] decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [11:0] decoder_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  isWFI = decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 175:{23,23}]
  Decoder decoder ( // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
    .clock(decoder_clock),
    .reset(decoder_reset),
    .io_in_ready(decoder_io_in_ready),
    .io_in_valid(decoder_io_in_valid),
    .io_in_bits_instr(decoder_io_in_bits_instr),
    .io_in_bits_pc(decoder_io_in_bits_pc),
    .io_in_bits_pnpc(decoder_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_1(decoder_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_12(decoder_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder_io_in_bits_brIdx),
    .io_in_bits_crossBoundaryFault(decoder_io_in_bits_crossBoundaryFault),
    .io_out_ready(decoder_io_out_ready),
    .io_out_valid(decoder_io_out_valid),
    .io_out_bits_cf_instr(decoder_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(decoder_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(decoder_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(decoder_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(decoder_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(decoder_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(decoder_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(decoder_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_src1Type(decoder_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(decoder_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_imm(decoder_io_out_bits_data_imm),
    .io_isWFI(decoder_io_isWFI),
    .io_sfence_vma_invalid(decoder_io_sfence_vma_invalid),
    .io_wfi_invalid(decoder_io_wfi_invalid),
    .intrVecIDU(decoder_intrVecIDU)
  );
  assign io_in_0_ready = decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign io_out_0_valid = decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_instr = decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pc = decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pnpc = decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_brIdx = decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_crossBoundaryFault = decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src1Type = decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src2Type = decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuType = decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfWen = decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfDest = decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_isNutCoreTrap = decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_data_imm = decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign isWFI_0 = isWFI;
  assign decoder_clock = clock;
  assign decoder_reset = reset;
  assign decoder_io_in_valid = io_in_0_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_instr = io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pc = io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_1 = io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_crossBoundaryFault = io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_out_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign decoder_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 171:33]
  assign decoder_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 172:26]
  assign decoder_intrVecIDU = intrVecIDU;
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [63:0] io_enq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [3:0]  io_enq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_deq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [63:0] io_deq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_0, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_2, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_3, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_4, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_5, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_6, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_7, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_8, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_9, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_10, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_11, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_12, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_13, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_14, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_15, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [3:0]  io_deq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_flush // @[src/main/scala/utils/FlushableQueue.scala 21:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pnpc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_0 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_1 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_2 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_3 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_4 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_5 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_6 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_7 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_8 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_9 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_10 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_11 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_12 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_13 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_14 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_15 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [3:0] ram_brIdx [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/utils/FlushableQueue.scala 28:41]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 29:33]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 30:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_220_clock;
  wire  line_220_reset;
  wire  line_220_valid;
  reg  line_220_valid_reg;
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_221_clock;
  wire  line_221_reset;
  wire  line_221_valid;
  reg  line_221_valid_reg;
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T = do_enq != do_deq; // @[src/main/scala/utils/FlushableQueue.scala 41:16]
  wire  line_222_clock;
  wire  line_222_reset;
  wire  line_222_valid;
  reg  line_222_valid_reg;
  wire  line_223_clock;
  wire  line_223_reset;
  wire  line_223_valid;
  reg  line_223_valid_reg;
  GEN_w1_line #(.COVER_INDEX(220)) line_220 (
    .clock(line_220_clock),
    .reset(line_220_reset),
    .valid(line_220_valid)
  );
  GEN_w1_line #(.COVER_INDEX(221)) line_221 (
    .clock(line_221_clock),
    .reset(line_221_reset),
    .valid(line_221_valid)
  );
  GEN_w1_line #(.COVER_INDEX(222)) line_222 (
    .clock(line_222_clock),
    .reset(line_222_reset),
    .valid(line_222_valid)
  );
  GEN_w1_line #(.COVER_INDEX(223)) line_223 (
    .clock(line_223_clock),
    .reset(line_223_reset),
    .valid(line_223_valid)
  );
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pnpc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pnpc_io_deq_bits_MPORT_data = ram_pnpc[ram_pnpc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign ram_pnpc_MPORT_addr = enq_ptr_value;
  assign ram_pnpc_MPORT_mask = 1'h1;
  assign ram_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_data = ram_exceptionVec_0[ram_exceptionVec_0_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_0_MPORT_data = 1'h0;
  assign ram_exceptionVec_0_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_0_MPORT_mask = 1'h1;
  assign ram_exceptionVec_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_data = ram_exceptionVec_1[ram_exceptionVec_1_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_1_MPORT_data = io_enq_bits_exceptionVec_1;
  assign ram_exceptionVec_1_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_1_MPORT_mask = 1'h1;
  assign ram_exceptionVec_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_data = ram_exceptionVec_2[ram_exceptionVec_2_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_2_MPORT_data = 1'h0;
  assign ram_exceptionVec_2_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_2_MPORT_mask = 1'h1;
  assign ram_exceptionVec_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_data = ram_exceptionVec_3[ram_exceptionVec_3_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_3_MPORT_data = 1'h0;
  assign ram_exceptionVec_3_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_3_MPORT_mask = 1'h1;
  assign ram_exceptionVec_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_data = ram_exceptionVec_4[ram_exceptionVec_4_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_4_MPORT_data = 1'h0;
  assign ram_exceptionVec_4_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_4_MPORT_mask = 1'h1;
  assign ram_exceptionVec_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_data = ram_exceptionVec_5[ram_exceptionVec_5_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_5_MPORT_data = 1'h0;
  assign ram_exceptionVec_5_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_5_MPORT_mask = 1'h1;
  assign ram_exceptionVec_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_data = ram_exceptionVec_6[ram_exceptionVec_6_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_6_MPORT_data = 1'h0;
  assign ram_exceptionVec_6_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_6_MPORT_mask = 1'h1;
  assign ram_exceptionVec_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_data = ram_exceptionVec_7[ram_exceptionVec_7_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_7_MPORT_data = 1'h0;
  assign ram_exceptionVec_7_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_7_MPORT_mask = 1'h1;
  assign ram_exceptionVec_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_data = ram_exceptionVec_8[ram_exceptionVec_8_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_8_MPORT_data = 1'h0;
  assign ram_exceptionVec_8_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_8_MPORT_mask = 1'h1;
  assign ram_exceptionVec_8_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_data = ram_exceptionVec_9[ram_exceptionVec_9_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_9_MPORT_data = 1'h0;
  assign ram_exceptionVec_9_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_9_MPORT_mask = 1'h1;
  assign ram_exceptionVec_9_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_data = ram_exceptionVec_10[ram_exceptionVec_10_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_10_MPORT_data = 1'h0;
  assign ram_exceptionVec_10_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_10_MPORT_mask = 1'h1;
  assign ram_exceptionVec_10_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_data = ram_exceptionVec_11[ram_exceptionVec_11_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_11_MPORT_data = 1'h0;
  assign ram_exceptionVec_11_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_11_MPORT_mask = 1'h1;
  assign ram_exceptionVec_11_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_data = ram_exceptionVec_12[ram_exceptionVec_12_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_12_MPORT_data = 1'h0;
  assign ram_exceptionVec_12_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_12_MPORT_mask = 1'h1;
  assign ram_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_data = ram_exceptionVec_13[ram_exceptionVec_13_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_13_MPORT_data = 1'h0;
  assign ram_exceptionVec_13_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_13_MPORT_mask = 1'h1;
  assign ram_exceptionVec_13_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_data = ram_exceptionVec_14[ram_exceptionVec_14_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_14_MPORT_data = 1'h0;
  assign ram_exceptionVec_14_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_14_MPORT_mask = 1'h1;
  assign ram_exceptionVec_14_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_data = ram_exceptionVec_15[ram_exceptionVec_15_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_15_MPORT_data = 1'h0;
  assign ram_exceptionVec_15_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_15_MPORT_mask = 1'h1;
  assign ram_exceptionVec_15_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx_io_deq_bits_MPORT_en = 1'h1;
  assign ram_brIdx_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_brIdx_io_deq_bits_MPORT_data = ram_brIdx[ram_brIdx_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign ram_brIdx_MPORT_addr = enq_ptr_value;
  assign ram_brIdx_MPORT_mask = 1'h1;
  assign ram_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_220_clock = clock;
  assign line_220_reset = reset;
  assign line_220_valid = do_enq ^ line_220_valid_reg;
  assign line_221_clock = clock;
  assign line_221_reset = reset;
  assign line_221_valid = do_deq ^ line_221_valid_reg;
  assign line_222_clock = clock;
  assign line_222_reset = reset;
  assign line_222_valid = _T ^ line_222_valid_reg;
  assign line_223_clock = clock;
  assign line_223_reset = reset;
  assign line_223_valid = io_flush ^ line_223_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/utils/FlushableQueue.scala 46:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/utils/FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_0 = ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_1 = ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_2 = ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_3 = ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_4 = ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_5 = ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_6 = ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_7 = ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_8 = ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_9 = ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_10 = ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_11 = ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_13 = ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_14 = ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_15 = ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  always @(posedge clock) begin
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pnpc_MPORT_en & ram_pnpc_MPORT_mask) begin
      ram_pnpc[ram_pnpc_MPORT_addr] <= ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_0_MPORT_en & ram_exceptionVec_0_MPORT_mask) begin
      ram_exceptionVec_0[ram_exceptionVec_0_MPORT_addr] <= ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_1_MPORT_en & ram_exceptionVec_1_MPORT_mask) begin
      ram_exceptionVec_1[ram_exceptionVec_1_MPORT_addr] <= ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_2_MPORT_en & ram_exceptionVec_2_MPORT_mask) begin
      ram_exceptionVec_2[ram_exceptionVec_2_MPORT_addr] <= ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_3_MPORT_en & ram_exceptionVec_3_MPORT_mask) begin
      ram_exceptionVec_3[ram_exceptionVec_3_MPORT_addr] <= ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_4_MPORT_en & ram_exceptionVec_4_MPORT_mask) begin
      ram_exceptionVec_4[ram_exceptionVec_4_MPORT_addr] <= ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_5_MPORT_en & ram_exceptionVec_5_MPORT_mask) begin
      ram_exceptionVec_5[ram_exceptionVec_5_MPORT_addr] <= ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_6_MPORT_en & ram_exceptionVec_6_MPORT_mask) begin
      ram_exceptionVec_6[ram_exceptionVec_6_MPORT_addr] <= ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_7_MPORT_en & ram_exceptionVec_7_MPORT_mask) begin
      ram_exceptionVec_7[ram_exceptionVec_7_MPORT_addr] <= ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_8_MPORT_en & ram_exceptionVec_8_MPORT_mask) begin
      ram_exceptionVec_8[ram_exceptionVec_8_MPORT_addr] <= ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_9_MPORT_en & ram_exceptionVec_9_MPORT_mask) begin
      ram_exceptionVec_9[ram_exceptionVec_9_MPORT_addr] <= ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_10_MPORT_en & ram_exceptionVec_10_MPORT_mask) begin
      ram_exceptionVec_10[ram_exceptionVec_10_MPORT_addr] <= ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_11_MPORT_en & ram_exceptionVec_11_MPORT_mask) begin
      ram_exceptionVec_11[ram_exceptionVec_11_MPORT_addr] <= ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_12_MPORT_en & ram_exceptionVec_12_MPORT_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12_MPORT_addr] <= ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_13_MPORT_en & ram_exceptionVec_13_MPORT_mask) begin
      ram_exceptionVec_13[ram_exceptionVec_13_MPORT_addr] <= ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_14_MPORT_en & ram_exceptionVec_14_MPORT_mask) begin
      ram_exceptionVec_14[ram_exceptionVec_14_MPORT_addr] <= ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_15_MPORT_en & ram_exceptionVec_15_MPORT_mask) begin
      ram_exceptionVec_15[ram_exceptionVec_15_MPORT_addr] <= ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_brIdx_MPORT_en & ram_brIdx_MPORT_mask) begin
      ram_brIdx[ram_brIdx_MPORT_addr] <= ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      enq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 64:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      deq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 65:21]
    end else if (do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 38:17]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/FlushableQueue.scala 26:35]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 67:16]
    end else if (do_enq != do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 41:28]
      maybe_full <= do_enq; // @[src/main/scala/utils/FlushableQueue.scala 42:16]
    end
    line_220_valid_reg <= do_enq;
    line_221_valid_reg <= do_deq;
    line_222_valid_reg <= _T;
    line_223_valid_reg <= io_flush;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_0[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_1[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_2[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_3[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_4[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_5[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_6[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_7[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_8[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_9[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_10[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_11[initvar] = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_13[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_14[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_15[initvar] = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_19[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  enq_ptr_value = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  deq_ptr_value = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  maybe_full = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_220_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_221_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_222_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_223_valid_reg = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (do_enq) begin
      cover(1'h1);
    end
    //
    if (do_deq) begin
      cover(1'h1);
    end
    //
    if (_T) begin
      cover(1'h1);
    end
    //
    if (io_flush) begin
      cover(1'h1);
    end
  end
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [86:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [86:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input         REG_actualTaken,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  output        isWFI,
  input         flushICache,
  input         flushTLB,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isMissPredict; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_actualTarget; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_actualTaken; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [6:0] ifu_REG_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [1:0] ifu_REG_btbType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isRVC; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushICache; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushTLB; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ibf_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_flush; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  idu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_isWFI_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [11:0] idu_intrVecIDU; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  ibf_io_in_q_clock; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_reset; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_flush; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  line_224_clock;
  wire  line_224_reset;
  wire  line_224_valid;
  reg  line_224_valid_reg;
  wire  _GEN_4 = _T_1 ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  line_225_clock;
  wire  line_225_reset;
  wire  line_225_valid;
  reg  line_225_valid_reg;
  wire  _GEN_5 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_4; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  wire  line_226_clock;
  wire  line_226_reset;
  wire  line_226_valid;
  reg  line_226_valid_reg;
  reg [63:0] idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  line_227_clock;
  wire  line_227_reset;
  wire  line_227_valid;
  reg  line_227_valid_reg;
  IFU_inorder ifu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ifu_io_out_bits_exceptionVec_1),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_iaf(ifu_io_iaf),
    .REG_valid(ifu_REG_valid),
    .REG_pc(ifu_REG_pc),
    .REG_isMissPredict(ifu_REG_isMissPredict),
    .REG_actualTarget(ifu_REG_actualTarget),
    .REG_actualTaken(ifu_REG_actualTaken),
    .REG_fuOpType(ifu_REG_fuOpType),
    .REG_btbType(ifu_REG_btbType),
    .REG_isRVC(ifu_REG_isRVC),
    .flushICache(ifu_flushICache),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_0(ibf_io_in_bits_exceptionVec_0),
    .io_in_bits_exceptionVec_1(ibf_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_2(ibf_io_in_bits_exceptionVec_2),
    .io_in_bits_exceptionVec_3(ibf_io_in_bits_exceptionVec_3),
    .io_in_bits_exceptionVec_4(ibf_io_in_bits_exceptionVec_4),
    .io_in_bits_exceptionVec_5(ibf_io_in_bits_exceptionVec_5),
    .io_in_bits_exceptionVec_6(ibf_io_in_bits_exceptionVec_6),
    .io_in_bits_exceptionVec_7(ibf_io_in_bits_exceptionVec_7),
    .io_in_bits_exceptionVec_8(ibf_io_in_bits_exceptionVec_8),
    .io_in_bits_exceptionVec_9(ibf_io_in_bits_exceptionVec_9),
    .io_in_bits_exceptionVec_10(ibf_io_in_bits_exceptionVec_10),
    .io_in_bits_exceptionVec_11(ibf_io_in_bits_exceptionVec_11),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_exceptionVec_13(ibf_io_in_bits_exceptionVec_13),
    .io_in_bits_exceptionVec_14(ibf_io_in_bits_exceptionVec_14),
    .io_in_bits_exceptionVec_15(ibf_io_in_bits_exceptionVec_15),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ibf_io_out_bits_exceptionVec_1),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossBoundaryFault(ibf_io_out_bits_crossBoundaryFault),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_1(idu_io_in_0_bits_exceptionVec_1),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossBoundaryFault(idu_io_in_0_bits_crossBoundaryFault),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(idu_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(idu_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_sfence_vma_invalid(idu_io_sfence_vma_invalid),
    .io_wfi_invalid(idu_io_wfi_invalid),
    .isWFI_0(idu_isWFI_0),
    .intrVecIDU(idu_intrVecIDU)
  );
  FlushableQueue ibf_io_in_q ( // @[src/main/scala/utils/FlushableQueue.scala 94:21]
    .clock(ibf_io_in_q_clock),
    .reset(ibf_io_in_q_reset),
    .io_enq_ready(ibf_io_in_q_io_enq_ready),
    .io_enq_valid(ibf_io_in_q_io_enq_valid),
    .io_enq_bits_instr(ibf_io_in_q_io_enq_bits_instr),
    .io_enq_bits_pc(ibf_io_in_q_io_enq_bits_pc),
    .io_enq_bits_pnpc(ibf_io_in_q_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_1(ibf_io_in_q_io_enq_bits_exceptionVec_1),
    .io_enq_bits_brIdx(ibf_io_in_q_io_enq_bits_brIdx),
    .io_deq_ready(ibf_io_in_q_io_deq_ready),
    .io_deq_valid(ibf_io_in_q_io_deq_valid),
    .io_deq_bits_instr(ibf_io_in_q_io_deq_bits_instr),
    .io_deq_bits_pc(ibf_io_in_q_io_deq_bits_pc),
    .io_deq_bits_pnpc(ibf_io_in_q_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_0(ibf_io_in_q_io_deq_bits_exceptionVec_0),
    .io_deq_bits_exceptionVec_1(ibf_io_in_q_io_deq_bits_exceptionVec_1),
    .io_deq_bits_exceptionVec_2(ibf_io_in_q_io_deq_bits_exceptionVec_2),
    .io_deq_bits_exceptionVec_3(ibf_io_in_q_io_deq_bits_exceptionVec_3),
    .io_deq_bits_exceptionVec_4(ibf_io_in_q_io_deq_bits_exceptionVec_4),
    .io_deq_bits_exceptionVec_5(ibf_io_in_q_io_deq_bits_exceptionVec_5),
    .io_deq_bits_exceptionVec_6(ibf_io_in_q_io_deq_bits_exceptionVec_6),
    .io_deq_bits_exceptionVec_7(ibf_io_in_q_io_deq_bits_exceptionVec_7),
    .io_deq_bits_exceptionVec_8(ibf_io_in_q_io_deq_bits_exceptionVec_8),
    .io_deq_bits_exceptionVec_9(ibf_io_in_q_io_deq_bits_exceptionVec_9),
    .io_deq_bits_exceptionVec_10(ibf_io_in_q_io_deq_bits_exceptionVec_10),
    .io_deq_bits_exceptionVec_11(ibf_io_in_q_io_deq_bits_exceptionVec_11),
    .io_deq_bits_exceptionVec_12(ibf_io_in_q_io_deq_bits_exceptionVec_12),
    .io_deq_bits_exceptionVec_13(ibf_io_in_q_io_deq_bits_exceptionVec_13),
    .io_deq_bits_exceptionVec_14(ibf_io_in_q_io_deq_bits_exceptionVec_14),
    .io_deq_bits_exceptionVec_15(ibf_io_in_q_io_deq_bits_exceptionVec_15),
    .io_deq_bits_brIdx(ibf_io_in_q_io_deq_bits_brIdx),
    .io_flush(ibf_io_in_q_io_flush)
  );
  GEN_w1_line #(.COVER_INDEX(224)) line_224 (
    .clock(line_224_clock),
    .reset(line_224_reset),
    .valid(line_224_valid)
  );
  GEN_w1_line #(.COVER_INDEX(225)) line_225 (
    .clock(line_225_clock),
    .reset(line_225_reset),
    .valid(line_225_valid)
  );
  GEN_w1_line #(.COVER_INDEX(226)) line_226 (
    .clock(line_226_clock),
    .reset(line_226_reset),
    .valid(line_226_valid)
  );
  GEN_w1_line #(.COVER_INDEX(227)) line_227 (
    .clock(line_227_clock),
    .reset(line_227_reset),
    .valid(line_227_valid)
  );
  assign line_224_clock = clock;
  assign line_224_reset = reset;
  assign line_224_valid = _T_1 ^ line_224_valid_reg;
  assign line_225_clock = clock;
  assign line_225_reset = reset;
  assign line_225_valid = _T_3 ^ line_225_valid_reg;
  assign line_226_clock = clock;
  assign line_226_reset = reset;
  assign line_226_valid = ifu_io_flushVec[1] ^ line_226_valid_reg;
  assign line_227_clock = clock;
  assign line_227_reset = reset;
  assign line_227_valid = _T_3 ^ line_227_valid_reg;
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_crossBoundaryFault = idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_isNutCoreTrap = idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_flushVec = ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:15]
  assign isWFI = idu_isWFI_0;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_out_ready = ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_iaf = io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 122:10]
  assign ifu_REG_valid = REG_valid;
  assign ifu_REG_pc = REG_pc;
  assign ifu_REG_isMissPredict = REG_isMissPredict;
  assign ifu_REG_actualTarget = REG_actualTarget;
  assign ifu_REG_actualTaken = REG_actualTaken;
  assign ifu_REG_fuOpType = REG_fuOpType;
  assign ifu_REG_btbType = REG_btbType;
  assign ifu_REG_isRVC = REG_isRVC;
  assign ifu_flushICache = flushICache;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = ibf_io_in_q_io_deq_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_instr = ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pc = ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pnpc = ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_0 = ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_1 = ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_2 = ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_3 = ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_4 = ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_5 = ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_6 = ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_7 = ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_8 = ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_9 = ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_10 = ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_11 = ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_12 = ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_13 = ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_14 = ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_15 = ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_brIdx = ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[src/main/scala/nutcore/frontend/Frontend.scala 116:34]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_1 = idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossBoundaryFault = idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign idu_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 113:29]
  assign idu_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:22]
  assign idu_intrVecIDU = intrVecIDU;
  assign ibf_io_in_q_clock = clock;
  assign ibf_io_in_q_reset = reset;
  assign ibf_io_in_q_io_enq_valid = ifu_io_out_valid; // @[src/main/scala/utils/FlushableQueue.scala 95:22]
  assign ibf_io_in_q_io_enq_bits_instr = ifu_io_out_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pc = ifu_io_out_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_exceptionVec_1 = ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_deq_ready = ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_q_io_flush = ifu_io_flushVec[0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:58]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_5;
    end
    line_224_valid_reg <= _T_1;
    line_225_valid_reg <= _T_3;
    line_226_valid_reg <= ifu_io_flushVec[1];
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_instr <= ibf_io_out_bits_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pc <= ibf_io_out_bits_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pnpc <= ibf_io_out_bits_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_1 <= ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_brIdx <= ibf_io_out_bits_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_crossBoundaryFault <= ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    line_227_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_224_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_225_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_226_valid_reg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc = _RAND_5[38:0];
  _RAND_6 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_12 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  idu_io_in_0_bits_r_crossBoundaryFault = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_227_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_3) begin
      cover(1'h1);
    end
    //
    if (ifu_io_flushVec[1]) begin
      cover(1'h1);
    end
    //
    if (_T_3) begin
      cover(1'h1);
    end
  end
endmodule
module DummyDPICWrapper(
  input         clock,
  input         reset,
  input  [63:0] io_bits_value_1, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_2, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_3, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_4, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_5, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_6, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_7, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_8, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_9, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_10, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_11, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_12, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_13, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_14, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_15, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_16, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_17, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_18, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_19, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_20, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_21, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_22, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_23, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_24, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_25, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_26, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_27, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_28, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_29, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_30, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_31 // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_0; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_1; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_2; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_3; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_4; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_5; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_6; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_7; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_8; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_9; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_10; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_11; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_12; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_13; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_14; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_15; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_16; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_17; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_18; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_19; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_20; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_21; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_22; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_23; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_24; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_25; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_26; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_27; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_28; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_29; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_30; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_31; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchIntRegState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_value_0(dpic_io_value_0),
    .io_value_1(dpic_io_value_1),
    .io_value_2(dpic_io_value_2),
    .io_value_3(dpic_io_value_3),
    .io_value_4(dpic_io_value_4),
    .io_value_5(dpic_io_value_5),
    .io_value_6(dpic_io_value_6),
    .io_value_7(dpic_io_value_7),
    .io_value_8(dpic_io_value_8),
    .io_value_9(dpic_io_value_9),
    .io_value_10(dpic_io_value_10),
    .io_value_11(dpic_io_value_11),
    .io_value_12(dpic_io_value_12),
    .io_value_13(dpic_io_value_13),
    .io_value_14(dpic_io_value_14),
    .io_value_15(dpic_io_value_15),
    .io_value_16(dpic_io_value_16),
    .io_value_17(dpic_io_value_17),
    .io_value_18(dpic_io_value_18),
    .io_value_19(dpic_io_value_19),
    .io_value_20(dpic_io_value_20),
    .io_value_21(dpic_io_value_21),
    .io_value_22(dpic_io_value_22),
    .io_value_23(dpic_io_value_23),
    .io_value_24(dpic_io_value_24),
    .io_value_25(dpic_io_value_25),
    .io_value_26(dpic_io_value_26),
    .io_value_27(dpic_io_value_27),
    .io_value_28(dpic_io_value_28),
    .io_value_29(dpic_io_value_29),
    .io_value_30(dpic_io_value_30),
    .io_value_31(dpic_io_value_31),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_value_0 = 64'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_1 = io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_2 = io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_3 = io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_4 = io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_5 = io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_6 = io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_7 = io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_8 = io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_9 = io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_10 = io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_11 = io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_12 = io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_13 = io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_14 = io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_15 = io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_16 = io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_17 = io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_18 = io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_19 = io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_20 = io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_21 = io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_22 = io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_23 = io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_24 = io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_25 = io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_26 = io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_27 = io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_28 = io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_29 = io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_30 = io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_31 = io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_flush // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  _src1ForwardNextCycle_T = ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _src1ForwardNextCycle_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 51:43]
  wire  _src1Forward_T_1 = dontForward1 ? ~src1DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _src1Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:34]
  wire  _src2Forward_T_1 = dontForward1 ? ~src2DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _src2Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:34]
  reg [31:0] busy; // @[src/main/scala/nutcore/RF.scala 38:21]
  wire [31:0] _src1Ready_T = busy >> io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/RF.scala 39:37]
  wire  src1Ready = ~_src1Ready_T[0] | src1ForwardNextCycle | src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 56:62]
  wire [31:0] _src2Ready_T = busy >> io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/RF.scala 39:37]
  wire  src2Ready = ~_src2Ready_T[0] | src2ForwardNextCycle | src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 57:62]
  reg [63:0] rf_0; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_1; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_2; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_3; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_4; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_5; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_6; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_7; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_8; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_9; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_10; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_11; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_12; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_13; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_14; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_15; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_16; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_17; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_18; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_19; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_20; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_21; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_22; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_23; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_24; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_25; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_26; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_27; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_28; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_29; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_30; // @[src/main/scala/nutcore/RF.scala 32:19]
  reg [63:0] rf_31; // @[src/main/scala/nutcore/RF.scala 32:19]
  wire  io_out_bits_data_src1_signBit = io_in_0_bits_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _io_out_bits_data_src1_T_1 = io_out_bits_data_src1_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_data_src1_T_2 = {_io_out_bits_data_src1_T_1,io_in_0_bits_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _io_out_bits_data_src1_T_3 = ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:21]
  wire  _io_out_bits_data_src1_T_4 = src1Forward & ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:18]
  wire  _io_out_bits_data_src1_T_9 = ~io_in_0_bits_ctrl_src1Type & _io_out_bits_data_src1_T_3 & ~src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 67:76]
  wire  line_228_clock;
  wire  line_228_reset;
  wire  line_228_valid;
  reg  line_228_valid_reg;
  wire  line_229_clock;
  wire  line_229_reset;
  wire  line_229_valid;
  reg  line_229_valid_reg;
  wire [63:0] _GEN_100 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_230_clock;
  wire  line_230_reset;
  wire  line_230_valid;
  reg  line_230_valid_reg;
  wire [63:0] _GEN_101 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? rf_2 : _GEN_100; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_231_clock;
  wire  line_231_reset;
  wire  line_231_valid;
  reg  line_231_valid_reg;
  wire [63:0] _GEN_102 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? rf_3 : _GEN_101; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_232_clock;
  wire  line_232_reset;
  wire  line_232_valid;
  reg  line_232_valid_reg;
  wire [63:0] _GEN_103 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? rf_4 : _GEN_102; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_233_clock;
  wire  line_233_reset;
  wire  line_233_valid;
  reg  line_233_valid_reg;
  wire [63:0] _GEN_104 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? rf_5 : _GEN_103; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_234_clock;
  wire  line_234_reset;
  wire  line_234_valid;
  reg  line_234_valid_reg;
  wire [63:0] _GEN_105 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? rf_6 : _GEN_104; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_235_clock;
  wire  line_235_reset;
  wire  line_235_valid;
  reg  line_235_valid_reg;
  wire [63:0] _GEN_106 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? rf_7 : _GEN_105; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_236_clock;
  wire  line_236_reset;
  wire  line_236_valid;
  reg  line_236_valid_reg;
  wire [63:0] _GEN_107 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? rf_8 : _GEN_106; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_237_clock;
  wire  line_237_reset;
  wire  line_237_valid;
  reg  line_237_valid_reg;
  wire [63:0] _GEN_108 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? rf_9 : _GEN_107; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_238_clock;
  wire  line_238_reset;
  wire  line_238_valid;
  reg  line_238_valid_reg;
  wire [63:0] _GEN_109 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? rf_10 : _GEN_108; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_239_clock;
  wire  line_239_reset;
  wire  line_239_valid;
  reg  line_239_valid_reg;
  wire [63:0] _GEN_110 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? rf_11 : _GEN_109; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_240_clock;
  wire  line_240_reset;
  wire  line_240_valid;
  reg  line_240_valid_reg;
  wire [63:0] _GEN_111 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? rf_12 : _GEN_110; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_241_clock;
  wire  line_241_reset;
  wire  line_241_valid;
  reg  line_241_valid_reg;
  wire [63:0] _GEN_112 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? rf_13 : _GEN_111; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_242_clock;
  wire  line_242_reset;
  wire  line_242_valid;
  reg  line_242_valid_reg;
  wire [63:0] _GEN_113 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? rf_14 : _GEN_112; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_243_clock;
  wire  line_243_reset;
  wire  line_243_valid;
  reg  line_243_valid_reg;
  wire [63:0] _GEN_114 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? rf_15 : _GEN_113; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_244_clock;
  wire  line_244_reset;
  wire  line_244_valid;
  reg  line_244_valid_reg;
  wire [63:0] _GEN_115 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? rf_16 : _GEN_114; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_245_clock;
  wire  line_245_reset;
  wire  line_245_valid;
  reg  line_245_valid_reg;
  wire [63:0] _GEN_116 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? rf_17 : _GEN_115; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_246_clock;
  wire  line_246_reset;
  wire  line_246_valid;
  reg  line_246_valid_reg;
  wire [63:0] _GEN_117 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? rf_18 : _GEN_116; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_247_clock;
  wire  line_247_reset;
  wire  line_247_valid;
  reg  line_247_valid_reg;
  wire [63:0] _GEN_118 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? rf_19 : _GEN_117; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_248_clock;
  wire  line_248_reset;
  wire  line_248_valid;
  reg  line_248_valid_reg;
  wire [63:0] _GEN_119 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? rf_20 : _GEN_118; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_249_clock;
  wire  line_249_reset;
  wire  line_249_valid;
  reg  line_249_valid_reg;
  wire [63:0] _GEN_120 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? rf_21 : _GEN_119; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_250_clock;
  wire  line_250_reset;
  wire  line_250_valid;
  reg  line_250_valid_reg;
  wire [63:0] _GEN_121 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? rf_22 : _GEN_120; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_251_clock;
  wire  line_251_reset;
  wire  line_251_valid;
  reg  line_251_valid_reg;
  wire [63:0] _GEN_122 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? rf_23 : _GEN_121; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_252_clock;
  wire  line_252_reset;
  wire  line_252_valid;
  reg  line_252_valid_reg;
  wire [63:0] _GEN_123 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? rf_24 : _GEN_122; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_253_clock;
  wire  line_253_reset;
  wire  line_253_valid;
  reg  line_253_valid_reg;
  wire [63:0] _GEN_124 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? rf_25 : _GEN_123; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_254_clock;
  wire  line_254_reset;
  wire  line_254_valid;
  reg  line_254_valid_reg;
  wire [63:0] _GEN_125 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? rf_26 : _GEN_124; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_255_clock;
  wire  line_255_reset;
  wire  line_255_valid;
  reg  line_255_valid_reg;
  wire [63:0] _GEN_126 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? rf_27 : _GEN_125; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_256_clock;
  wire  line_256_reset;
  wire  line_256_valid;
  reg  line_256_valid_reg;
  wire [63:0] _GEN_127 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? rf_28 : _GEN_126; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_257_clock;
  wire  line_257_reset;
  wire  line_257_valid;
  reg  line_257_valid_reg;
  wire [63:0] _GEN_128 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? rf_29 : _GEN_127; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_258_clock;
  wire  line_258_reset;
  wire  line_258_valid;
  reg  line_258_valid_reg;
  wire [63:0] _GEN_129 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? rf_30 : _GEN_128; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_259_clock;
  wire  line_259_reset;
  wire  line_259_valid;
  reg  line_259_valid_reg;
  wire [63:0] _GEN_130 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? rf_31 : _GEN_129; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire [63:0] _io_out_bits_data_src1_T_11 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : _GEN_130; // @[src/main/scala/nutcore/RF.scala 33:36]
  wire [63:0] _io_out_bits_data_src1_T_12 = io_in_0_bits_ctrl_src1Type ? _io_out_bits_data_src1_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_13 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_14 = _io_out_bits_data_src1_T_4 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_15 = _io_out_bits_data_src1_T_9 ? _io_out_bits_data_src1_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_16 = _io_out_bits_data_src1_T_12 | _io_out_bits_data_src1_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_17 = _io_out_bits_data_src1_T_16 | _io_out_bits_data_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_bits_data_src2_T_1 = ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:21]
  wire  _io_out_bits_data_src2_T_2 = src2Forward & ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:18]
  wire  _io_out_bits_data_src2_T_7 = ~io_in_0_bits_ctrl_src2Type & _io_out_bits_data_src2_T_1 & ~src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 73:77]
  wire  line_260_clock;
  wire  line_260_reset;
  wire  line_260_valid;
  reg  line_260_valid_reg;
  wire  line_261_clock;
  wire  line_261_reset;
  wire  line_261_valid;
  reg  line_261_valid_reg;
  wire [63:0] _GEN_132 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_262_clock;
  wire  line_262_reset;
  wire  line_262_valid;
  reg  line_262_valid_reg;
  wire [63:0] _GEN_133 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? rf_2 : _GEN_132; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_263_clock;
  wire  line_263_reset;
  wire  line_263_valid;
  reg  line_263_valid_reg;
  wire [63:0] _GEN_134 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? rf_3 : _GEN_133; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_264_clock;
  wire  line_264_reset;
  wire  line_264_valid;
  reg  line_264_valid_reg;
  wire [63:0] _GEN_135 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? rf_4 : _GEN_134; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_265_clock;
  wire  line_265_reset;
  wire  line_265_valid;
  reg  line_265_valid_reg;
  wire [63:0] _GEN_136 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? rf_5 : _GEN_135; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_266_clock;
  wire  line_266_reset;
  wire  line_266_valid;
  reg  line_266_valid_reg;
  wire [63:0] _GEN_137 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? rf_6 : _GEN_136; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_267_clock;
  wire  line_267_reset;
  wire  line_267_valid;
  reg  line_267_valid_reg;
  wire [63:0] _GEN_138 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? rf_7 : _GEN_137; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_268_clock;
  wire  line_268_reset;
  wire  line_268_valid;
  reg  line_268_valid_reg;
  wire [63:0] _GEN_139 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? rf_8 : _GEN_138; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_269_clock;
  wire  line_269_reset;
  wire  line_269_valid;
  reg  line_269_valid_reg;
  wire [63:0] _GEN_140 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? rf_9 : _GEN_139; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_270_clock;
  wire  line_270_reset;
  wire  line_270_valid;
  reg  line_270_valid_reg;
  wire [63:0] _GEN_141 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? rf_10 : _GEN_140; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_271_clock;
  wire  line_271_reset;
  wire  line_271_valid;
  reg  line_271_valid_reg;
  wire [63:0] _GEN_142 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? rf_11 : _GEN_141; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_272_clock;
  wire  line_272_reset;
  wire  line_272_valid;
  reg  line_272_valid_reg;
  wire [63:0] _GEN_143 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? rf_12 : _GEN_142; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_273_clock;
  wire  line_273_reset;
  wire  line_273_valid;
  reg  line_273_valid_reg;
  wire [63:0] _GEN_144 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? rf_13 : _GEN_143; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_274_clock;
  wire  line_274_reset;
  wire  line_274_valid;
  reg  line_274_valid_reg;
  wire [63:0] _GEN_145 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? rf_14 : _GEN_144; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_275_clock;
  wire  line_275_reset;
  wire  line_275_valid;
  reg  line_275_valid_reg;
  wire [63:0] _GEN_146 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? rf_15 : _GEN_145; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_276_clock;
  wire  line_276_reset;
  wire  line_276_valid;
  reg  line_276_valid_reg;
  wire [63:0] _GEN_147 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? rf_16 : _GEN_146; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_277_clock;
  wire  line_277_reset;
  wire  line_277_valid;
  reg  line_277_valid_reg;
  wire [63:0] _GEN_148 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? rf_17 : _GEN_147; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_278_clock;
  wire  line_278_reset;
  wire  line_278_valid;
  reg  line_278_valid_reg;
  wire [63:0] _GEN_149 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? rf_18 : _GEN_148; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_279_clock;
  wire  line_279_reset;
  wire  line_279_valid;
  reg  line_279_valid_reg;
  wire [63:0] _GEN_150 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? rf_19 : _GEN_149; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_280_clock;
  wire  line_280_reset;
  wire  line_280_valid;
  reg  line_280_valid_reg;
  wire [63:0] _GEN_151 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? rf_20 : _GEN_150; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_281_clock;
  wire  line_281_reset;
  wire  line_281_valid;
  reg  line_281_valid_reg;
  wire [63:0] _GEN_152 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? rf_21 : _GEN_151; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_282_clock;
  wire  line_282_reset;
  wire  line_282_valid;
  reg  line_282_valid_reg;
  wire [63:0] _GEN_153 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? rf_22 : _GEN_152; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_283_clock;
  wire  line_283_reset;
  wire  line_283_valid;
  reg  line_283_valid_reg;
  wire [63:0] _GEN_154 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? rf_23 : _GEN_153; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_284_clock;
  wire  line_284_reset;
  wire  line_284_valid;
  reg  line_284_valid_reg;
  wire [63:0] _GEN_155 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? rf_24 : _GEN_154; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_285_clock;
  wire  line_285_reset;
  wire  line_285_valid;
  reg  line_285_valid_reg;
  wire [63:0] _GEN_156 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? rf_25 : _GEN_155; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_286_clock;
  wire  line_286_reset;
  wire  line_286_valid;
  reg  line_286_valid_reg;
  wire [63:0] _GEN_157 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? rf_26 : _GEN_156; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_287_clock;
  wire  line_287_reset;
  wire  line_287_valid;
  reg  line_287_valid_reg;
  wire [63:0] _GEN_158 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? rf_27 : _GEN_157; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_288_clock;
  wire  line_288_reset;
  wire  line_288_valid;
  reg  line_288_valid_reg;
  wire [63:0] _GEN_159 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? rf_28 : _GEN_158; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_289_clock;
  wire  line_289_reset;
  wire  line_289_valid;
  reg  line_289_valid_reg;
  wire [63:0] _GEN_160 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? rf_29 : _GEN_159; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_290_clock;
  wire  line_290_reset;
  wire  line_290_valid;
  reg  line_290_valid_reg;
  wire [63:0] _GEN_161 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? rf_30 : _GEN_160; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire  line_291_clock;
  wire  line_291_reset;
  wire  line_291_valid;
  reg  line_291_valid_reg;
  wire [63:0] _GEN_162 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? rf_31 : _GEN_161; // @[src/main/scala/nutcore/RF.scala 33:{36,36}]
  wire [63:0] _io_out_bits_data_src2_T_9 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : _GEN_162; // @[src/main/scala/nutcore/RF.scala 33:36]
  wire [63:0] _io_out_bits_data_src2_T_10 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_11 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_12 = _io_out_bits_data_src2_T_2 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_13 = _io_out_bits_data_src2_T_7 ? _io_out_bits_data_src2_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_14 = _io_out_bits_data_src2_T_10 | _io_out_bits_data_src2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_15 = _io_out_bits_data_src2_T_14 | _io_out_bits_data_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  line_292_clock;
  wire  line_292_reset;
  wire  line_292_valid;
  reg  line_292_valid_reg;
  wire  _GEN_64 = 5'h0 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_293_clock;
  wire  line_293_reset;
  wire  line_293_valid;
  reg  line_293_valid_reg;
  wire  _GEN_65 = 5'h1 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_294_clock;
  wire  line_294_reset;
  wire  line_294_valid;
  reg  line_294_valid_reg;
  wire  _GEN_66 = 5'h2 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_295_clock;
  wire  line_295_reset;
  wire  line_295_valid;
  reg  line_295_valid_reg;
  wire  _GEN_67 = 5'h3 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_296_clock;
  wire  line_296_reset;
  wire  line_296_valid;
  reg  line_296_valid_reg;
  wire  _GEN_68 = 5'h4 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_297_clock;
  wire  line_297_reset;
  wire  line_297_valid;
  reg  line_297_valid_reg;
  wire  _GEN_69 = 5'h5 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_298_clock;
  wire  line_298_reset;
  wire  line_298_valid;
  reg  line_298_valid_reg;
  wire  _GEN_70 = 5'h6 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_299_clock;
  wire  line_299_reset;
  wire  line_299_valid;
  reg  line_299_valid_reg;
  wire  _GEN_71 = 5'h7 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_300_clock;
  wire  line_300_reset;
  wire  line_300_valid;
  reg  line_300_valid_reg;
  wire  _GEN_72 = 5'h8 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_301_clock;
  wire  line_301_reset;
  wire  line_301_valid;
  reg  line_301_valid_reg;
  wire  _GEN_73 = 5'h9 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_302_clock;
  wire  line_302_reset;
  wire  line_302_valid;
  reg  line_302_valid_reg;
  wire  _GEN_74 = 5'ha == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_303_clock;
  wire  line_303_reset;
  wire  line_303_valid;
  reg  line_303_valid_reg;
  wire  _GEN_75 = 5'hb == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_304_clock;
  wire  line_304_reset;
  wire  line_304_valid;
  reg  line_304_valid_reg;
  wire  _GEN_76 = 5'hc == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_305_clock;
  wire  line_305_reset;
  wire  line_305_valid;
  reg  line_305_valid_reg;
  wire  _GEN_77 = 5'hd == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_306_clock;
  wire  line_306_reset;
  wire  line_306_valid;
  reg  line_306_valid_reg;
  wire  _GEN_78 = 5'he == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_307_clock;
  wire  line_307_reset;
  wire  line_307_valid;
  reg  line_307_valid_reg;
  wire  _GEN_79 = 5'hf == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_308_clock;
  wire  line_308_reset;
  wire  line_308_valid;
  reg  line_308_valid_reg;
  wire  _GEN_80 = 5'h10 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_309_clock;
  wire  line_309_reset;
  wire  line_309_valid;
  reg  line_309_valid_reg;
  wire  _GEN_81 = 5'h11 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_310_clock;
  wire  line_310_reset;
  wire  line_310_valid;
  reg  line_310_valid_reg;
  wire  _GEN_82 = 5'h12 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_311_clock;
  wire  line_311_reset;
  wire  line_311_valid;
  reg  line_311_valid_reg;
  wire  _GEN_83 = 5'h13 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_312_clock;
  wire  line_312_reset;
  wire  line_312_valid;
  reg  line_312_valid_reg;
  wire  _GEN_84 = 5'h14 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_313_clock;
  wire  line_313_reset;
  wire  line_313_valid;
  reg  line_313_valid_reg;
  wire  _GEN_85 = 5'h15 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_314_clock;
  wire  line_314_reset;
  wire  line_314_valid;
  reg  line_314_valid_reg;
  wire  _GEN_86 = 5'h16 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_315_clock;
  wire  line_315_reset;
  wire  line_315_valid;
  reg  line_315_valid_reg;
  wire  _GEN_87 = 5'h17 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_316_clock;
  wire  line_316_reset;
  wire  line_316_valid;
  reg  line_316_valid_reg;
  wire  _GEN_88 = 5'h18 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_317_clock;
  wire  line_317_reset;
  wire  line_317_valid;
  reg  line_317_valid_reg;
  wire  _GEN_89 = 5'h19 == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_318_clock;
  wire  line_318_reset;
  wire  line_318_valid;
  reg  line_318_valid_reg;
  wire  _GEN_90 = 5'h1a == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_319_clock;
  wire  line_319_reset;
  wire  line_319_valid;
  reg  line_319_valid_reg;
  wire  _GEN_91 = 5'h1b == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_320_clock;
  wire  line_320_reset;
  wire  line_320_valid;
  reg  line_320_valid_reg;
  wire  _GEN_92 = 5'h1c == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_321_clock;
  wire  line_321_reset;
  wire  line_321_valid;
  reg  line_321_valid_reg;
  wire  _GEN_93 = 5'h1d == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_322_clock;
  wire  line_322_reset;
  wire  line_322_valid;
  reg  line_322_valid_reg;
  wire  _GEN_94 = 5'h1e == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_323_clock;
  wire  line_323_reset;
  wire  line_323_valid;
  reg  line_323_valid_reg;
  wire  _GEN_95 = 5'h1f == io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 34:50]
  wire  line_324_clock;
  wire  line_324_reset;
  wire  line_324_valid;
  reg  line_324_valid_reg;
  wire  _wbClearMask_T_3 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire [62:0] _wbClearMask_T_6 = 63'h1 << io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 40:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_wbClearMask_T_3 ? _wbClearMask_T_6[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 85:24]
  wire  _isuFireSetMask_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [62:0] _isuFireSetMask_T_1 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/RF.scala 40:39]
  wire [31:0] isuFireSetMask = _isuFireSetMask_T ? _isuFireSetMask_T_1[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 87:27]
  wire  line_325_clock;
  wire  line_325_reset;
  wire  line_325_valid;
  reg  line_325_valid_reg;
  wire  line_326_clock;
  wire  line_326_reset;
  wire  line_326_valid;
  reg  line_326_valid_reg;
  wire [31:0] _busy_T_5 = ~wbClearMask; // @[src/main/scala/nutcore/RF.scala 46:26]
  wire [31:0] _busy_T_6 = busy & _busy_T_5; // @[src/main/scala/nutcore/RF.scala 46:24]
  wire [31:0] _busy_T_7 = _busy_T_6 | isuFireSetMask; // @[src/main/scala/nutcore/RF.scala 46:38]
  wire [31:0] _busy_T_9 = {_busy_T_7[31:1],1'h0}; // @[src/main/scala/nutcore/RF.scala 46:16]
  wire  _T_3 = io_in_0_valid & ~io_out_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 97:40]
  wire  _T_6 = io_out_valid & ~_isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 98:38]
  wire  _T_7 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  DummyDPICWrapper difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_value_1(difftest_module_io_bits_value_1),
    .io_bits_value_2(difftest_module_io_bits_value_2),
    .io_bits_value_3(difftest_module_io_bits_value_3),
    .io_bits_value_4(difftest_module_io_bits_value_4),
    .io_bits_value_5(difftest_module_io_bits_value_5),
    .io_bits_value_6(difftest_module_io_bits_value_6),
    .io_bits_value_7(difftest_module_io_bits_value_7),
    .io_bits_value_8(difftest_module_io_bits_value_8),
    .io_bits_value_9(difftest_module_io_bits_value_9),
    .io_bits_value_10(difftest_module_io_bits_value_10),
    .io_bits_value_11(difftest_module_io_bits_value_11),
    .io_bits_value_12(difftest_module_io_bits_value_12),
    .io_bits_value_13(difftest_module_io_bits_value_13),
    .io_bits_value_14(difftest_module_io_bits_value_14),
    .io_bits_value_15(difftest_module_io_bits_value_15),
    .io_bits_value_16(difftest_module_io_bits_value_16),
    .io_bits_value_17(difftest_module_io_bits_value_17),
    .io_bits_value_18(difftest_module_io_bits_value_18),
    .io_bits_value_19(difftest_module_io_bits_value_19),
    .io_bits_value_20(difftest_module_io_bits_value_20),
    .io_bits_value_21(difftest_module_io_bits_value_21),
    .io_bits_value_22(difftest_module_io_bits_value_22),
    .io_bits_value_23(difftest_module_io_bits_value_23),
    .io_bits_value_24(difftest_module_io_bits_value_24),
    .io_bits_value_25(difftest_module_io_bits_value_25),
    .io_bits_value_26(difftest_module_io_bits_value_26),
    .io_bits_value_27(difftest_module_io_bits_value_27),
    .io_bits_value_28(difftest_module_io_bits_value_28),
    .io_bits_value_29(difftest_module_io_bits_value_29),
    .io_bits_value_30(difftest_module_io_bits_value_30),
    .io_bits_value_31(difftest_module_io_bits_value_31)
  );
  GEN_w1_line #(.COVER_INDEX(228)) line_228 (
    .clock(line_228_clock),
    .reset(line_228_reset),
    .valid(line_228_valid)
  );
  GEN_w1_line #(.COVER_INDEX(229)) line_229 (
    .clock(line_229_clock),
    .reset(line_229_reset),
    .valid(line_229_valid)
  );
  GEN_w1_line #(.COVER_INDEX(230)) line_230 (
    .clock(line_230_clock),
    .reset(line_230_reset),
    .valid(line_230_valid)
  );
  GEN_w1_line #(.COVER_INDEX(231)) line_231 (
    .clock(line_231_clock),
    .reset(line_231_reset),
    .valid(line_231_valid)
  );
  GEN_w1_line #(.COVER_INDEX(232)) line_232 (
    .clock(line_232_clock),
    .reset(line_232_reset),
    .valid(line_232_valid)
  );
  GEN_w1_line #(.COVER_INDEX(233)) line_233 (
    .clock(line_233_clock),
    .reset(line_233_reset),
    .valid(line_233_valid)
  );
  GEN_w1_line #(.COVER_INDEX(234)) line_234 (
    .clock(line_234_clock),
    .reset(line_234_reset),
    .valid(line_234_valid)
  );
  GEN_w1_line #(.COVER_INDEX(235)) line_235 (
    .clock(line_235_clock),
    .reset(line_235_reset),
    .valid(line_235_valid)
  );
  GEN_w1_line #(.COVER_INDEX(236)) line_236 (
    .clock(line_236_clock),
    .reset(line_236_reset),
    .valid(line_236_valid)
  );
  GEN_w1_line #(.COVER_INDEX(237)) line_237 (
    .clock(line_237_clock),
    .reset(line_237_reset),
    .valid(line_237_valid)
  );
  GEN_w1_line #(.COVER_INDEX(238)) line_238 (
    .clock(line_238_clock),
    .reset(line_238_reset),
    .valid(line_238_valid)
  );
  GEN_w1_line #(.COVER_INDEX(239)) line_239 (
    .clock(line_239_clock),
    .reset(line_239_reset),
    .valid(line_239_valid)
  );
  GEN_w1_line #(.COVER_INDEX(240)) line_240 (
    .clock(line_240_clock),
    .reset(line_240_reset),
    .valid(line_240_valid)
  );
  GEN_w1_line #(.COVER_INDEX(241)) line_241 (
    .clock(line_241_clock),
    .reset(line_241_reset),
    .valid(line_241_valid)
  );
  GEN_w1_line #(.COVER_INDEX(242)) line_242 (
    .clock(line_242_clock),
    .reset(line_242_reset),
    .valid(line_242_valid)
  );
  GEN_w1_line #(.COVER_INDEX(243)) line_243 (
    .clock(line_243_clock),
    .reset(line_243_reset),
    .valid(line_243_valid)
  );
  GEN_w1_line #(.COVER_INDEX(244)) line_244 (
    .clock(line_244_clock),
    .reset(line_244_reset),
    .valid(line_244_valid)
  );
  GEN_w1_line #(.COVER_INDEX(245)) line_245 (
    .clock(line_245_clock),
    .reset(line_245_reset),
    .valid(line_245_valid)
  );
  GEN_w1_line #(.COVER_INDEX(246)) line_246 (
    .clock(line_246_clock),
    .reset(line_246_reset),
    .valid(line_246_valid)
  );
  GEN_w1_line #(.COVER_INDEX(247)) line_247 (
    .clock(line_247_clock),
    .reset(line_247_reset),
    .valid(line_247_valid)
  );
  GEN_w1_line #(.COVER_INDEX(248)) line_248 (
    .clock(line_248_clock),
    .reset(line_248_reset),
    .valid(line_248_valid)
  );
  GEN_w1_line #(.COVER_INDEX(249)) line_249 (
    .clock(line_249_clock),
    .reset(line_249_reset),
    .valid(line_249_valid)
  );
  GEN_w1_line #(.COVER_INDEX(250)) line_250 (
    .clock(line_250_clock),
    .reset(line_250_reset),
    .valid(line_250_valid)
  );
  GEN_w1_line #(.COVER_INDEX(251)) line_251 (
    .clock(line_251_clock),
    .reset(line_251_reset),
    .valid(line_251_valid)
  );
  GEN_w1_line #(.COVER_INDEX(252)) line_252 (
    .clock(line_252_clock),
    .reset(line_252_reset),
    .valid(line_252_valid)
  );
  GEN_w1_line #(.COVER_INDEX(253)) line_253 (
    .clock(line_253_clock),
    .reset(line_253_reset),
    .valid(line_253_valid)
  );
  GEN_w1_line #(.COVER_INDEX(254)) line_254 (
    .clock(line_254_clock),
    .reset(line_254_reset),
    .valid(line_254_valid)
  );
  GEN_w1_line #(.COVER_INDEX(255)) line_255 (
    .clock(line_255_clock),
    .reset(line_255_reset),
    .valid(line_255_valid)
  );
  GEN_w1_line #(.COVER_INDEX(256)) line_256 (
    .clock(line_256_clock),
    .reset(line_256_reset),
    .valid(line_256_valid)
  );
  GEN_w1_line #(.COVER_INDEX(257)) line_257 (
    .clock(line_257_clock),
    .reset(line_257_reset),
    .valid(line_257_valid)
  );
  GEN_w1_line #(.COVER_INDEX(258)) line_258 (
    .clock(line_258_clock),
    .reset(line_258_reset),
    .valid(line_258_valid)
  );
  GEN_w1_line #(.COVER_INDEX(259)) line_259 (
    .clock(line_259_clock),
    .reset(line_259_reset),
    .valid(line_259_valid)
  );
  GEN_w1_line #(.COVER_INDEX(260)) line_260 (
    .clock(line_260_clock),
    .reset(line_260_reset),
    .valid(line_260_valid)
  );
  GEN_w1_line #(.COVER_INDEX(261)) line_261 (
    .clock(line_261_clock),
    .reset(line_261_reset),
    .valid(line_261_valid)
  );
  GEN_w1_line #(.COVER_INDEX(262)) line_262 (
    .clock(line_262_clock),
    .reset(line_262_reset),
    .valid(line_262_valid)
  );
  GEN_w1_line #(.COVER_INDEX(263)) line_263 (
    .clock(line_263_clock),
    .reset(line_263_reset),
    .valid(line_263_valid)
  );
  GEN_w1_line #(.COVER_INDEX(264)) line_264 (
    .clock(line_264_clock),
    .reset(line_264_reset),
    .valid(line_264_valid)
  );
  GEN_w1_line #(.COVER_INDEX(265)) line_265 (
    .clock(line_265_clock),
    .reset(line_265_reset),
    .valid(line_265_valid)
  );
  GEN_w1_line #(.COVER_INDEX(266)) line_266 (
    .clock(line_266_clock),
    .reset(line_266_reset),
    .valid(line_266_valid)
  );
  GEN_w1_line #(.COVER_INDEX(267)) line_267 (
    .clock(line_267_clock),
    .reset(line_267_reset),
    .valid(line_267_valid)
  );
  GEN_w1_line #(.COVER_INDEX(268)) line_268 (
    .clock(line_268_clock),
    .reset(line_268_reset),
    .valid(line_268_valid)
  );
  GEN_w1_line #(.COVER_INDEX(269)) line_269 (
    .clock(line_269_clock),
    .reset(line_269_reset),
    .valid(line_269_valid)
  );
  GEN_w1_line #(.COVER_INDEX(270)) line_270 (
    .clock(line_270_clock),
    .reset(line_270_reset),
    .valid(line_270_valid)
  );
  GEN_w1_line #(.COVER_INDEX(271)) line_271 (
    .clock(line_271_clock),
    .reset(line_271_reset),
    .valid(line_271_valid)
  );
  GEN_w1_line #(.COVER_INDEX(272)) line_272 (
    .clock(line_272_clock),
    .reset(line_272_reset),
    .valid(line_272_valid)
  );
  GEN_w1_line #(.COVER_INDEX(273)) line_273 (
    .clock(line_273_clock),
    .reset(line_273_reset),
    .valid(line_273_valid)
  );
  GEN_w1_line #(.COVER_INDEX(274)) line_274 (
    .clock(line_274_clock),
    .reset(line_274_reset),
    .valid(line_274_valid)
  );
  GEN_w1_line #(.COVER_INDEX(275)) line_275 (
    .clock(line_275_clock),
    .reset(line_275_reset),
    .valid(line_275_valid)
  );
  GEN_w1_line #(.COVER_INDEX(276)) line_276 (
    .clock(line_276_clock),
    .reset(line_276_reset),
    .valid(line_276_valid)
  );
  GEN_w1_line #(.COVER_INDEX(277)) line_277 (
    .clock(line_277_clock),
    .reset(line_277_reset),
    .valid(line_277_valid)
  );
  GEN_w1_line #(.COVER_INDEX(278)) line_278 (
    .clock(line_278_clock),
    .reset(line_278_reset),
    .valid(line_278_valid)
  );
  GEN_w1_line #(.COVER_INDEX(279)) line_279 (
    .clock(line_279_clock),
    .reset(line_279_reset),
    .valid(line_279_valid)
  );
  GEN_w1_line #(.COVER_INDEX(280)) line_280 (
    .clock(line_280_clock),
    .reset(line_280_reset),
    .valid(line_280_valid)
  );
  GEN_w1_line #(.COVER_INDEX(281)) line_281 (
    .clock(line_281_clock),
    .reset(line_281_reset),
    .valid(line_281_valid)
  );
  GEN_w1_line #(.COVER_INDEX(282)) line_282 (
    .clock(line_282_clock),
    .reset(line_282_reset),
    .valid(line_282_valid)
  );
  GEN_w1_line #(.COVER_INDEX(283)) line_283 (
    .clock(line_283_clock),
    .reset(line_283_reset),
    .valid(line_283_valid)
  );
  GEN_w1_line #(.COVER_INDEX(284)) line_284 (
    .clock(line_284_clock),
    .reset(line_284_reset),
    .valid(line_284_valid)
  );
  GEN_w1_line #(.COVER_INDEX(285)) line_285 (
    .clock(line_285_clock),
    .reset(line_285_reset),
    .valid(line_285_valid)
  );
  GEN_w1_line #(.COVER_INDEX(286)) line_286 (
    .clock(line_286_clock),
    .reset(line_286_reset),
    .valid(line_286_valid)
  );
  GEN_w1_line #(.COVER_INDEX(287)) line_287 (
    .clock(line_287_clock),
    .reset(line_287_reset),
    .valid(line_287_valid)
  );
  GEN_w1_line #(.COVER_INDEX(288)) line_288 (
    .clock(line_288_clock),
    .reset(line_288_reset),
    .valid(line_288_valid)
  );
  GEN_w1_line #(.COVER_INDEX(289)) line_289 (
    .clock(line_289_clock),
    .reset(line_289_reset),
    .valid(line_289_valid)
  );
  GEN_w1_line #(.COVER_INDEX(290)) line_290 (
    .clock(line_290_clock),
    .reset(line_290_reset),
    .valid(line_290_valid)
  );
  GEN_w1_line #(.COVER_INDEX(291)) line_291 (
    .clock(line_291_clock),
    .reset(line_291_reset),
    .valid(line_291_valid)
  );
  GEN_w1_line #(.COVER_INDEX(292)) line_292 (
    .clock(line_292_clock),
    .reset(line_292_reset),
    .valid(line_292_valid)
  );
  GEN_w1_line #(.COVER_INDEX(293)) line_293 (
    .clock(line_293_clock),
    .reset(line_293_reset),
    .valid(line_293_valid)
  );
  GEN_w1_line #(.COVER_INDEX(294)) line_294 (
    .clock(line_294_clock),
    .reset(line_294_reset),
    .valid(line_294_valid)
  );
  GEN_w1_line #(.COVER_INDEX(295)) line_295 (
    .clock(line_295_clock),
    .reset(line_295_reset),
    .valid(line_295_valid)
  );
  GEN_w1_line #(.COVER_INDEX(296)) line_296 (
    .clock(line_296_clock),
    .reset(line_296_reset),
    .valid(line_296_valid)
  );
  GEN_w1_line #(.COVER_INDEX(297)) line_297 (
    .clock(line_297_clock),
    .reset(line_297_reset),
    .valid(line_297_valid)
  );
  GEN_w1_line #(.COVER_INDEX(298)) line_298 (
    .clock(line_298_clock),
    .reset(line_298_reset),
    .valid(line_298_valid)
  );
  GEN_w1_line #(.COVER_INDEX(299)) line_299 (
    .clock(line_299_clock),
    .reset(line_299_reset),
    .valid(line_299_valid)
  );
  GEN_w1_line #(.COVER_INDEX(300)) line_300 (
    .clock(line_300_clock),
    .reset(line_300_reset),
    .valid(line_300_valid)
  );
  GEN_w1_line #(.COVER_INDEX(301)) line_301 (
    .clock(line_301_clock),
    .reset(line_301_reset),
    .valid(line_301_valid)
  );
  GEN_w1_line #(.COVER_INDEX(302)) line_302 (
    .clock(line_302_clock),
    .reset(line_302_reset),
    .valid(line_302_valid)
  );
  GEN_w1_line #(.COVER_INDEX(303)) line_303 (
    .clock(line_303_clock),
    .reset(line_303_reset),
    .valid(line_303_valid)
  );
  GEN_w1_line #(.COVER_INDEX(304)) line_304 (
    .clock(line_304_clock),
    .reset(line_304_reset),
    .valid(line_304_valid)
  );
  GEN_w1_line #(.COVER_INDEX(305)) line_305 (
    .clock(line_305_clock),
    .reset(line_305_reset),
    .valid(line_305_valid)
  );
  GEN_w1_line #(.COVER_INDEX(306)) line_306 (
    .clock(line_306_clock),
    .reset(line_306_reset),
    .valid(line_306_valid)
  );
  GEN_w1_line #(.COVER_INDEX(307)) line_307 (
    .clock(line_307_clock),
    .reset(line_307_reset),
    .valid(line_307_valid)
  );
  GEN_w1_line #(.COVER_INDEX(308)) line_308 (
    .clock(line_308_clock),
    .reset(line_308_reset),
    .valid(line_308_valid)
  );
  GEN_w1_line #(.COVER_INDEX(309)) line_309 (
    .clock(line_309_clock),
    .reset(line_309_reset),
    .valid(line_309_valid)
  );
  GEN_w1_line #(.COVER_INDEX(310)) line_310 (
    .clock(line_310_clock),
    .reset(line_310_reset),
    .valid(line_310_valid)
  );
  GEN_w1_line #(.COVER_INDEX(311)) line_311 (
    .clock(line_311_clock),
    .reset(line_311_reset),
    .valid(line_311_valid)
  );
  GEN_w1_line #(.COVER_INDEX(312)) line_312 (
    .clock(line_312_clock),
    .reset(line_312_reset),
    .valid(line_312_valid)
  );
  GEN_w1_line #(.COVER_INDEX(313)) line_313 (
    .clock(line_313_clock),
    .reset(line_313_reset),
    .valid(line_313_valid)
  );
  GEN_w1_line #(.COVER_INDEX(314)) line_314 (
    .clock(line_314_clock),
    .reset(line_314_reset),
    .valid(line_314_valid)
  );
  GEN_w1_line #(.COVER_INDEX(315)) line_315 (
    .clock(line_315_clock),
    .reset(line_315_reset),
    .valid(line_315_valid)
  );
  GEN_w1_line #(.COVER_INDEX(316)) line_316 (
    .clock(line_316_clock),
    .reset(line_316_reset),
    .valid(line_316_valid)
  );
  GEN_w1_line #(.COVER_INDEX(317)) line_317 (
    .clock(line_317_clock),
    .reset(line_317_reset),
    .valid(line_317_valid)
  );
  GEN_w1_line #(.COVER_INDEX(318)) line_318 (
    .clock(line_318_clock),
    .reset(line_318_reset),
    .valid(line_318_valid)
  );
  GEN_w1_line #(.COVER_INDEX(319)) line_319 (
    .clock(line_319_clock),
    .reset(line_319_reset),
    .valid(line_319_valid)
  );
  GEN_w1_line #(.COVER_INDEX(320)) line_320 (
    .clock(line_320_clock),
    .reset(line_320_reset),
    .valid(line_320_valid)
  );
  GEN_w1_line #(.COVER_INDEX(321)) line_321 (
    .clock(line_321_clock),
    .reset(line_321_reset),
    .valid(line_321_valid)
  );
  GEN_w1_line #(.COVER_INDEX(322)) line_322 (
    .clock(line_322_clock),
    .reset(line_322_reset),
    .valid(line_322_valid)
  );
  GEN_w1_line #(.COVER_INDEX(323)) line_323 (
    .clock(line_323_clock),
    .reset(line_323_reset),
    .valid(line_323_valid)
  );
  GEN_w1_line #(.COVER_INDEX(324)) line_324 (
    .clock(line_324_clock),
    .reset(line_324_reset),
    .valid(line_324_valid)
  );
  GEN_w1_line #(.COVER_INDEX(325)) line_325 (
    .clock(line_325_clock),
    .reset(line_325_reset),
    .valid(line_325_valid)
  );
  GEN_w1_line #(.COVER_INDEX(326)) line_326 (
    .clock(line_326_clock),
    .reset(line_326_reset),
    .valid(line_326_valid)
  );
  assign line_228_clock = clock;
  assign line_228_reset = reset;
  assign line_228_valid = 5'h0 == io_in_0_bits_ctrl_rfSrc1 ^ line_228_valid_reg;
  assign line_229_clock = clock;
  assign line_229_reset = reset;
  assign line_229_valid = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ^ line_229_valid_reg;
  assign line_230_clock = clock;
  assign line_230_reset = reset;
  assign line_230_valid = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ^ line_230_valid_reg;
  assign line_231_clock = clock;
  assign line_231_reset = reset;
  assign line_231_valid = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ^ line_231_valid_reg;
  assign line_232_clock = clock;
  assign line_232_reset = reset;
  assign line_232_valid = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ^ line_232_valid_reg;
  assign line_233_clock = clock;
  assign line_233_reset = reset;
  assign line_233_valid = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ^ line_233_valid_reg;
  assign line_234_clock = clock;
  assign line_234_reset = reset;
  assign line_234_valid = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ^ line_234_valid_reg;
  assign line_235_clock = clock;
  assign line_235_reset = reset;
  assign line_235_valid = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ^ line_235_valid_reg;
  assign line_236_clock = clock;
  assign line_236_reset = reset;
  assign line_236_valid = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ^ line_236_valid_reg;
  assign line_237_clock = clock;
  assign line_237_reset = reset;
  assign line_237_valid = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ^ line_237_valid_reg;
  assign line_238_clock = clock;
  assign line_238_reset = reset;
  assign line_238_valid = 5'ha == io_in_0_bits_ctrl_rfSrc1 ^ line_238_valid_reg;
  assign line_239_clock = clock;
  assign line_239_reset = reset;
  assign line_239_valid = 5'hb == io_in_0_bits_ctrl_rfSrc1 ^ line_239_valid_reg;
  assign line_240_clock = clock;
  assign line_240_reset = reset;
  assign line_240_valid = 5'hc == io_in_0_bits_ctrl_rfSrc1 ^ line_240_valid_reg;
  assign line_241_clock = clock;
  assign line_241_reset = reset;
  assign line_241_valid = 5'hd == io_in_0_bits_ctrl_rfSrc1 ^ line_241_valid_reg;
  assign line_242_clock = clock;
  assign line_242_reset = reset;
  assign line_242_valid = 5'he == io_in_0_bits_ctrl_rfSrc1 ^ line_242_valid_reg;
  assign line_243_clock = clock;
  assign line_243_reset = reset;
  assign line_243_valid = 5'hf == io_in_0_bits_ctrl_rfSrc1 ^ line_243_valid_reg;
  assign line_244_clock = clock;
  assign line_244_reset = reset;
  assign line_244_valid = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ^ line_244_valid_reg;
  assign line_245_clock = clock;
  assign line_245_reset = reset;
  assign line_245_valid = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ^ line_245_valid_reg;
  assign line_246_clock = clock;
  assign line_246_reset = reset;
  assign line_246_valid = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ^ line_246_valid_reg;
  assign line_247_clock = clock;
  assign line_247_reset = reset;
  assign line_247_valid = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ^ line_247_valid_reg;
  assign line_248_clock = clock;
  assign line_248_reset = reset;
  assign line_248_valid = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ^ line_248_valid_reg;
  assign line_249_clock = clock;
  assign line_249_reset = reset;
  assign line_249_valid = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ^ line_249_valid_reg;
  assign line_250_clock = clock;
  assign line_250_reset = reset;
  assign line_250_valid = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ^ line_250_valid_reg;
  assign line_251_clock = clock;
  assign line_251_reset = reset;
  assign line_251_valid = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ^ line_251_valid_reg;
  assign line_252_clock = clock;
  assign line_252_reset = reset;
  assign line_252_valid = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ^ line_252_valid_reg;
  assign line_253_clock = clock;
  assign line_253_reset = reset;
  assign line_253_valid = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ^ line_253_valid_reg;
  assign line_254_clock = clock;
  assign line_254_reset = reset;
  assign line_254_valid = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ^ line_254_valid_reg;
  assign line_255_clock = clock;
  assign line_255_reset = reset;
  assign line_255_valid = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ^ line_255_valid_reg;
  assign line_256_clock = clock;
  assign line_256_reset = reset;
  assign line_256_valid = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ^ line_256_valid_reg;
  assign line_257_clock = clock;
  assign line_257_reset = reset;
  assign line_257_valid = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ^ line_257_valid_reg;
  assign line_258_clock = clock;
  assign line_258_reset = reset;
  assign line_258_valid = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ^ line_258_valid_reg;
  assign line_259_clock = clock;
  assign line_259_reset = reset;
  assign line_259_valid = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ^ line_259_valid_reg;
  assign line_260_clock = clock;
  assign line_260_reset = reset;
  assign line_260_valid = 5'h0 == io_in_0_bits_ctrl_rfSrc2 ^ line_260_valid_reg;
  assign line_261_clock = clock;
  assign line_261_reset = reset;
  assign line_261_valid = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ^ line_261_valid_reg;
  assign line_262_clock = clock;
  assign line_262_reset = reset;
  assign line_262_valid = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ^ line_262_valid_reg;
  assign line_263_clock = clock;
  assign line_263_reset = reset;
  assign line_263_valid = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ^ line_263_valid_reg;
  assign line_264_clock = clock;
  assign line_264_reset = reset;
  assign line_264_valid = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ^ line_264_valid_reg;
  assign line_265_clock = clock;
  assign line_265_reset = reset;
  assign line_265_valid = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ^ line_265_valid_reg;
  assign line_266_clock = clock;
  assign line_266_reset = reset;
  assign line_266_valid = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ^ line_266_valid_reg;
  assign line_267_clock = clock;
  assign line_267_reset = reset;
  assign line_267_valid = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ^ line_267_valid_reg;
  assign line_268_clock = clock;
  assign line_268_reset = reset;
  assign line_268_valid = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ^ line_268_valid_reg;
  assign line_269_clock = clock;
  assign line_269_reset = reset;
  assign line_269_valid = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ^ line_269_valid_reg;
  assign line_270_clock = clock;
  assign line_270_reset = reset;
  assign line_270_valid = 5'ha == io_in_0_bits_ctrl_rfSrc2 ^ line_270_valid_reg;
  assign line_271_clock = clock;
  assign line_271_reset = reset;
  assign line_271_valid = 5'hb == io_in_0_bits_ctrl_rfSrc2 ^ line_271_valid_reg;
  assign line_272_clock = clock;
  assign line_272_reset = reset;
  assign line_272_valid = 5'hc == io_in_0_bits_ctrl_rfSrc2 ^ line_272_valid_reg;
  assign line_273_clock = clock;
  assign line_273_reset = reset;
  assign line_273_valid = 5'hd == io_in_0_bits_ctrl_rfSrc2 ^ line_273_valid_reg;
  assign line_274_clock = clock;
  assign line_274_reset = reset;
  assign line_274_valid = 5'he == io_in_0_bits_ctrl_rfSrc2 ^ line_274_valid_reg;
  assign line_275_clock = clock;
  assign line_275_reset = reset;
  assign line_275_valid = 5'hf == io_in_0_bits_ctrl_rfSrc2 ^ line_275_valid_reg;
  assign line_276_clock = clock;
  assign line_276_reset = reset;
  assign line_276_valid = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ^ line_276_valid_reg;
  assign line_277_clock = clock;
  assign line_277_reset = reset;
  assign line_277_valid = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ^ line_277_valid_reg;
  assign line_278_clock = clock;
  assign line_278_reset = reset;
  assign line_278_valid = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ^ line_278_valid_reg;
  assign line_279_clock = clock;
  assign line_279_reset = reset;
  assign line_279_valid = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ^ line_279_valid_reg;
  assign line_280_clock = clock;
  assign line_280_reset = reset;
  assign line_280_valid = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ^ line_280_valid_reg;
  assign line_281_clock = clock;
  assign line_281_reset = reset;
  assign line_281_valid = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ^ line_281_valid_reg;
  assign line_282_clock = clock;
  assign line_282_reset = reset;
  assign line_282_valid = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ^ line_282_valid_reg;
  assign line_283_clock = clock;
  assign line_283_reset = reset;
  assign line_283_valid = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ^ line_283_valid_reg;
  assign line_284_clock = clock;
  assign line_284_reset = reset;
  assign line_284_valid = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ^ line_284_valid_reg;
  assign line_285_clock = clock;
  assign line_285_reset = reset;
  assign line_285_valid = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ^ line_285_valid_reg;
  assign line_286_clock = clock;
  assign line_286_reset = reset;
  assign line_286_valid = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ^ line_286_valid_reg;
  assign line_287_clock = clock;
  assign line_287_reset = reset;
  assign line_287_valid = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ^ line_287_valid_reg;
  assign line_288_clock = clock;
  assign line_288_reset = reset;
  assign line_288_valid = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ^ line_288_valid_reg;
  assign line_289_clock = clock;
  assign line_289_reset = reset;
  assign line_289_valid = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ^ line_289_valid_reg;
  assign line_290_clock = clock;
  assign line_290_reset = reset;
  assign line_290_valid = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ^ line_290_valid_reg;
  assign line_291_clock = clock;
  assign line_291_reset = reset;
  assign line_291_valid = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ^ line_291_valid_reg;
  assign line_292_clock = clock;
  assign line_292_reset = reset;
  assign line_292_valid = io_wb_rfWen ^ line_292_valid_reg;
  assign line_293_clock = clock;
  assign line_293_reset = reset;
  assign line_293_valid = 5'h0 == io_wb_rfDest ^ line_293_valid_reg;
  assign line_294_clock = clock;
  assign line_294_reset = reset;
  assign line_294_valid = 5'h1 == io_wb_rfDest ^ line_294_valid_reg;
  assign line_295_clock = clock;
  assign line_295_reset = reset;
  assign line_295_valid = 5'h2 == io_wb_rfDest ^ line_295_valid_reg;
  assign line_296_clock = clock;
  assign line_296_reset = reset;
  assign line_296_valid = 5'h3 == io_wb_rfDest ^ line_296_valid_reg;
  assign line_297_clock = clock;
  assign line_297_reset = reset;
  assign line_297_valid = 5'h4 == io_wb_rfDest ^ line_297_valid_reg;
  assign line_298_clock = clock;
  assign line_298_reset = reset;
  assign line_298_valid = 5'h5 == io_wb_rfDest ^ line_298_valid_reg;
  assign line_299_clock = clock;
  assign line_299_reset = reset;
  assign line_299_valid = 5'h6 == io_wb_rfDest ^ line_299_valid_reg;
  assign line_300_clock = clock;
  assign line_300_reset = reset;
  assign line_300_valid = 5'h7 == io_wb_rfDest ^ line_300_valid_reg;
  assign line_301_clock = clock;
  assign line_301_reset = reset;
  assign line_301_valid = 5'h8 == io_wb_rfDest ^ line_301_valid_reg;
  assign line_302_clock = clock;
  assign line_302_reset = reset;
  assign line_302_valid = 5'h9 == io_wb_rfDest ^ line_302_valid_reg;
  assign line_303_clock = clock;
  assign line_303_reset = reset;
  assign line_303_valid = 5'ha == io_wb_rfDest ^ line_303_valid_reg;
  assign line_304_clock = clock;
  assign line_304_reset = reset;
  assign line_304_valid = 5'hb == io_wb_rfDest ^ line_304_valid_reg;
  assign line_305_clock = clock;
  assign line_305_reset = reset;
  assign line_305_valid = 5'hc == io_wb_rfDest ^ line_305_valid_reg;
  assign line_306_clock = clock;
  assign line_306_reset = reset;
  assign line_306_valid = 5'hd == io_wb_rfDest ^ line_306_valid_reg;
  assign line_307_clock = clock;
  assign line_307_reset = reset;
  assign line_307_valid = 5'he == io_wb_rfDest ^ line_307_valid_reg;
  assign line_308_clock = clock;
  assign line_308_reset = reset;
  assign line_308_valid = 5'hf == io_wb_rfDest ^ line_308_valid_reg;
  assign line_309_clock = clock;
  assign line_309_reset = reset;
  assign line_309_valid = 5'h10 == io_wb_rfDest ^ line_309_valid_reg;
  assign line_310_clock = clock;
  assign line_310_reset = reset;
  assign line_310_valid = 5'h11 == io_wb_rfDest ^ line_310_valid_reg;
  assign line_311_clock = clock;
  assign line_311_reset = reset;
  assign line_311_valid = 5'h12 == io_wb_rfDest ^ line_311_valid_reg;
  assign line_312_clock = clock;
  assign line_312_reset = reset;
  assign line_312_valid = 5'h13 == io_wb_rfDest ^ line_312_valid_reg;
  assign line_313_clock = clock;
  assign line_313_reset = reset;
  assign line_313_valid = 5'h14 == io_wb_rfDest ^ line_313_valid_reg;
  assign line_314_clock = clock;
  assign line_314_reset = reset;
  assign line_314_valid = 5'h15 == io_wb_rfDest ^ line_314_valid_reg;
  assign line_315_clock = clock;
  assign line_315_reset = reset;
  assign line_315_valid = 5'h16 == io_wb_rfDest ^ line_315_valid_reg;
  assign line_316_clock = clock;
  assign line_316_reset = reset;
  assign line_316_valid = 5'h17 == io_wb_rfDest ^ line_316_valid_reg;
  assign line_317_clock = clock;
  assign line_317_reset = reset;
  assign line_317_valid = 5'h18 == io_wb_rfDest ^ line_317_valid_reg;
  assign line_318_clock = clock;
  assign line_318_reset = reset;
  assign line_318_valid = 5'h19 == io_wb_rfDest ^ line_318_valid_reg;
  assign line_319_clock = clock;
  assign line_319_reset = reset;
  assign line_319_valid = 5'h1a == io_wb_rfDest ^ line_319_valid_reg;
  assign line_320_clock = clock;
  assign line_320_reset = reset;
  assign line_320_valid = 5'h1b == io_wb_rfDest ^ line_320_valid_reg;
  assign line_321_clock = clock;
  assign line_321_reset = reset;
  assign line_321_valid = 5'h1c == io_wb_rfDest ^ line_321_valid_reg;
  assign line_322_clock = clock;
  assign line_322_reset = reset;
  assign line_322_valid = 5'h1d == io_wb_rfDest ^ line_322_valid_reg;
  assign line_323_clock = clock;
  assign line_323_reset = reset;
  assign line_323_valid = 5'h1e == io_wb_rfDest ^ line_323_valid_reg;
  assign line_324_clock = clock;
  assign line_324_reset = reset;
  assign line_324_valid = 5'h1f == io_wb_rfDest ^ line_324_valid_reg;
  assign line_325_clock = clock;
  assign line_325_reset = reset;
  assign line_325_valid = io_flush ^ line_325_valid_reg;
  assign line_326_clock = clock;
  assign line_326_reset = reset;
  assign line_326_valid = io_flush ^ line_326_valid_reg;
  assign io_in_0_ready = ~io_in_0_valid | _isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[src/main/scala/nutcore/backend/seq/ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_data_src1 = _io_out_bits_data_src1_T_17 | _io_out_bits_data_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_src2 = _io_out_bits_data_src2_T_15 | _io_out_bits_data_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/ISU.scala 75:25]
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_value_1 = rf_1; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_2 = rf_2; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_3 = rf_3; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_4 = rf_4; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_5 = rf_5; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_6 = rf_6; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_7 = rf_7; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_8 = rf_8; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_9 = rf_9; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_10 = rf_10; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_11 = rf_11; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_12 = rf_12; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_13 = rf_13; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_14 = rf_14; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_15 = rf_15; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_16 = rf_16; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_17 = rf_17; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_18 = rf_18; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_19 = rf_19; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_20 = rf_20; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_21 = rf_21; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_22 = rf_22; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_23 = rf_23; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_24 = rf_24; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_25 = rf_25; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_26 = rf_26; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_27 = rf_27; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_28 = rf_28; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_29 = rf_29; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_30 = rf_30; // @[src/main/scala/nutcore/RF.scala 33:36]
  assign difftest_module_io_bits_value_31 = rf_31; // @[src/main/scala/nutcore/RF.scala 33:36]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 38:21]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 38:21]
    end else if (io_flush) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 88:19]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 46:10]
    end else begin
      busy <= _busy_T_9; // @[src/main/scala/nutcore/RF.scala 46:10]
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h0 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_0 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_1 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_1 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_2 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h2 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_2 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_3 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h3 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_3 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_4 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h4 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_4 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_5 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h5 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_5 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_6 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h6 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_6 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_7 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h7 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_7 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_8 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h8 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_8 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_9 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h9 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_9 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_10 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'ha == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_10 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_11 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hb == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_11 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_12 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hc == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_12 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_13 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hd == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_13 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_14 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'he == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_14 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_15 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hf == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_15 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_16 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h10 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_16 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_17 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h11 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_17 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_18 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h12 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_18 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_19 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h13 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_19 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_20 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h14 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_20 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_21 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h15 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_21 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_22 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h16 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_22 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_23 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h17 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_23 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_24 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h18 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_24 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_25 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h19 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_25 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_26 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1a == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_26 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_27 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1b == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_27 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_28 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1c == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_28 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_29 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1d == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_29 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_30 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1e == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_30 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 32:19]
      rf_31 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 32:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1f == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 34:50]
        rf_31 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 34:50]
      end
    end
    line_228_valid_reg <= 5'h0 == io_in_0_bits_ctrl_rfSrc1;
    line_229_valid_reg <= 5'h1 == io_in_0_bits_ctrl_rfSrc1;
    line_230_valid_reg <= 5'h2 == io_in_0_bits_ctrl_rfSrc1;
    line_231_valid_reg <= 5'h3 == io_in_0_bits_ctrl_rfSrc1;
    line_232_valid_reg <= 5'h4 == io_in_0_bits_ctrl_rfSrc1;
    line_233_valid_reg <= 5'h5 == io_in_0_bits_ctrl_rfSrc1;
    line_234_valid_reg <= 5'h6 == io_in_0_bits_ctrl_rfSrc1;
    line_235_valid_reg <= 5'h7 == io_in_0_bits_ctrl_rfSrc1;
    line_236_valid_reg <= 5'h8 == io_in_0_bits_ctrl_rfSrc1;
    line_237_valid_reg <= 5'h9 == io_in_0_bits_ctrl_rfSrc1;
    line_238_valid_reg <= 5'ha == io_in_0_bits_ctrl_rfSrc1;
    line_239_valid_reg <= 5'hb == io_in_0_bits_ctrl_rfSrc1;
    line_240_valid_reg <= 5'hc == io_in_0_bits_ctrl_rfSrc1;
    line_241_valid_reg <= 5'hd == io_in_0_bits_ctrl_rfSrc1;
    line_242_valid_reg <= 5'he == io_in_0_bits_ctrl_rfSrc1;
    line_243_valid_reg <= 5'hf == io_in_0_bits_ctrl_rfSrc1;
    line_244_valid_reg <= 5'h10 == io_in_0_bits_ctrl_rfSrc1;
    line_245_valid_reg <= 5'h11 == io_in_0_bits_ctrl_rfSrc1;
    line_246_valid_reg <= 5'h12 == io_in_0_bits_ctrl_rfSrc1;
    line_247_valid_reg <= 5'h13 == io_in_0_bits_ctrl_rfSrc1;
    line_248_valid_reg <= 5'h14 == io_in_0_bits_ctrl_rfSrc1;
    line_249_valid_reg <= 5'h15 == io_in_0_bits_ctrl_rfSrc1;
    line_250_valid_reg <= 5'h16 == io_in_0_bits_ctrl_rfSrc1;
    line_251_valid_reg <= 5'h17 == io_in_0_bits_ctrl_rfSrc1;
    line_252_valid_reg <= 5'h18 == io_in_0_bits_ctrl_rfSrc1;
    line_253_valid_reg <= 5'h19 == io_in_0_bits_ctrl_rfSrc1;
    line_254_valid_reg <= 5'h1a == io_in_0_bits_ctrl_rfSrc1;
    line_255_valid_reg <= 5'h1b == io_in_0_bits_ctrl_rfSrc1;
    line_256_valid_reg <= 5'h1c == io_in_0_bits_ctrl_rfSrc1;
    line_257_valid_reg <= 5'h1d == io_in_0_bits_ctrl_rfSrc1;
    line_258_valid_reg <= 5'h1e == io_in_0_bits_ctrl_rfSrc1;
    line_259_valid_reg <= 5'h1f == io_in_0_bits_ctrl_rfSrc1;
    line_260_valid_reg <= 5'h0 == io_in_0_bits_ctrl_rfSrc2;
    line_261_valid_reg <= 5'h1 == io_in_0_bits_ctrl_rfSrc2;
    line_262_valid_reg <= 5'h2 == io_in_0_bits_ctrl_rfSrc2;
    line_263_valid_reg <= 5'h3 == io_in_0_bits_ctrl_rfSrc2;
    line_264_valid_reg <= 5'h4 == io_in_0_bits_ctrl_rfSrc2;
    line_265_valid_reg <= 5'h5 == io_in_0_bits_ctrl_rfSrc2;
    line_266_valid_reg <= 5'h6 == io_in_0_bits_ctrl_rfSrc2;
    line_267_valid_reg <= 5'h7 == io_in_0_bits_ctrl_rfSrc2;
    line_268_valid_reg <= 5'h8 == io_in_0_bits_ctrl_rfSrc2;
    line_269_valid_reg <= 5'h9 == io_in_0_bits_ctrl_rfSrc2;
    line_270_valid_reg <= 5'ha == io_in_0_bits_ctrl_rfSrc2;
    line_271_valid_reg <= 5'hb == io_in_0_bits_ctrl_rfSrc2;
    line_272_valid_reg <= 5'hc == io_in_0_bits_ctrl_rfSrc2;
    line_273_valid_reg <= 5'hd == io_in_0_bits_ctrl_rfSrc2;
    line_274_valid_reg <= 5'he == io_in_0_bits_ctrl_rfSrc2;
    line_275_valid_reg <= 5'hf == io_in_0_bits_ctrl_rfSrc2;
    line_276_valid_reg <= 5'h10 == io_in_0_bits_ctrl_rfSrc2;
    line_277_valid_reg <= 5'h11 == io_in_0_bits_ctrl_rfSrc2;
    line_278_valid_reg <= 5'h12 == io_in_0_bits_ctrl_rfSrc2;
    line_279_valid_reg <= 5'h13 == io_in_0_bits_ctrl_rfSrc2;
    line_280_valid_reg <= 5'h14 == io_in_0_bits_ctrl_rfSrc2;
    line_281_valid_reg <= 5'h15 == io_in_0_bits_ctrl_rfSrc2;
    line_282_valid_reg <= 5'h16 == io_in_0_bits_ctrl_rfSrc2;
    line_283_valid_reg <= 5'h17 == io_in_0_bits_ctrl_rfSrc2;
    line_284_valid_reg <= 5'h18 == io_in_0_bits_ctrl_rfSrc2;
    line_285_valid_reg <= 5'h19 == io_in_0_bits_ctrl_rfSrc2;
    line_286_valid_reg <= 5'h1a == io_in_0_bits_ctrl_rfSrc2;
    line_287_valid_reg <= 5'h1b == io_in_0_bits_ctrl_rfSrc2;
    line_288_valid_reg <= 5'h1c == io_in_0_bits_ctrl_rfSrc2;
    line_289_valid_reg <= 5'h1d == io_in_0_bits_ctrl_rfSrc2;
    line_290_valid_reg <= 5'h1e == io_in_0_bits_ctrl_rfSrc2;
    line_291_valid_reg <= 5'h1f == io_in_0_bits_ctrl_rfSrc2;
    line_292_valid_reg <= io_wb_rfWen;
    line_293_valid_reg <= 5'h0 == io_wb_rfDest;
    line_294_valid_reg <= 5'h1 == io_wb_rfDest;
    line_295_valid_reg <= 5'h2 == io_wb_rfDest;
    line_296_valid_reg <= 5'h3 == io_wb_rfDest;
    line_297_valid_reg <= 5'h4 == io_wb_rfDest;
    line_298_valid_reg <= 5'h5 == io_wb_rfDest;
    line_299_valid_reg <= 5'h6 == io_wb_rfDest;
    line_300_valid_reg <= 5'h7 == io_wb_rfDest;
    line_301_valid_reg <= 5'h8 == io_wb_rfDest;
    line_302_valid_reg <= 5'h9 == io_wb_rfDest;
    line_303_valid_reg <= 5'ha == io_wb_rfDest;
    line_304_valid_reg <= 5'hb == io_wb_rfDest;
    line_305_valid_reg <= 5'hc == io_wb_rfDest;
    line_306_valid_reg <= 5'hd == io_wb_rfDest;
    line_307_valid_reg <= 5'he == io_wb_rfDest;
    line_308_valid_reg <= 5'hf == io_wb_rfDest;
    line_309_valid_reg <= 5'h10 == io_wb_rfDest;
    line_310_valid_reg <= 5'h11 == io_wb_rfDest;
    line_311_valid_reg <= 5'h12 == io_wb_rfDest;
    line_312_valid_reg <= 5'h13 == io_wb_rfDest;
    line_313_valid_reg <= 5'h14 == io_wb_rfDest;
    line_314_valid_reg <= 5'h15 == io_wb_rfDest;
    line_315_valid_reg <= 5'h16 == io_wb_rfDest;
    line_316_valid_reg <= 5'h17 == io_wb_rfDest;
    line_317_valid_reg <= 5'h18 == io_wb_rfDest;
    line_318_valid_reg <= 5'h19 == io_wb_rfDest;
    line_319_valid_reg <= 5'h1a == io_wb_rfDest;
    line_320_valid_reg <= 5'h1b == io_wb_rfDest;
    line_321_valid_reg <= 5'h1c == io_wb_rfDest;
    line_322_valid_reg <= 5'h1d == io_wb_rfDest;
    line_323_valid_reg <= 5'h1e == io_wb_rfDest;
    line_324_valid_reg <= 5'h1f == io_wb_rfDest;
    line_325_valid_reg <= io_flush;
    line_326_valid_reg <= io_flush;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  rf_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  rf_31 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  line_228_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_229_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_230_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_231_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_232_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_233_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_234_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_235_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_236_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_237_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_238_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_239_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_240_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_241_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_242_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_243_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_244_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_245_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_246_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_247_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_248_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_249_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_250_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_251_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_252_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_253_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_254_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_255_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_256_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_257_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_258_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_259_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_260_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_261_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_262_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_263_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_264_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_265_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_266_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_267_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_268_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_269_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_270_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_271_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_272_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_273_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_274_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_275_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_276_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_277_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_278_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_279_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_280_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_281_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_282_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_283_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_284_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_285_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_286_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_287_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_288_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_289_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_290_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_291_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_292_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_293_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_294_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_295_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_296_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_297_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_298_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_299_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_300_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_301_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_302_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_303_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_304_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_305_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_306_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_307_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_308_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_309_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_310_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_311_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_312_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_313_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_314_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_315_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_316_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_317_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_318_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_319_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_320_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_321_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_322_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_323_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_324_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_325_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_326_valid_reg = _RAND_131[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (5'h0 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h2 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h3 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h4 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h5 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h6 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h7 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h8 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h9 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'ha == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'hb == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'hc == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'hd == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'he == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'hf == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h10 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h11 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h12 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h13 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h14 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h15 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h16 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h17 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h18 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h19 == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1a == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1b == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1c == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1d == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1e == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h1f == io_in_0_bits_ctrl_rfSrc1) begin
      cover(1'h1);
    end
    //
    if (5'h0 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h2 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h3 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h4 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h5 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h6 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h7 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h8 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h9 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'ha == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'hb == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'hc == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'hd == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'he == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'hf == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h10 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h11 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h12 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h13 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h14 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h15 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h16 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h17 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h18 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h19 == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1a == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1b == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1c == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1d == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1e == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (5'h1f == io_in_0_bits_ctrl_rfSrc2) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_64) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_65) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_66) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_67) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_68) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_69) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_70) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_71) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_72) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_73) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_74) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_75) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_76) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_77) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_78) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_79) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_80) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_81) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_82) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_83) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_84) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_85) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_86) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_87) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_88) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_89) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_90) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_91) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_92) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_93) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_94) begin
      cover(1'h1);
    end
    //
    if (io_wb_rfWen & _GEN_95) begin
      cover(1'h1);
    end
    //
    if (io_flush) begin
      cover(1'h1);
    end
    //
    if (~io_flush) begin
      cover(1'h1);
    end
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pnpc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [3:0]  io_cfIn_brIdx, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_offset, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_iVmEnable, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_jumpIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_jumpIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_jumpIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output        REG_0_actualTaken,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 89:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:39]
  wire [63:0] _adderRes_T_1 = io_in_bits_src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:33]
  wire [64:0] _adderRes_T_2 = io_in_bits_src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:24]
  wire [64:0] _GEN_9 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_9; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 91:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 92:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/ALU.scala 93:28]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  shsrc1_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _shsrc1_T_4 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _shsrc1_T_5 = {_shsrc1_T_4,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _shsrc1_T_7 = 7'h25 == io_in_bits_func ? _shsrc1_T_2 : io_in_bits_src1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:18]
  wire [126:0] _GEN_8 = {{63'd0}, shsrc1}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [126:0] _res_T_1 = _GEN_8 << shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 105:32]
  wire [63:0] _res_T_6 = io_in_bits_src1 | io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:30]
  wire [63:0] _res_T_7 = io_in_bits_src1 & io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 107:30]
  wire [63:0] _res_T_8 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:32]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:49]
  wire [64:0] _res_T_12 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_1[63:0]} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_3} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_4} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_5} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_7} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  aluRes_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _aluRes_T_2 = aluRes_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _aluRes_T_3 = {_aluRes_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _aluRes_T_3} : res; // @[src/main/scala/nutcore/backend/fu/ALU.scala 110:19]
  wire  _T_1 = ~(|xorRes); // @[src/main/scala/nutcore/backend/fu/ALU.scala 113:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _taken_T_1 = 2'h0 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_2 = 2'h2 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_3 = 2'h3 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_8 = _taken_T_1 & _T_1 | _taken_T_2 & slt | _taken_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  taken = _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
  wire  target_signBit = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _target_T = target_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _target_T_1 = {_target_T,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _target_T_3 = _target_T_1 + io_offset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:56]
  wire [63:0] _target_T_5 = {adderRes[63:1],1'h0}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:72]
  wire [63:0] target = isBranch ? _target_T_3 : _target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
  wire  _predictWrong_T_1 = ~taken & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
  wire  _T_8 = ~reset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
  wire  line_327_clock;
  wire  line_327_reset;
  wire  line_327_valid;
  reg  line_327_valid_reg;
  wire  _T_9 = ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
  wire  line_328_clock;
  wire  line_328_reset;
  wire  line_328_valid;
  reg  line_328_valid_reg;
  wire  _T_12 = ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 125:55]
  wire [38:0] _io_redirect_target_T_3 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:71]
  wire [38:0] _io_redirect_target_T_5 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:89]
  wire [38:0] _io_redirect_target_T_6 = isRVC ? _io_redirect_target_T_3 : _io_redirect_target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:52]
  wire [63:0] _io_redirect_target_T_7 = _predictWrong_T_1 ? {{25'd0}, _io_redirect_target_T_6} : target; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:28]
  wire  _io_redirect_valid_T = io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:30]
  wire  _io_redirect_valid_T_1 = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  wire [63:0] _io_out_bits_T_4 = _target_T_1 + 64'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:71]
  wire [63:0] _io_out_bits_T_8 = _target_T_1 + 64'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:108]
  wire [63:0] _io_out_bits_T_9 = _T_12 ? _io_out_bits_T_4 : _io_out_bits_T_8; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:32]
  wire [64:0] _io_out_bits_T_10 = isBru ? {{1'd0}, _io_out_bits_T_9} : aluRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:21]
  reg  hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
  wire  addrNotLegal_signBit = target[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,target[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  addrNotLegal = io_iVmEnable ? target != _addrNotLegal_T_2 : |target[63:39]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 139:25]
  wire  isIllegalJumpAddr = io_redirect_valid & ~isBranch & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/ALU.scala 140:58]
  wire  line_329_clock;
  wire  line_329_reset;
  wire  line_329_valid;
  reg  line_329_valid_reg;
  wire  line_330_clock;
  wire  line_330_reset;
  wire  line_330_valid;
  reg  line_330_valid_reg;
  wire  _T_15 = io_jumpIsIllegal_ready & io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_331_clock;
  wire  line_331_reset;
  wire  line_331_valid;
  reg  line_331_valid_reg;
  wire  _GEN_6 = _T_15 ? 1'h0 : hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:38 144:24 138:35]
  wire  _GEN_7 = isIllegalJumpAddr | _GEN_6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 141:28 142:24]
  reg [63:0] io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
  wire  line_332_clock;
  wire  line_332_reset;
  wire  line_332_valid;
  reg  line_332_valid_reg;
  wire  _T_21 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:180]
  wire  _T_22 = io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:214]
  wire  _T_23 = io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:239]
  wire  _T_32 = 7'h5c == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_33 = 7'h5e == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_34 = 7'h58 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_35 = 7'h5a == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [1:0] _T_43 = _T_33 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_45 = _T_35 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_10 = {{1'd0}, _T_32}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_52 = _GEN_10 | _T_43; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_11 = {{1'd0}, _T_34}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_53 = _T_52 | _GEN_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [6:0] REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [1:0] REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  right = _io_redirect_valid_T & ~predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:32]
  wire  _T_55 = right & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:33]
  wire  _T_56 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 179:33]
  wire  _T_60 = _T_56 & io_cfIn_pc[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:45]
  wire  _T_61 = _T_56 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:73]
  wire  _T_67 = _T_60 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 181:73]
  wire  _T_71 = _T_56 & io_cfIn_pc[2:0] == 3'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:45]
  wire  _T_72 = _T_56 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:73]
  wire  _T_78 = _T_71 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 183:73]
  wire  _T_82 = _T_56 & io_cfIn_pc[2:0] == 3'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:45]
  wire  _T_83 = _T_56 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:73]
  wire  _T_89 = _T_82 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 185:73]
  wire  _T_93 = _T_56 & io_cfIn_pc[2:0] == 3'h6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:45]
  wire  _T_94 = _T_56 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:73]
  wire  _T_100 = _T_93 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 187:73]
  wire  _T_104 = right & _T_21; // @[src/main/scala/nutcore/backend/fu/ALU.scala 188:33]
  wire  _T_108 = _io_redirect_valid_T_1 & _T_21; // @[src/main/scala/nutcore/backend/fu/ALU.scala 189:33]
  wire  _T_110 = right & _T_22; // @[src/main/scala/nutcore/backend/fu/ALU.scala 190:33]
  wire  _T_112 = _io_redirect_valid_T_1 & _T_22; // @[src/main/scala/nutcore/backend/fu/ALU.scala 191:33]
  wire  _T_114 = right & _T_23; // @[src/main/scala/nutcore/backend/fu/ALU.scala 192:33]
  wire  _T_116 = _io_redirect_valid_T_1 & _T_23; // @[src/main/scala/nutcore/backend/fu/ALU.scala 193:33]
  GEN_w1_line #(.COVER_INDEX(327)) line_327 (
    .clock(line_327_clock),
    .reset(line_327_reset),
    .valid(line_327_valid)
  );
  GEN_w1_line #(.COVER_INDEX(328)) line_328 (
    .clock(line_328_clock),
    .reset(line_328_reset),
    .valid(line_328_valid)
  );
  GEN_w1_line #(.COVER_INDEX(329)) line_329 (
    .clock(line_329_clock),
    .reset(line_329_reset),
    .valid(line_329_valid)
  );
  GEN_w1_line #(.COVER_INDEX(330)) line_330 (
    .clock(line_330_clock),
    .reset(line_330_reset),
    .valid(line_330_valid)
  );
  GEN_w1_line #(.COVER_INDEX(331)) line_331 (
    .clock(line_331_clock),
    .reset(line_331_reset),
    .valid(line_331_valid)
  );
  GEN_w1_line #(.COVER_INDEX(332)) line_332 (
    .clock(line_332_clock),
    .reset(line_332_reset),
    .valid(line_332_valid)
  );
  assign line_327_clock = clock;
  assign line_327_reset = reset;
  assign line_327_valid = _T_8 ^ line_327_valid_reg;
  assign line_328_clock = clock;
  assign line_328_reset = reset;
  assign line_328_valid = _T_9 ^ line_328_valid_reg;
  assign line_329_clock = clock;
  assign line_329_reset = reset;
  assign line_329_valid = isIllegalJumpAddr ^ line_329_valid_reg;
  assign line_330_clock = clock;
  assign line_330_reset = reset;
  assign line_330_valid = isIllegalJumpAddr ^ line_330_valid_reg;
  assign line_331_clock = clock;
  assign line_331_reset = reset;
  assign line_331_valid = _T_15 ^ line_331_valid_reg;
  assign line_332_clock = clock;
  assign line_332_reset = reset;
  assign line_332_valid = isIllegalJumpAddr ^ line_332_valid_reg;
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 161:16]
  assign io_out_bits = _io_out_bits_T_10[63:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:15]
  assign io_redirect_target = _io_redirect_target_T_7[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:22]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  assign io_jumpIsIllegal_valid = hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 146:26]
  assign io_jumpIsIllegal_bits = io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:25]
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_actualTaken = REG_actualTaken;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  always @(posedge clock) begin
    line_327_valid_reg <= _T_8;
    line_328_valid_reg <= _T_9;
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
      hasIllegalJumpAddr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
    end else begin
      hasIllegalJumpAddr <= _GEN_7;
    end
    line_329_valid_reg <= isIllegalJumpAddr;
    line_330_valid_reg <= isIllegalJumpAddr;
    line_331_valid_reg <= _T_15;
    if (isIllegalJumpAddr) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
      if (isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
        io_jumpIsIllegal_bits_r <= _target_T_3;
      end else begin
        io_jumpIsIllegal_bits_r <= _target_T_5;
      end
    end
    line_332_valid_reg <= isIllegalJumpAddr;
    REG_valid <= io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 164:31]
    REG_pc <= io_cfIn_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 165:19]
    if (~taken & isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= target[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 167:29]
    REG_actualTaken <= _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
    REG_fuOpType <= io_in_bits_func; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 169:25]
    REG_btbType <= _T_53 | _T_45; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:124 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_327_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_328_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hasIllegalJumpAddr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_329_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_330_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_331_valid_reg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  io_jumpIsIllegal_bits_r = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  line_332_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG_valid = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  REG_pc = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  REG_actualTarget = _RAND_11[38:0];
  _RAND_12 = {1{`RANDOM}};
  REG_actualTaken = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_fuOpType = _RAND_13[6:0];
  _RAND_14 = {1{`RANDOM}};
  REG_btbType = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  REG_isRVC = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_8) begin
      cover(1'h1);
    end
    //
    if (_T_8 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
    end
    //
    if (isIllegalJumpAddr) begin
      cover(1'h1);
    end
    //
    if (~isIllegalJumpAddr) begin
      cover(1'h1);
    end
    //
    if (~isIllegalJumpAddr & _T_15) begin
      cover(1'h1);
    end
    //
    if (isIllegalJumpAddr) begin
      cover(1'h1);
    end
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_resp_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         DTLBPF,
  input         scIsSuccess_0,
  input         vmEnable_0,
  input         ISAMO2,
  input         DTLBFINISH,
  input         DTLBAF
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  _io_vaddr_T = io__in_ready & io__in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_333_clock;
  wire  line_333_reset;
  wire  line_333_valid;
  reg  line_333_valid_reg;
  reg [63:0] addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 423:23]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 424:30]
  reg [1:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
  wire [5:0] vaddrPF_lo_lo = {io__vaddr[58] != io__vaddr[38],io__vaddr[59] != io__vaddr[38],io__vaddr[60] != io__vaddr[
    38],io__vaddr[61] != io__vaddr[38],io__vaddr[62] != io__vaddr[38],io__vaddr[63] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [11:0] vaddrPF_lo = {io__vaddr[52] != io__vaddr[38],io__vaddr[53] != io__vaddr[38],io__vaddr[54] != io__vaddr[38]
    ,io__vaddr[55] != io__vaddr[38],io__vaddr[56] != io__vaddr[38],io__vaddr[57] != io__vaddr[38],vaddrPF_lo_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [5:0] vaddrPF_hi_lo = {io__vaddr[46] != io__vaddr[38],io__vaddr[47] != io__vaddr[38],io__vaddr[48] != io__vaddr[
    38],io__vaddr[49] != io__vaddr[38],io__vaddr[50] != io__vaddr[38],io__vaddr[51] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [24:0] _vaddrPF_T_76 = {io__vaddr[39] != io__vaddr[38],io__vaddr[40] != io__vaddr[38],io__vaddr[41] != io__vaddr[
    38],io__vaddr[42] != io__vaddr[38],io__vaddr[43] != io__vaddr[38],io__vaddr[44] != io__vaddr[38],io__vaddr[45] !=
    io__vaddr[38],vaddrPF_hi_lo,vaddrPF_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire  vaddrPF = io__in_valid & vmEnable_0 & |_vaddrPF_T_76; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:37]
  wire  dtlbHasException = DTLBPF | DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 446:33]
  wire  _T = 2'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
  wire  line_334_clock;
  wire  line_334_reset;
  wire  line_334_valid;
  reg  line_334_valid_reg;
  wire  _T_1 = io__dmem_req_ready & io__dmem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_2 = _T_1 & vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:29]
  wire  line_335_clock;
  wire  line_335_reset;
  wire  line_335_valid;
  reg  line_335_valid_reg;
  wire  _T_4 = ~vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:32]
  wire  _T_5 = _T_1 & ~vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:29]
  wire  line_336_clock;
  wire  line_336_reset;
  wire  line_336_valid;
  reg  line_336_valid_reg;
  wire  line_337_clock;
  wire  line_337_reset;
  wire  line_337_valid;
  reg  line_337_valid_reg;
  wire  _T_6 = 2'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
  wire  line_338_clock;
  wire  line_338_reset;
  wire  line_338_valid;
  reg  line_338_valid_reg;
  wire  _T_9 = DTLBFINISH & (dtlbHasException | ~scIsSuccess_0); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 454:24]
  wire  line_339_clock;
  wire  line_339_reset;
  wire  line_339_valid;
  reg  line_339_valid_reg;
  wire [1:0] _GEN_20 = DTLBFINISH & (dtlbHasException | ~scIsSuccess_0) ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 454:{63,71}]
  wire  _T_12 = DTLBFINISH & ~dtlbHasException & scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:45]
  wire  line_340_clock;
  wire  line_340_reset;
  wire  line_340_valid;
  reg  line_340_valid_reg;
  wire  line_341_clock;
  wire  line_341_reset;
  wire  line_341_valid;
  reg  line_341_valid_reg;
  wire  _T_13 = 2'h2 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
  wire  line_342_clock;
  wire  line_342_reset;
  wire  line_342_valid;
  reg  line_342_valid_reg;
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_343_clock;
  wire  line_343_reset;
  wire  line_343_valid;
  reg  line_343_valid_reg;
  wire [1:0] _state_T = partialLoad ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 457:62]
  wire [1:0] _GEN_22 = _T_14 ? _state_T : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 457:{48,56}]
  wire  line_344_clock;
  wire  line_344_reset;
  wire  line_344_valid;
  reg  line_344_valid_reg;
  wire  _T_15 = 2'h3 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
  wire  line_345_clock;
  wire  line_345_reset;
  wire  line_345_valid;
  reg  line_345_valid_reg;
  wire [1:0] _GEN_23 = 2'h3 == state ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18 427:22 458:32]
  wire [63:0] _reqWdata_T_3 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]
    ,io__wdata[7:0],io__wdata[7:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 399:22]
  wire [63:0] _reqWdata_T_6 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 400:22]
  wire [63:0] _reqWdata_T_8 = {io__wdata[31:0],io__wdata[31:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 401:22]
  wire  _reqWdata_T_9 = 2'h0 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_10 = 2'h1 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_11 = 2'h2 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_12 = 2'h3 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _reqWdata_T_13 = _reqWdata_T_9 ? _reqWdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_14 = _reqWdata_T_10 ? _reqWdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_15 = _reqWdata_T_11 ? _reqWdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_16 = _reqWdata_T_12 ? io__wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_17 = _reqWdata_T_13 | _reqWdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_18 = _reqWdata_T_17 | _reqWdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_5 = _reqWdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_6 = _reqWdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_7 = _reqWdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_31 = {{1'd0}, _reqWdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_8 = _GEN_31 | _reqWmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_32 = {{2'd0}, _reqWmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_9 = _GEN_32 | _reqWmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_33 = {{4'd0}, _reqWmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_10 = _GEN_33 | _reqWmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_41 = {{7'd0}, _reqWmask_T_10}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire [14:0] reqWmask = _GEN_41 << io__in_bits_src1[2:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire  hasException = io__loadAccessFault | io__storeAccessFault | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 476:64]
  wire  _io_dmem_req_valid_T = state == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:37]
  wire  _io_out_valid_T_3 = state == 2'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 483:13]
  wire  _io_out_valid_T_6 = _T_14 & state == 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 484:22]
  wire  _io_out_valid_T_7 = partialLoad ? _io_out_valid_T_3 : _io_out_valid_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 482:8]
  reg [63:0] rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
  wire  _rdataSel64_T_9 = 3'h0 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_10 = 3'h1 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_11 = 3'h2 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_12 = 3'h3 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_13 = 3'h4 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_14 = 3'h5 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_15 = 3'h6 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_16 = 3'h7 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataSel64_T_17 = _rdataSel64_T_9 ? rdataLatch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdataSel64_T_18 = _rdataSel64_T_10 ? rdataLatch[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdataSel64_T_19 = _rdataSel64_T_11 ? rdataLatch[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdataSel64_T_20 = _rdataSel64_T_12 ? rdataLatch[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdataSel64_T_21 = _rdataSel64_T_13 ? rdataLatch[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdataSel64_T_22 = _rdataSel64_T_14 ? rdataLatch[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdataSel64_T_23 = _rdataSel64_T_15 ? rdataLatch[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdataSel64_T_24 = _rdataSel64_T_16 ? rdataLatch[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_34 = {{8'd0}, _rdataSel64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_25 = _rdataSel64_T_17 | _GEN_34; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_35 = {{16'd0}, _rdataSel64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_26 = _rdataSel64_T_25 | _GEN_35; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_36 = {{24'd0}, _rdataSel64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_27 = _rdataSel64_T_26 | _GEN_36; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_37 = {{32'd0}, _rdataSel64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_28 = _rdataSel64_T_27 | _GEN_37; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_38 = {{40'd0}, _rdataSel64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_29 = _rdataSel64_T_28 | _GEN_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_39 = {{48'd0}, _rdataSel64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_30 = _rdataSel64_T_29 | _GEN_39; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_40 = {{56'd0}, _rdataSel64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataSel64 = _rdataSel64_T_30 | _GEN_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdataPartialLoad_signBit = rdataSel64[7]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [55:0] _rdataPartialLoad_T_1 = rdataPartialLoad_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_2 = {_rdataPartialLoad_T_1,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_1 = rdataSel64[15]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [47:0] _rdataPartialLoad_T_4 = rdataPartialLoad_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_5 = {_rdataPartialLoad_T_4,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_2 = rdataSel64[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _rdataPartialLoad_T_7 = rdataPartialLoad_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_8 = {_rdataPartialLoad_T_7,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _rdataPartialLoad_T_10 = {56'h0,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_12 = {48'h0,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_14 = {32'h0,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdataPartialLoad_T_15 = 7'h0 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_16 = 7'h1 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_17 = 7'h2 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_18 = 7'h4 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_19 = 7'h5 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_20 = 7'h6 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataPartialLoad_T_21 = _rdataPartialLoad_T_15 ? _rdataPartialLoad_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_22 = _rdataPartialLoad_T_16 ? _rdataPartialLoad_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_23 = _rdataPartialLoad_T_17 ? _rdataPartialLoad_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_24 = _rdataPartialLoad_T_18 ? _rdataPartialLoad_T_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_25 = _rdataPartialLoad_T_19 ? _rdataPartialLoad_T_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_26 = _rdataPartialLoad_T_20 ? _rdataPartialLoad_T_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_27 = _rdataPartialLoad_T_21 | _rdataPartialLoad_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_28 = _rdataPartialLoad_T_27 | _rdataPartialLoad_T_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_29 = _rdataPartialLoad_T_28 | _rdataPartialLoad_T_24; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_30 = _rdataPartialLoad_T_29 | _rdataPartialLoad_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataPartialLoad = _rdataPartialLoad_T_30 | _rdataPartialLoad_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_loadAccessFault_T_1 = io__in_valid & _T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:32]
  wire  _io_loadAccessFault_T_7 = io__in_bits_src1 >= 64'h38000000 & io__in_bits_src1 < 64'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_10 = io__in_bits_src1 >= 64'h3c000000 & io__in_bits_src1 < 64'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_13 = io__in_bits_src1 >= 64'h40600000 & io__in_bits_src1 < 64'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_16 = io__in_bits_src1 >= 64'h50000000 & io__in_bits_src1 < 64'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_19 = io__in_bits_src1 >= 64'h40001000 & io__in_bits_src1 < 64'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_22 = io__in_bits_src1 >= 64'h40000000 & io__in_bits_src1 < 64'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_25 = io__in_bits_src1 >= 64'h40002000 & io__in_bits_src1 < 64'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_28 = io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _io_loadAccessFault_T_29 = {_io_loadAccessFault_T_28,_io_loadAccessFault_T_25,_io_loadAccessFault_T_22,
    _io_loadAccessFault_T_19,_io_loadAccessFault_T_16,_io_loadAccessFault_T_13,_io_loadAccessFault_T_10,
    _io_loadAccessFault_T_7}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _io_loadAccessFault_T_30 = |_io_loadAccessFault_T_29; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _io_loadAccessFault_T_31 = ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:71]
  wire  _io_storeAccessFault_T_33 = |(io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _T_30 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_31 = io__dmem_req_valid & _T_30; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  wire  _T_33 = _T_31 & _T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 534:39]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_346_clock;
  wire  line_346_reset;
  wire  line_346_valid;
  reg  line_346_valid_reg;
  wire  _GEN_27 = _T_31 | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_347_clock;
  wire  line_347_reset;
  wire  line_347_valid;
  reg  line_347_valid_reg;
  wire  _T_42 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  reg  r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_348_clock;
  wire  line_348_reset;
  wire  line_348_valid;
  reg  line_348_valid_reg;
  wire  _GEN_29 = _T_42 | r_1; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_349_clock;
  wire  line_349_reset;
  wire  line_349_valid;
  reg  line_349_valid_reg;
  GEN_w1_line #(.COVER_INDEX(333)) line_333 (
    .clock(line_333_clock),
    .reset(line_333_reset),
    .valid(line_333_valid)
  );
  GEN_w1_line #(.COVER_INDEX(334)) line_334 (
    .clock(line_334_clock),
    .reset(line_334_reset),
    .valid(line_334_valid)
  );
  GEN_w1_line #(.COVER_INDEX(335)) line_335 (
    .clock(line_335_clock),
    .reset(line_335_reset),
    .valid(line_335_valid)
  );
  GEN_w1_line #(.COVER_INDEX(336)) line_336 (
    .clock(line_336_clock),
    .reset(line_336_reset),
    .valid(line_336_valid)
  );
  GEN_w1_line #(.COVER_INDEX(337)) line_337 (
    .clock(line_337_clock),
    .reset(line_337_reset),
    .valid(line_337_valid)
  );
  GEN_w1_line #(.COVER_INDEX(338)) line_338 (
    .clock(line_338_clock),
    .reset(line_338_reset),
    .valid(line_338_valid)
  );
  GEN_w1_line #(.COVER_INDEX(339)) line_339 (
    .clock(line_339_clock),
    .reset(line_339_reset),
    .valid(line_339_valid)
  );
  GEN_w1_line #(.COVER_INDEX(340)) line_340 (
    .clock(line_340_clock),
    .reset(line_340_reset),
    .valid(line_340_valid)
  );
  GEN_w1_line #(.COVER_INDEX(341)) line_341 (
    .clock(line_341_clock),
    .reset(line_341_reset),
    .valid(line_341_valid)
  );
  GEN_w1_line #(.COVER_INDEX(342)) line_342 (
    .clock(line_342_clock),
    .reset(line_342_reset),
    .valid(line_342_valid)
  );
  GEN_w1_line #(.COVER_INDEX(343)) line_343 (
    .clock(line_343_clock),
    .reset(line_343_reset),
    .valid(line_343_valid)
  );
  GEN_w1_line #(.COVER_INDEX(344)) line_344 (
    .clock(line_344_clock),
    .reset(line_344_reset),
    .valid(line_344_valid)
  );
  GEN_w1_line #(.COVER_INDEX(345)) line_345 (
    .clock(line_345_clock),
    .reset(line_345_reset),
    .valid(line_345_valid)
  );
  GEN_w1_line #(.COVER_INDEX(346)) line_346 (
    .clock(line_346_clock),
    .reset(line_346_reset),
    .valid(line_346_valid)
  );
  GEN_w1_line #(.COVER_INDEX(347)) line_347 (
    .clock(line_347_clock),
    .reset(line_347_reset),
    .valid(line_347_valid)
  );
  GEN_w1_line #(.COVER_INDEX(348)) line_348 (
    .clock(line_348_clock),
    .reset(line_348_reset),
    .valid(line_348_valid)
  );
  GEN_w1_line #(.COVER_INDEX(349)) line_349 (
    .clock(line_349_clock),
    .reset(line_349_reset),
    .valid(line_349_valid)
  );
  assign line_333_clock = clock;
  assign line_333_reset = reset;
  assign line_333_valid = _io_vaddr_T ^ line_333_valid_reg;
  assign line_334_clock = clock;
  assign line_334_reset = reset;
  assign line_334_valid = _T ^ line_334_valid_reg;
  assign line_335_clock = clock;
  assign line_335_reset = reset;
  assign line_335_valid = _T_2 ^ line_335_valid_reg;
  assign line_336_clock = clock;
  assign line_336_reset = reset;
  assign line_336_valid = _T_5 ^ line_336_valid_reg;
  assign line_337_clock = clock;
  assign line_337_reset = reset;
  assign line_337_valid = _T ^ line_337_valid_reg;
  assign line_338_clock = clock;
  assign line_338_reset = reset;
  assign line_338_valid = _T_6 ^ line_338_valid_reg;
  assign line_339_clock = clock;
  assign line_339_reset = reset;
  assign line_339_valid = _T_9 ^ line_339_valid_reg;
  assign line_340_clock = clock;
  assign line_340_reset = reset;
  assign line_340_valid = _T_12 ^ line_340_valid_reg;
  assign line_341_clock = clock;
  assign line_341_reset = reset;
  assign line_341_valid = _T_6 ^ line_341_valid_reg;
  assign line_342_clock = clock;
  assign line_342_reset = reset;
  assign line_342_valid = _T_13 ^ line_342_valid_reg;
  assign line_343_clock = clock;
  assign line_343_reset = reset;
  assign line_343_valid = _T_14 ^ line_343_valid_reg;
  assign line_344_clock = clock;
  assign line_344_reset = reset;
  assign line_344_valid = _T_13 ^ line_344_valid_reg;
  assign line_345_clock = clock;
  assign line_345_reset = reset;
  assign line_345_valid = _T_15 ^ line_345_valid_reg;
  assign line_346_clock = clock;
  assign line_346_reset = reset;
  assign line_346_valid = _T_31 ^ line_346_valid_reg;
  assign line_347_clock = clock;
  assign line_347_reset = reset;
  assign line_347_valid = _T_14 ^ line_347_valid_reg;
  assign line_348_clock = clock;
  assign line_348_reset = reset;
  assign line_348_valid = _T_42 ^ line_348_valid_reg;
  assign line_349_clock = clock;
  assign line_349_reset = reset;
  assign line_349_valid = _T_14 ^ line_349_valid_reg;
  assign io__in_ready = _io_dmem_req_valid_T | dtlbHasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 487:37]
  assign io__out_valid = dtlbHasException & state != 2'h0 | hasException | _io_out_valid_T_7; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 480:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 520:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:49]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 466:68]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _reqWdata_T_18 | _reqWdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__dmem_resp_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 478:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 443:23]
  assign io__dtlbAF = DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 431:24]
  assign io__vaddr = _io_vaddr_T ? io__in_bits_src1 : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io__loadAccessFault = io__in_valid & _T_4 & ~(isStore | ISAMO2) & ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:68]
  assign io__storeAccessFault = _io_loadAccessFault_T_1 & (isStore & _io_loadAccessFault_T_31 | ISAMO2 & ~
    _io_storeAccessFault_T_33); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 532:45]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= io__in_bits_src1; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_333_valid_reg <= _io_vaddr_T;
    addrLatch <= io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
      state <= 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    end else if (2'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (_T_1 & ~vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:45]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:53]
      end else if (_T_1 & vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:45]
        state <= 2'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:53]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (DTLBFINISH & ~dtlbHasException & scIsSuccess_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:61]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:69]
      end else begin
        state <= _GEN_20;
      end
    end else if (2'h2 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      state <= _GEN_22;
    end else begin
      state <= _GEN_23;
    end
    line_334_valid_reg <= _T;
    line_335_valid_reg <= _T_2;
    line_336_valid_reg <= _T_5;
    line_337_valid_reg <= _T;
    line_338_valid_reg <= _T_6;
    line_339_valid_reg <= _T_9;
    line_340_valid_reg <= _T_12;
    line_341_valid_reg <= _T_6;
    line_342_valid_reg <= _T_13;
    line_343_valid_reg <= _T_14;
    line_344_valid_reg <= _T_13;
    line_345_valid_reg <= _T_15;
    rdataLatch <= io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_27;
    end
    line_346_valid_reg <= _T_31;
    line_347_valid_reg <= _T_14;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r_1 <= _GEN_29;
    end
    line_348_valid_reg <= _T_42;
    line_349_valid_reg <= _T_14;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  line_333_valid_reg = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  addrLatch = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  line_334_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_335_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_336_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_337_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_338_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_339_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_340_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_341_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_342_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_343_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_344_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_345_valid_reg = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  rdataLatch = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_346_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_347_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_348_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_349_valid_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_io_vaddr_T) begin
      cover(1'h1);
    end
    //
    if (_T) begin
      cover(1'h1);
    end
    //
    if (_T & _T_2) begin
      cover(1'h1);
    end
    //
    if (_T & _T_5) begin
      cover(1'h1);
    end
    //
    if (~_T) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_6) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_6 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_6 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_6) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_6 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_6 & _T_13 & _T_14) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_6 & ~_T_13) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_6 & ~_T_13 & _T_15) begin
      cover(1'h1);
    end
    //
    if (_T_31) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
    //
    if (_T_42) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
  end
endmodule
module AtomALU(
  input         clock,
  input         reset,
  input  [63:0] io_src1, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [63:0] io_src2, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [6:0]  io_func, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input         io_isWordOp, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  output [63:0] io_result // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
);
  wire  src1_signBit = io_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src1_T_1 = src1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src1_T_2 = {_src1_T_1,io_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src1 = io_isWordOp ? _src1_T_2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 183:17]
  wire  src2_signBit = io_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src2_T_1 = src2_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src2_T_2 = {_src2_T_1,io_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src2 = io_isWordOp ? _src2_T_2 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 184:17]
  wire  isAdderSub = ~io_func[6]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 186:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:39]
  wire [63:0] _adderRes_T_1 = src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:33]
  wire [64:0] _adderRes_T_2 = src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [63:0] xorRes = src1 ^ src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 188:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 189:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/LSU.scala 190:28]
  wire [63:0] _res_T_1 = src1 & src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 196:32]
  wire [63:0] _res_T_2 = src1 | src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 197:32]
  wire [63:0] _res_T_4 = slt ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 198:29]
  wire [63:0] _res_T_6 = slt ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 199:29]
  wire [63:0] _res_T_8 = sltu ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 200:29]
  wire [63:0] _res_T_10 = sltu ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 201:29]
  wire [64:0] _res_T_12 = 6'h22 == io_func[5:0] ? {{1'd0}, src2} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 6'h25 == io_func[5:0] ? {{1'd0}, _res_T_1} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 6'h26 == io_func[5:0] ? {{1'd0}, _res_T_2} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 6'h37 == io_func[5:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 6'h30 == io_func[5:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 6'h31 == io_func[5:0] ? {{1'd0}, _res_T_8} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  assign io_result = res[63:0]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 204:13]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src2, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [31:0] io__instr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        setLr_0,
  input         lr_0,
  output        scInflight_0,
  output        amoReq_0,
  input  [63:0] lr_addr,
  input  [55:0] dtlb_paddr,
  input         _T_12_0,
  input         scIsSuccess_0,
  output        setLrVal_0,
  input         vmEnable,
  input         DTLBFINISH,
  input         lsuMMIO_0,
  input         _T_13_1,
  output [63:0] setLrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__vaddr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_ISAMO2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBFINISH; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  atomALU_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  atomALU_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [6:0] atomALU_io_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  atomALU_io_isWordOp; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  isAtomic = io__in_bits_func[5]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 54:38]
  wire  _isAmo_T_1 = io__in_bits_func == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _isAmo_T_4 = io__in_bits_func == 7'h21; // @[src/main/scala/nutcore/backend/fu/LSU.scala 58:37]
  wire  isAmo = isAtomic & ~_isAmo_T_1 & ~_isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/LSU.scala 59:61]
  wire [63:0] _in_vaddr_T_1 = io__in_bits_src1 + io__in_bits_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:43]
  wire [63:0] in_vaddr = isAtomic ? io__in_bits_src1 : _in_vaddr_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
  wire [1:0] _in_func_T_1 = io__instr[12] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:34]
  wire [1:0] in_func = isAtomic ? _in_func_T_1 : io__in_bits_func[1:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:20]
  wire  _addrAligned_T_1 = ~in_vaddr[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 69:29]
  wire  _addrAligned_T_3 = in_vaddr[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 70:32]
  wire  _addrAligned_T_5 = in_vaddr[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 71:32]
  wire  _addrAligned_T_6 = 2'h0 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_7 = 2'h1 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_8 = 2'h2 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_9 = 2'h3 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  addrAligned = _addrAligned_T_6 | _addrAligned_T_7 & _addrAligned_T_1 | _addrAligned_T_8 & _addrAligned_T_3 |
    _addrAligned_T_9 & _addrAligned_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  hasAddrMisaligned = io__in_valid & ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 73:36]
  wire  _io_loadAddrMisaligned_T_4 = ~io__in_bits_func[3] & ~isAtomic; // @[src/main/scala/nutcore/backend/fu/LSU.scala 56:49]
  wire  _hasScAccessFault_T_1 = ~vmEnable; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:46]
  wire  _hasScAccessFault_T_6 = |(in_vaddr >= 64'h80000000 & in_vaddr < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  hasScAccessFault = io__in_valid & _isAmo_T_4 & ~vmEnable & ~_hasScAccessFault_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:58]
  wire  valid = io__in_valid & addrAligned & ~hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 86:39]
  wire  _io_vaddr_T_2 = hasAddrMisaligned | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 91:44]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_350_clock;
  wire  line_350_reset;
  wire  line_350_valid;
  reg  line_350_valid_reg;
  wire [63:0] _GEN_28 = _io_vaddr_T_2 ? in_vaddr : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  atomReq = valid & isAtomic; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 97:23]
  wire  amoReq = valid & isAmo; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:22]
  wire  lrReq = valid & _isAmo_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 99:21]
  wire  scReq = valid & _isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 100:21]
  wire [2:0] funct3 = io__instr[14:12]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 108:24]
  wire  scInvalid = scReq & (io__in_bits_src1 != lr_addr | ~lr_0) & _hasScAccessFault_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 126:53]
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
  reg [63:0] atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
  reg [63:0] atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
  wire  _T = 3'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_351_clock;
  wire  line_351_reset;
  wire  line_351_valid;
  reg  line_351_valid_reg;
  wire  line_352_clock;
  wire  line_352_reset;
  wire  line_352_valid;
  reg  line_352_valid_reg;
  wire  _lsExecUnit_io_in_valid_T = ~atomReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 184:48]
  wire  _io_in_ready_T_1 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_353_clock;
  wire  line_353_reset;
  wire  line_353_valid;
  reg  line_353_valid_reg;
  wire [2:0] _GEN_30 = amoReq ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 192:15 195:{19,26}]
  wire  line_354_clock;
  wire  line_354_reset;
  wire  line_354_valid;
  reg  line_354_valid_reg;
  wire [2:0] _GEN_31 = lrReq ? 3'h3 : _GEN_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 196:{18,25}]
  wire  line_355_clock;
  wire  line_355_reset;
  wire  line_355_valid;
  reg  line_355_valid_reg;
  wire [2:0] _state_T = scInvalid ? 3'h0 : 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:31]
  wire  line_356_clock;
  wire  line_356_reset;
  wire  line_356_valid;
  reg  line_356_valid_reg;
  wire  _T_1 = 3'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_357_clock;
  wire  line_357_reset;
  wire  line_357_valid;
  reg  line_357_valid_reg;
  wire  _T_10 = ~reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
  wire  line_358_clock;
  wire  line_358_reset;
  wire  line_358_valid;
  reg  line_358_valid_reg;
  wire  _T_11 = ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
  wire  line_359_clock;
  wire  line_359_reset;
  wire  line_359_valid;
  reg  line_359_valid_reg;
  wire  line_360_clock;
  wire  line_360_reset;
  wire  line_360_valid;
  reg  line_360_valid_reg;
  wire [2:0] _GEN_33 = io__out_valid ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22 211:{26,33}]
  wire  line_361_clock;
  wire  line_361_reset;
  wire  line_361_valid;
  reg  line_361_valid_reg;
  wire  _T_13 = 3'h5 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_362_clock;
  wire  line_362_reset;
  wire  line_362_valid;
  reg  line_362_valid_reg;
  wire [1:0] _lsExecUnit_io_in_bits_func_T = funct3[0] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 231:40]
  wire  line_363_clock;
  wire  line_363_reset;
  wire  line_363_valid;
  reg  line_363_valid_reg;
  wire [2:0] _GEN_34 = _io_in_ready_T_1 ? 3'h6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 235:37 236:15 132:22]
  wire  line_364_clock;
  wire  line_364_reset;
  wire  line_364_valid;
  reg  line_364_valid_reg;
  wire  _T_15 = 3'h6 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_365_clock;
  wire  line_365_reset;
  wire  line_365_valid;
  reg  line_365_valid_reg;
  wire  line_366_clock;
  wire  line_366_reset;
  wire  line_366_valid;
  reg  line_366_valid_reg;
  wire  _T_16 = 3'h7 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_367_clock;
  wire  line_367_reset;
  wire  line_367_valid;
  reg  line_367_valid_reg;
  wire [3:0] _lsExecUnit_io_in_bits_func_T_1 = funct3[0] ? 4'hb : 4'ha; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 262:40]
  wire  line_368_clock;
  wire  line_368_reset;
  wire  line_368_valid;
  reg  line_368_valid_reg;
  wire [2:0] _GEN_35 = _io_in_ready_T_1 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 266:37 267:15 132:22]
  wire  line_369_clock;
  wire  line_369_reset;
  wire  line_369_valid;
  reg  line_369_valid_reg;
  wire  _T_18 = 3'h3 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_370_clock;
  wire  line_370_reset;
  wire  line_370_valid;
  reg  line_370_valid_reg;
  wire  line_371_clock;
  wire  line_371_reset;
  wire  line_371_valid;
  reg  line_371_valid_reg;
  wire  line_372_clock;
  wire  line_372_reset;
  wire  line_372_valid;
  reg  line_372_valid_reg;
  wire  _T_20 = 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  line_373_clock;
  wire  line_373_reset;
  wire  line_373_valid;
  reg  line_373_valid_reg;
  wire  _io_in_ready_T_7 = ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 292:63]
  wire  _io_in_ready_T_8 = _io_in_ready_T_1 | ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 292:60]
  wire  line_374_clock;
  wire  line_374_reset;
  wire  line_374_valid;
  reg  line_374_valid_reg;
  wire [2:0] _GEN_37 = _io_in_ready_T_8 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 294:51 295:15 132:22]
  wire  _GEN_43 = 3'h4 == state & (_io_in_ready_T_1 | ~scIsSuccess_0); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 167:30 292:34]
  wire [2:0] _GEN_45 = 3'h4 == state ? _GEN_37 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 132:22]
  wire  _GEN_46 = 3'h3 == state | 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 272:34]
  wire [3:0] _GEN_49 = 3'h3 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _lsExecUnit_io_in_bits_func_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 276:34]
  wire  _GEN_51 = 3'h3 == state ? _io_in_ready_T_1 : _GEN_43; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 278:34]
  wire [2:0] _GEN_53 = 3'h3 == state ? _GEN_35 : _GEN_45; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_54 = 3'h7 == state | _GEN_46; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 258:34]
  wire [3:0] _GEN_57 = 3'h7 == state ? _lsExecUnit_io_in_bits_func_T_1 : _GEN_49; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 262:34]
  wire [63:0] _GEN_58 = 3'h7 == state ? atomMemReg : io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 263:34]
  wire  _GEN_59 = 3'h7 == state ? _io_in_ready_T_1 : _GEN_51; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 264:34]
  wire [2:0] _GEN_61 = 3'h7 == state ? _GEN_35 : _GEN_53; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_62 = 3'h6 == state ? 1'h0 : _GEN_54; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 244:34]
  wire  _GEN_63 = 3'h6 == state ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 245:34]
  wire  _GEN_67 = 3'h6 == state ? 1'h0 : _GEN_59; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 250:34]
  wire [2:0] _GEN_69 = 3'h6 == state ? 3'h7 : _GEN_61; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 252:13]
  wire  _GEN_71 = 3'h5 == state | _GEN_62; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 227:34]
  wire  _GEN_72 = 3'h5 == state | _GEN_63; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 228:34]
  wire [3:0] _GEN_74 = 3'h5 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _GEN_57; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 231:34]
  wire  _GEN_76 = 3'h5 == state ? 1'h0 : _GEN_67; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 233:34]
  wire [2:0] _GEN_78 = 3'h5 == state ? _GEN_34 : _GEN_69; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_81 = 3'h1 == state | _GEN_71; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 202:34]
  wire  _GEN_82 = 3'h1 == state | _GEN_72; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 203:34]
  wire [6:0] _GEN_84 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_74}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 206:34]
  wire [63:0] _GEN_85 = 3'h1 == state ? io__wdata : _GEN_58; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 207:34]
  wire  _GEN_87 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_76; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 209:34]
  wire  _GEN_97 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_87; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 191:36]
  wire  _hasException_T_1 = lsExecUnit_io__dtlbAF | lsExecUnit_io__dtlbPF | io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 300:67]
  wire  _hasException_T_3 = _hasException_T_1 | io__storeAddrMisaligned | io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 301:53]
  wire  hasException = _hasException_T_3 | io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 302:24]
  wire  line_375_clock;
  wire  line_375_reset;
  wire  line_375_valid;
  reg  line_375_valid_reg;
  wire [31:0] lr_paddr = dtlb_paddr[31:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 316:26]
  wire  _io_out_bits_T_1 = scInvalid | _io_in_ready_T_7; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:39]
  wire [63:0] _io_out_bits_T_3 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:59]
  reg  mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
  wire  _T_25 = ~mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:9]
  wire  line_376_clock;
  wire  line_376_reset;
  wire  line_376_valid;
  reg  line_376_valid_reg;
  wire  line_377_clock;
  wire  line_377_reset;
  wire  line_377_valid;
  reg  line_377_valid_reg;
  wire  setLr = io__out_valid & (lrReq | scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 318:24]
  wire  setLrVal = lrReq & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 319:21]
  wire [63:0] setLrAddr = vmEnable ? {{32'd0}, lr_paddr} : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 320:19]
  wire  scInflight = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 143:23]
  LSExecUnit lsExecUnit ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_ready(lsExecUnit_io__in_ready),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__dtlbAF(lsExecUnit_io__dtlbAF),
    .io__vaddr(lsExecUnit_io__vaddr),
    .io__loadAccessFault(lsExecUnit_io__loadAccessFault),
    .io__storeAccessFault(lsExecUnit_io__storeAccessFault),
    .DTLBPF(lsExecUnit_DTLBPF),
    .scIsSuccess_0(lsExecUnit_scIsSuccess_0),
    .vmEnable_0(lsExecUnit_vmEnable_0),
    .ISAMO2(lsExecUnit_ISAMO2),
    .DTLBFINISH(lsExecUnit_DTLBFINISH),
    .DTLBAF(lsExecUnit_DTLBAF)
  );
  AtomALU atomALU ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
    .clock(atomALU_clock),
    .reset(atomALU_reset),
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  GEN_w1_line #(.COVER_INDEX(350)) line_350 (
    .clock(line_350_clock),
    .reset(line_350_reset),
    .valid(line_350_valid)
  );
  GEN_w1_line #(.COVER_INDEX(351)) line_351 (
    .clock(line_351_clock),
    .reset(line_351_reset),
    .valid(line_351_valid)
  );
  GEN_w1_line #(.COVER_INDEX(352)) line_352 (
    .clock(line_352_clock),
    .reset(line_352_reset),
    .valid(line_352_valid)
  );
  GEN_w1_line #(.COVER_INDEX(353)) line_353 (
    .clock(line_353_clock),
    .reset(line_353_reset),
    .valid(line_353_valid)
  );
  GEN_w1_line #(.COVER_INDEX(354)) line_354 (
    .clock(line_354_clock),
    .reset(line_354_reset),
    .valid(line_354_valid)
  );
  GEN_w1_line #(.COVER_INDEX(355)) line_355 (
    .clock(line_355_clock),
    .reset(line_355_reset),
    .valid(line_355_valid)
  );
  GEN_w1_line #(.COVER_INDEX(356)) line_356 (
    .clock(line_356_clock),
    .reset(line_356_reset),
    .valid(line_356_valid)
  );
  GEN_w1_line #(.COVER_INDEX(357)) line_357 (
    .clock(line_357_clock),
    .reset(line_357_reset),
    .valid(line_357_valid)
  );
  GEN_w1_line #(.COVER_INDEX(358)) line_358 (
    .clock(line_358_clock),
    .reset(line_358_reset),
    .valid(line_358_valid)
  );
  GEN_w1_line #(.COVER_INDEX(359)) line_359 (
    .clock(line_359_clock),
    .reset(line_359_reset),
    .valid(line_359_valid)
  );
  GEN_w1_line #(.COVER_INDEX(360)) line_360 (
    .clock(line_360_clock),
    .reset(line_360_reset),
    .valid(line_360_valid)
  );
  GEN_w1_line #(.COVER_INDEX(361)) line_361 (
    .clock(line_361_clock),
    .reset(line_361_reset),
    .valid(line_361_valid)
  );
  GEN_w1_line #(.COVER_INDEX(362)) line_362 (
    .clock(line_362_clock),
    .reset(line_362_reset),
    .valid(line_362_valid)
  );
  GEN_w1_line #(.COVER_INDEX(363)) line_363 (
    .clock(line_363_clock),
    .reset(line_363_reset),
    .valid(line_363_valid)
  );
  GEN_w1_line #(.COVER_INDEX(364)) line_364 (
    .clock(line_364_clock),
    .reset(line_364_reset),
    .valid(line_364_valid)
  );
  GEN_w1_line #(.COVER_INDEX(365)) line_365 (
    .clock(line_365_clock),
    .reset(line_365_reset),
    .valid(line_365_valid)
  );
  GEN_w1_line #(.COVER_INDEX(366)) line_366 (
    .clock(line_366_clock),
    .reset(line_366_reset),
    .valid(line_366_valid)
  );
  GEN_w1_line #(.COVER_INDEX(367)) line_367 (
    .clock(line_367_clock),
    .reset(line_367_reset),
    .valid(line_367_valid)
  );
  GEN_w1_line #(.COVER_INDEX(368)) line_368 (
    .clock(line_368_clock),
    .reset(line_368_reset),
    .valid(line_368_valid)
  );
  GEN_w1_line #(.COVER_INDEX(369)) line_369 (
    .clock(line_369_clock),
    .reset(line_369_reset),
    .valid(line_369_valid)
  );
  GEN_w1_line #(.COVER_INDEX(370)) line_370 (
    .clock(line_370_clock),
    .reset(line_370_reset),
    .valid(line_370_valid)
  );
  GEN_w1_line #(.COVER_INDEX(371)) line_371 (
    .clock(line_371_clock),
    .reset(line_371_reset),
    .valid(line_371_valid)
  );
  GEN_w1_line #(.COVER_INDEX(372)) line_372 (
    .clock(line_372_clock),
    .reset(line_372_reset),
    .valid(line_372_valid)
  );
  GEN_w1_line #(.COVER_INDEX(373)) line_373 (
    .clock(line_373_clock),
    .reset(line_373_reset),
    .valid(line_373_valid)
  );
  GEN_w1_line #(.COVER_INDEX(374)) line_374 (
    .clock(line_374_clock),
    .reset(line_374_reset),
    .valid(line_374_valid)
  );
  GEN_w1_line #(.COVER_INDEX(375)) line_375 (
    .clock(line_375_clock),
    .reset(line_375_reset),
    .valid(line_375_valid)
  );
  GEN_w1_line #(.COVER_INDEX(376)) line_376 (
    .clock(line_376_clock),
    .reset(line_376_reset),
    .valid(line_376_valid)
  );
  GEN_w1_line #(.COVER_INDEX(377)) line_377 (
    .clock(line_377_clock),
    .reset(line_377_reset),
    .valid(line_377_valid)
  );
  assign line_350_clock = clock;
  assign line_350_reset = reset;
  assign line_350_valid = _io_vaddr_T_2 ^ line_350_valid_reg;
  assign line_351_clock = clock;
  assign line_351_reset = reset;
  assign line_351_valid = _T ^ line_351_valid_reg;
  assign line_352_clock = clock;
  assign line_352_reset = reset;
  assign line_352_valid = valid ^ line_352_valid_reg;
  assign line_353_clock = clock;
  assign line_353_reset = reset;
  assign line_353_valid = amoReq ^ line_353_valid_reg;
  assign line_354_clock = clock;
  assign line_354_reset = reset;
  assign line_354_valid = lrReq ^ line_354_valid_reg;
  assign line_355_clock = clock;
  assign line_355_reset = reset;
  assign line_355_valid = scReq ^ line_355_valid_reg;
  assign line_356_clock = clock;
  assign line_356_reset = reset;
  assign line_356_valid = _T ^ line_356_valid_reg;
  assign line_357_clock = clock;
  assign line_357_reset = reset;
  assign line_357_valid = _T_1 ^ line_357_valid_reg;
  assign line_358_clock = clock;
  assign line_358_reset = reset;
  assign line_358_valid = _T_10 ^ line_358_valid_reg;
  assign line_359_clock = clock;
  assign line_359_reset = reset;
  assign line_359_valid = _T_11 ^ line_359_valid_reg;
  assign line_360_clock = clock;
  assign line_360_reset = reset;
  assign line_360_valid = io__out_valid ^ line_360_valid_reg;
  assign line_361_clock = clock;
  assign line_361_reset = reset;
  assign line_361_valid = _T_1 ^ line_361_valid_reg;
  assign line_362_clock = clock;
  assign line_362_reset = reset;
  assign line_362_valid = _T_13 ^ line_362_valid_reg;
  assign line_363_clock = clock;
  assign line_363_reset = reset;
  assign line_363_valid = _io_in_ready_T_1 ^ line_363_valid_reg;
  assign line_364_clock = clock;
  assign line_364_reset = reset;
  assign line_364_valid = _T_13 ^ line_364_valid_reg;
  assign line_365_clock = clock;
  assign line_365_reset = reset;
  assign line_365_valid = _T_15 ^ line_365_valid_reg;
  assign line_366_clock = clock;
  assign line_366_reset = reset;
  assign line_366_valid = _T_15 ^ line_366_valid_reg;
  assign line_367_clock = clock;
  assign line_367_reset = reset;
  assign line_367_valid = _T_16 ^ line_367_valid_reg;
  assign line_368_clock = clock;
  assign line_368_reset = reset;
  assign line_368_valid = _io_in_ready_T_1 ^ line_368_valid_reg;
  assign line_369_clock = clock;
  assign line_369_reset = reset;
  assign line_369_valid = _T_16 ^ line_369_valid_reg;
  assign line_370_clock = clock;
  assign line_370_reset = reset;
  assign line_370_valid = _T_18 ^ line_370_valid_reg;
  assign line_371_clock = clock;
  assign line_371_reset = reset;
  assign line_371_valid = _io_in_ready_T_1 ^ line_371_valid_reg;
  assign line_372_clock = clock;
  assign line_372_reset = reset;
  assign line_372_valid = _T_18 ^ line_372_valid_reg;
  assign line_373_clock = clock;
  assign line_373_reset = reset;
  assign line_373_valid = _T_20 ^ line_373_valid_reg;
  assign line_374_clock = clock;
  assign line_374_reset = reset;
  assign line_374_valid = _io_in_ready_T_8 ^ line_374_valid_reg;
  assign line_375_clock = clock;
  assign line_375_reset = reset;
  assign line_375_valid = hasException ^ line_375_valid_reg;
  assign line_376_clock = clock;
  assign line_376_reset = reset;
  assign line_376_valid = _T_25 ^ line_376_valid_reg;
  assign line_377_clock = clock;
  assign line_377_reset = reset;
  assign line_377_valid = io__out_valid ^ line_377_valid_reg;
  assign io__out_valid = hasException | _GEN_97; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23 305:18]
  assign io__out_bits = scReq ? {{63'd0}, _io_out_bits_T_1} : _io_out_bits_T_3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:21]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__isMMIO = mmioReg & io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 332:24]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 94:13]
  assign io__dtlbAF = lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:13]
  assign io__vaddr = io__loadAddrMisaligned | io__storeAddrMisaligned | hasScAccessFault ? _GEN_28 :
    lsExecUnit_io__vaddr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 90:18]
  assign io__loadAddrMisaligned = hasAddrMisaligned & (_io_loadAddrMisaligned_T_4 | _isAmo_T_1); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 74:46]
  assign io__storeAddrMisaligned = hasAddrMisaligned & (io__in_bits_func[3] | isAmo | _isAmo_T_4); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 75:47]
  assign io__loadAccessFault = lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 334:22]
  assign io__storeAccessFault = lsExecUnit_io__storeAccessFault | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:57]
  assign setLr_0 = setLr;
  assign scInflight_0 = scInflight;
  assign amoReq_0 = amoReq;
  assign setLrVal_0 = setLrVal;
  assign setLrAddr_0 = setLrAddr;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? valid & ~atomReq : _GEN_81; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 184:36]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _in_vaddr_T_1 : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 186:36]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_84; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 188:36]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_82; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 185:36]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_85; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 189:36]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_DTLBPF = _T_12_0;
  assign lsExecUnit_scIsSuccess_0 = scIsSuccess_0;
  assign lsExecUnit_vmEnable_0 = vmEnable;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign lsExecUnit_DTLBAF = _T_13_1;
  assign atomALU_clock = clock;
  assign atomALU_reset = reset;
  assign atomALU_io_src1 = atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 136:19]
  assign atomALU_io_src2 = io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 137:19]
  assign atomALU_io_func = io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 138:19]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 110:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T_2) begin // @[src/main/scala/utils/Hold.scala 23:65]
      if (isAtomic) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
        io_vaddr_r <= io__in_bits_src1;
      end else begin
        io_vaddr_r <= _in_vaddr_T_1;
      end
    end
    line_350_valid_reg <= _io_vaddr_T_2;
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 304:11]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (scReq) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:18]
        state <= _state_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:25]
      end else begin
        state <= _GEN_31;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      state <= _GEN_33;
    end else begin
      state <= _GEN_78;
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 239:18]
        end else if (3'h6 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 253:18]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomRegReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 240:18]
        end
      end
    end
    line_351_valid_reg <= _T;
    line_352_valid_reg <= valid;
    line_353_valid_reg <= amoReq;
    line_354_valid_reg <= lrReq;
    line_355_valid_reg <= scReq;
    line_356_valid_reg <= _T;
    line_357_valid_reg <= _T_1;
    line_358_valid_reg <= _T_10;
    line_359_valid_reg <= _T_11;
    line_360_valid_reg <= io__out_valid;
    line_361_valid_reg <= _T_1;
    line_362_valid_reg <= _T_13;
    line_363_valid_reg <= _io_in_ready_T_1;
    line_364_valid_reg <= _T_13;
    line_365_valid_reg <= _T_15;
    line_366_valid_reg <= _T_15;
    line_367_valid_reg <= _T_16;
    line_368_valid_reg <= _io_in_ready_T_1;
    line_369_valid_reg <= _T_16;
    line_370_valid_reg <= _T_18;
    line_371_valid_reg <= _io_in_ready_T_1;
    line_372_valid_reg <= _T_18;
    line_373_valid_reg <= _T_20;
    line_374_valid_reg <= _io_in_ready_T_8;
    line_375_valid_reg <= hasException;
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
    end else if (io__out_valid) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:23]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:33]
    end else if (~mmioReg) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:19]
      mmioReg <= lsuMMIO_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:29]
    end
    line_376_valid_reg <= _T_25;
    line_377_valid_reg <= io__out_valid;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & _T_1 & _T_10 & ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:210 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  line_350_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  atomMemReg = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  atomRegReg = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  line_351_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_352_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_353_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_354_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_355_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_356_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_357_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_358_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_359_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_360_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_361_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_362_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_363_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_364_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_365_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_366_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_367_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_368_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_369_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_370_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_371_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_372_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_373_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_374_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_375_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mmioReg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_376_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_377_valid_reg = _RAND_32[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_io_vaddr_T_2) begin
      cover(1'h1);
    end
    //
    if (_T) begin
      cover(1'h1);
    end
    //
    if (_T & valid) begin
      cover(1'h1);
    end
    //
    if (_T & amoReq) begin
      cover(1'h1);
    end
    //
    if (_T & lrReq) begin
      cover(1'h1);
    end
    //
    if (_T & scReq) begin
      cover(1'h1);
    end
    //
    if (~_T) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_1) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_1 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_1 & _T_10 & _T_11) begin
      cover(1'h1);
    end
    //
    if (~_T & _T_1 & ~reset) begin
      assert(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
    end
    //
    if (~_T & _T_1 & io__out_valid) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & _T_13 & _io_in_ready_T_1) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & _T_15) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & _T_16) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & _T_16 & _io_in_ready_T_1) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16 & _T_18) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16 & _T_18 & _io_in_ready_T_1) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16 & ~_T_18) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16 & ~_T_18 & _T_20) begin
      cover(1'h1);
    end
    //
    if (~_T & ~_T_1 & ~_T_13 & ~_T_15 & ~_T_16 & ~_T_18 & _T_20 & _io_in_ready_T_8) begin
      cover(1'h1);
    end
    //
    if (hasException) begin
      cover(1'h1);
    end
    //
    if (_T_25) begin
      cover(1'h1);
    end
    //
    if (io__out_valid) begin
      cover(1'h1);
    end
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output [129:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [64:0] mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [129:0] io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg [129:0] io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg [129:0] io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg  io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg  io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg  io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  _T_1 = io_in_valid & ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 63:21]
  wire  line_378_clock;
  wire  line_378_reset;
  wire  line_378_valid;
  reg  line_378_valid_reg;
  wire  _GEN_2 = io_in_valid & ~busy | busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21 63:{31,38}]
  wire  line_379_clock;
  wire  line_379_reset;
  wire  line_379_valid;
  reg  line_379_valid_reg;
  GEN_w1_line #(.COVER_INDEX(378)) line_378 (
    .clock(line_378_clock),
    .reset(line_378_reset),
    .valid(line_378_valid)
  );
  GEN_w1_line #(.COVER_INDEX(379)) line_379 (
    .clock(line_379_clock),
    .reset(line_379_reset),
    .valid(line_379_valid)
  );
  assign line_378_clock = clock;
  assign line_378_reset = reset;
  assign line_378_valid = _T_1 ^ line_378_valid_reg;
  assign line_379_clock = clock;
  assign line_379_reset = reset;
  assign line_379_valid = io_out_valid ^ line_379_valid_reg;
  assign io_in_ready = ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 65:49]
  assign io_out_valid = io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 60:16]
  assign io_out_bits = io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 59:37]
  always @(posedge clock) begin
    mulRes_REG <= io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    mulRes_REG_1 <= io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    io_out_bits_REG <= $signed(mulRes_REG) * $signed(mulRes_REG_1); // @[src/main/scala/nutcore/backend/fu/MDU.scala 58:49]
    io_out_bits_REG_1 <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_bits_REG_2 <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    io_out_valid_REG <= io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    io_out_valid_REG_1 <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    io_out_valid_REG_2 <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_valid_REG_3 <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end else if (io_out_valid) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:23]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:30]
    end else begin
      busy <= _GEN_2;
    end
    line_378_valid_reg <= _T_1;
    line_379_valid_reg <= io_out_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  mulRes_REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  mulRes_REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  io_out_bits_REG = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  io_out_bits_REG_1 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  io_out_bits_REG_2 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_378_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_379_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (io_out_valid) begin
      cover(1'h1);
    end
  end
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_sign, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output [127:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  _newReq_T_1 = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  newReq = state == 3'h0 & _newReq_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 81:18]
  reg [128:0] shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_1 = 64'h0 - io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_1 : io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_3 = 64'h0 - io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  reg  aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  wire  line_380_clock;
  wire  line_380_reset;
  wire  line_380_valid;
  reg  line_380_valid_reg;
  reg  qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  wire  line_381_clock;
  wire  line_381_reset;
  wire  line_381_valid;
  reg  line_381_valid_reg;
  reg [63:0] bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire  line_382_clock;
  wire  line_382_reset;
  wire  line_382_valid;
  reg  line_382_valid_reg;
  wire [64:0] _aValx2Reg_T = {aVal,1'h0}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:32]
  reg [64:0] aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  wire  line_383_clock;
  wire  line_383_reset;
  wire  line_383_valid;
  reg  line_383_valid_reg;
  reg [5:0] cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_384_clock;
  wire  line_384_reset;
  wire  line_384_valid;
  reg  line_384_valid_reg;
  wire  line_385_clock;
  wire  line_385_reset;
  wire  line_385_valid;
  reg  line_385_valid_reg;
  wire  _T_4 = state == 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:22]
  wire  line_386_clock;
  wire  line_386_reset;
  wire  line_386_valid;
  reg  line_386_valid_reg;
  wire [31:0] canSkipShift_hi = bReg[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo = bReg[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi = |canSkipShift_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_1 = canSkipShift_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_1 = canSkipShift_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_1 = |canSkipShift_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_2 = canSkipShift_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_2 = canSkipShift_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_2 = |canSkipShift_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_3 = canSkipShift_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_3 = canSkipShift_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_3 = |canSkipShift_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_3 = canSkipShift_hi_3[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_4 = canSkipShift_hi_3[3] ? 2'h3 : _canSkipShift_T_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_8 = canSkipShift_lo_3[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_9 = canSkipShift_lo_3[3] ? 2'h3 : _canSkipShift_T_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_10 = canSkipShift_useHi_3 ? _canSkipShift_T_4 : _canSkipShift_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_11 = {canSkipShift_useHi_3,_canSkipShift_T_10}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_4 = canSkipShift_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_4 = canSkipShift_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_4 = |canSkipShift_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_15 = canSkipShift_hi_4[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_16 = canSkipShift_hi_4[3] ? 2'h3 : _canSkipShift_T_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_20 = canSkipShift_lo_4[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_21 = canSkipShift_lo_4[3] ? 2'h3 : _canSkipShift_T_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_22 = canSkipShift_useHi_4 ? _canSkipShift_T_16 : _canSkipShift_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_23 = {canSkipShift_useHi_4,_canSkipShift_T_22}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_24 = canSkipShift_useHi_2 ? _canSkipShift_T_11 : _canSkipShift_T_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_25 = {canSkipShift_useHi_2,_canSkipShift_T_24}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_5 = canSkipShift_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_5 = canSkipShift_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_5 = |canSkipShift_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_6 = canSkipShift_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_6 = canSkipShift_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_6 = |canSkipShift_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_29 = canSkipShift_hi_6[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_30 = canSkipShift_hi_6[3] ? 2'h3 : _canSkipShift_T_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_34 = canSkipShift_lo_6[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_35 = canSkipShift_lo_6[3] ? 2'h3 : _canSkipShift_T_34; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_36 = canSkipShift_useHi_6 ? _canSkipShift_T_30 : _canSkipShift_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_37 = {canSkipShift_useHi_6,_canSkipShift_T_36}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_7 = canSkipShift_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_7 = canSkipShift_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_7 = |canSkipShift_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_41 = canSkipShift_hi_7[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_42 = canSkipShift_hi_7[3] ? 2'h3 : _canSkipShift_T_41; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_46 = canSkipShift_lo_7[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_47 = canSkipShift_lo_7[3] ? 2'h3 : _canSkipShift_T_46; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_48 = canSkipShift_useHi_7 ? _canSkipShift_T_42 : _canSkipShift_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_49 = {canSkipShift_useHi_7,_canSkipShift_T_48}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_50 = canSkipShift_useHi_5 ? _canSkipShift_T_37 : _canSkipShift_T_49; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_51 = {canSkipShift_useHi_5,_canSkipShift_T_50}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_52 = canSkipShift_useHi_1 ? _canSkipShift_T_25 : _canSkipShift_T_51; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_53 = {canSkipShift_useHi_1,_canSkipShift_T_52}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_8 = canSkipShift_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_8 = canSkipShift_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_8 = |canSkipShift_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_9 = canSkipShift_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_9 = canSkipShift_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_9 = |canSkipShift_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_10 = canSkipShift_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_10 = canSkipShift_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_10 = |canSkipShift_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_57 = canSkipShift_hi_10[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_58 = canSkipShift_hi_10[3] ? 2'h3 : _canSkipShift_T_57; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_62 = canSkipShift_lo_10[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_63 = canSkipShift_lo_10[3] ? 2'h3 : _canSkipShift_T_62; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_64 = canSkipShift_useHi_10 ? _canSkipShift_T_58 : _canSkipShift_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_65 = {canSkipShift_useHi_10,_canSkipShift_T_64}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_11 = canSkipShift_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_11 = canSkipShift_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_11 = |canSkipShift_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_69 = canSkipShift_hi_11[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_70 = canSkipShift_hi_11[3] ? 2'h3 : _canSkipShift_T_69; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_74 = canSkipShift_lo_11[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_75 = canSkipShift_lo_11[3] ? 2'h3 : _canSkipShift_T_74; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_76 = canSkipShift_useHi_11 ? _canSkipShift_T_70 : _canSkipShift_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_77 = {canSkipShift_useHi_11,_canSkipShift_T_76}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_78 = canSkipShift_useHi_9 ? _canSkipShift_T_65 : _canSkipShift_T_77; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_79 = {canSkipShift_useHi_9,_canSkipShift_T_78}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_12 = canSkipShift_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_12 = canSkipShift_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_12 = |canSkipShift_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_13 = canSkipShift_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_13 = canSkipShift_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_13 = |canSkipShift_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_83 = canSkipShift_hi_13[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_84 = canSkipShift_hi_13[3] ? 2'h3 : _canSkipShift_T_83; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_88 = canSkipShift_lo_13[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_89 = canSkipShift_lo_13[3] ? 2'h3 : _canSkipShift_T_88; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_90 = canSkipShift_useHi_13 ? _canSkipShift_T_84 : _canSkipShift_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_91 = {canSkipShift_useHi_13,_canSkipShift_T_90}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_14 = canSkipShift_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_14 = canSkipShift_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_14 = |canSkipShift_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_95 = canSkipShift_hi_14[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_96 = canSkipShift_hi_14[3] ? 2'h3 : _canSkipShift_T_95; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_100 = canSkipShift_lo_14[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_101 = canSkipShift_lo_14[3] ? 2'h3 : _canSkipShift_T_100; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_102 = canSkipShift_useHi_14 ? _canSkipShift_T_96 : _canSkipShift_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_103 = {canSkipShift_useHi_14,_canSkipShift_T_102}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_104 = canSkipShift_useHi_12 ? _canSkipShift_T_91 : _canSkipShift_T_103; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_105 = {canSkipShift_useHi_12,_canSkipShift_T_104}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_106 = canSkipShift_useHi_8 ? _canSkipShift_T_79 : _canSkipShift_T_105; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_107 = {canSkipShift_useHi_8,_canSkipShift_T_106}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_108 = canSkipShift_useHi ? _canSkipShift_T_53 : _canSkipShift_T_107; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_109 = {canSkipShift_useHi,_canSkipShift_T_108}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] _GEN_32 = {{1'd0}, _canSkipShift_T_109}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire [6:0] _canSkipShift_T_110 = 7'h40 | _GEN_32; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire  canSkipShift_hi_15 = aValx2Reg[64]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [63:0] canSkipShift_lo_15 = aValx2Reg[63:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_15 = |canSkipShift_hi_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [31:0] canSkipShift_hi_16 = canSkipShift_lo_15[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo_16 = canSkipShift_lo_15[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_16 = |canSkipShift_hi_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_17 = canSkipShift_hi_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_17 = canSkipShift_hi_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_17 = |canSkipShift_hi_17; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_18 = canSkipShift_hi_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_18 = canSkipShift_hi_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_18 = |canSkipShift_hi_18; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_19 = canSkipShift_hi_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_19 = canSkipShift_hi_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_19 = |canSkipShift_hi_19; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_114 = canSkipShift_hi_19[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_115 = canSkipShift_hi_19[3] ? 2'h3 : _canSkipShift_T_114; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_119 = canSkipShift_lo_19[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_120 = canSkipShift_lo_19[3] ? 2'h3 : _canSkipShift_T_119; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_121 = canSkipShift_useHi_19 ? _canSkipShift_T_115 : _canSkipShift_T_120; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_122 = {canSkipShift_useHi_19,_canSkipShift_T_121}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_20 = canSkipShift_lo_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_20 = canSkipShift_lo_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_20 = |canSkipShift_hi_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_126 = canSkipShift_hi_20[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_127 = canSkipShift_hi_20[3] ? 2'h3 : _canSkipShift_T_126; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_131 = canSkipShift_lo_20[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_132 = canSkipShift_lo_20[3] ? 2'h3 : _canSkipShift_T_131; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_133 = canSkipShift_useHi_20 ? _canSkipShift_T_127 : _canSkipShift_T_132; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_134 = {canSkipShift_useHi_20,_canSkipShift_T_133}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_135 = canSkipShift_useHi_18 ? _canSkipShift_T_122 : _canSkipShift_T_134; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_136 = {canSkipShift_useHi_18,_canSkipShift_T_135}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_21 = canSkipShift_lo_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_21 = canSkipShift_lo_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_21 = |canSkipShift_hi_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_22 = canSkipShift_hi_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_22 = canSkipShift_hi_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_22 = |canSkipShift_hi_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_140 = canSkipShift_hi_22[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_141 = canSkipShift_hi_22[3] ? 2'h3 : _canSkipShift_T_140; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_145 = canSkipShift_lo_22[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_146 = canSkipShift_lo_22[3] ? 2'h3 : _canSkipShift_T_145; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_147 = canSkipShift_useHi_22 ? _canSkipShift_T_141 : _canSkipShift_T_146; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_148 = {canSkipShift_useHi_22,_canSkipShift_T_147}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_23 = canSkipShift_lo_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_23 = canSkipShift_lo_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_23 = |canSkipShift_hi_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_152 = canSkipShift_hi_23[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_153 = canSkipShift_hi_23[3] ? 2'h3 : _canSkipShift_T_152; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_157 = canSkipShift_lo_23[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_158 = canSkipShift_lo_23[3] ? 2'h3 : _canSkipShift_T_157; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_159 = canSkipShift_useHi_23 ? _canSkipShift_T_153 : _canSkipShift_T_158; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_160 = {canSkipShift_useHi_23,_canSkipShift_T_159}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_161 = canSkipShift_useHi_21 ? _canSkipShift_T_148 : _canSkipShift_T_160; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_162 = {canSkipShift_useHi_21,_canSkipShift_T_161}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_163 = canSkipShift_useHi_17 ? _canSkipShift_T_136 : _canSkipShift_T_162; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_164 = {canSkipShift_useHi_17,_canSkipShift_T_163}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_24 = canSkipShift_lo_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_24 = canSkipShift_lo_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_24 = |canSkipShift_hi_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_25 = canSkipShift_hi_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_25 = canSkipShift_hi_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_25 = |canSkipShift_hi_25; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_26 = canSkipShift_hi_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_26 = canSkipShift_hi_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_26 = |canSkipShift_hi_26; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_168 = canSkipShift_hi_26[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_169 = canSkipShift_hi_26[3] ? 2'h3 : _canSkipShift_T_168; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_173 = canSkipShift_lo_26[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_174 = canSkipShift_lo_26[3] ? 2'h3 : _canSkipShift_T_173; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_175 = canSkipShift_useHi_26 ? _canSkipShift_T_169 : _canSkipShift_T_174; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_176 = {canSkipShift_useHi_26,_canSkipShift_T_175}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_27 = canSkipShift_lo_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_27 = canSkipShift_lo_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_27 = |canSkipShift_hi_27; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_180 = canSkipShift_hi_27[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_181 = canSkipShift_hi_27[3] ? 2'h3 : _canSkipShift_T_180; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_185 = canSkipShift_lo_27[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_186 = canSkipShift_lo_27[3] ? 2'h3 : _canSkipShift_T_185; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_187 = canSkipShift_useHi_27 ? _canSkipShift_T_181 : _canSkipShift_T_186; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_188 = {canSkipShift_useHi_27,_canSkipShift_T_187}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_189 = canSkipShift_useHi_25 ? _canSkipShift_T_176 : _canSkipShift_T_188; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_190 = {canSkipShift_useHi_25,_canSkipShift_T_189}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_28 = canSkipShift_lo_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_28 = canSkipShift_lo_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_28 = |canSkipShift_hi_28; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_29 = canSkipShift_hi_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_29 = canSkipShift_hi_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_29 = |canSkipShift_hi_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_194 = canSkipShift_hi_29[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_195 = canSkipShift_hi_29[3] ? 2'h3 : _canSkipShift_T_194; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_199 = canSkipShift_lo_29[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_200 = canSkipShift_lo_29[3] ? 2'h3 : _canSkipShift_T_199; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_201 = canSkipShift_useHi_29 ? _canSkipShift_T_195 : _canSkipShift_T_200; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_202 = {canSkipShift_useHi_29,_canSkipShift_T_201}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_30 = canSkipShift_lo_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_30 = canSkipShift_lo_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_30 = |canSkipShift_hi_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_206 = canSkipShift_hi_30[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_207 = canSkipShift_hi_30[3] ? 2'h3 : _canSkipShift_T_206; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_211 = canSkipShift_lo_30[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_212 = canSkipShift_lo_30[3] ? 2'h3 : _canSkipShift_T_211; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_213 = canSkipShift_useHi_30 ? _canSkipShift_T_207 : _canSkipShift_T_212; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_214 = {canSkipShift_useHi_30,_canSkipShift_T_213}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_215 = canSkipShift_useHi_28 ? _canSkipShift_T_202 : _canSkipShift_T_214; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_216 = {canSkipShift_useHi_28,_canSkipShift_T_215}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_217 = canSkipShift_useHi_24 ? _canSkipShift_T_190 : _canSkipShift_T_216; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_218 = {canSkipShift_useHi_24,_canSkipShift_T_217}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_219 = canSkipShift_useHi_16 ? _canSkipShift_T_164 : _canSkipShift_T_218; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_220 = {canSkipShift_useHi_16,_canSkipShift_T_219}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _canSkipShift_T_221 = canSkipShift_useHi_15 ? 6'h0 : _canSkipShift_T_220; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [6:0] _canSkipShift_T_222 = {canSkipShift_useHi_15,_canSkipShift_T_221}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] canSkipShift = _canSkipShift_T_110 - _canSkipShift_T_222; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:45]
  wire [6:0] _value_T_1 = canSkipShift >= 7'h3f ? 7'h3f : canSkipShift; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:21]
  wire  line_387_clock;
  wire  line_387_reset;
  wire  line_387_valid;
  reg  line_387_valid_reg;
  wire  _T_5 = state == 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:22]
  wire  line_388_clock;
  wire  line_388_reset;
  wire  line_388_valid;
  reg  line_388_valid_reg;
  wire [127:0] _GEN_14 = {{63'd0}, aValx2Reg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [127:0] _shiftReg_T = _GEN_14 << cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire  line_389_clock;
  wire  line_389_reset;
  wire  line_389_valid;
  reg  line_389_valid_reg;
  wire  _T_6 = state == 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:22]
  wire  line_390_clock;
  wire  line_390_reset;
  wire  line_390_valid;
  reg  line_390_valid_reg;
  wire [64:0] _GEN_33 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire  enough = hi >= _GEN_33; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire [64:0] _shiftReg_T_2 = hi - _GEN_33; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_3 = enough ? _shiftReg_T_2 : hi; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:24]
  wire [128:0] _shiftReg_T_5 = {_shiftReg_T_3[63:0],lo,enough}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:20]
  wire  wrap = cnt_value == 6'h3f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [5:0] _value_T_4 = cnt_value + 6'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_391_clock;
  wire  line_391_reset;
  wire  line_391_valid;
  reg  line_391_valid_reg;
  wire [2:0] _GEN_18 = wrap ? 3'h4 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 118:{36,44} 77:22]
  wire  line_392_clock;
  wire  line_392_reset;
  wire  line_392_valid;
  reg  line_392_valid_reg;
  wire  _T_8 = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:22]
  wire  line_393_clock;
  wire  line_393_reset;
  wire  line_393_valid;
  reg  line_393_valid_reg;
  wire [2:0] _GEN_19 = state == 3'h4 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_21 = state == 3'h3 ? _value_T_4 : cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_22 = state == 3'h3 ? _GEN_18 : _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
  wire [5:0] _GEN_25 = state == 3'h2 ? cnt_value : _GEN_21; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [6:0] _GEN_26 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_25}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:15 97:34]
  wire [6:0] _GEN_30 = newReq ? {{1'd0}, cnt_value} : _GEN_26; // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] r = hi[64:1]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 123:13]
  wire [63:0] _resQ_T_1 = 64'h0 - lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _resQ_T_1 : lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:17]
  wire [63:0] _resR_T_1 = 64'h0 - r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _resR_T_1 : r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:17]
  wire [6:0] _GEN_35 = reset ? 7'h0 : _GEN_30; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  GEN_w1_line #(.COVER_INDEX(380)) line_380 (
    .clock(line_380_clock),
    .reset(line_380_reset),
    .valid(line_380_valid)
  );
  GEN_w1_line #(.COVER_INDEX(381)) line_381 (
    .clock(line_381_clock),
    .reset(line_381_reset),
    .valid(line_381_valid)
  );
  GEN_w1_line #(.COVER_INDEX(382)) line_382 (
    .clock(line_382_clock),
    .reset(line_382_reset),
    .valid(line_382_valid)
  );
  GEN_w1_line #(.COVER_INDEX(383)) line_383 (
    .clock(line_383_clock),
    .reset(line_383_reset),
    .valid(line_383_valid)
  );
  GEN_w1_line #(.COVER_INDEX(384)) line_384 (
    .clock(line_384_clock),
    .reset(line_384_reset),
    .valid(line_384_valid)
  );
  GEN_w1_line #(.COVER_INDEX(385)) line_385 (
    .clock(line_385_clock),
    .reset(line_385_reset),
    .valid(line_385_valid)
  );
  GEN_w1_line #(.COVER_INDEX(386)) line_386 (
    .clock(line_386_clock),
    .reset(line_386_reset),
    .valid(line_386_valid)
  );
  GEN_w1_line #(.COVER_INDEX(387)) line_387 (
    .clock(line_387_clock),
    .reset(line_387_reset),
    .valid(line_387_valid)
  );
  GEN_w1_line #(.COVER_INDEX(388)) line_388 (
    .clock(line_388_clock),
    .reset(line_388_reset),
    .valid(line_388_valid)
  );
  GEN_w1_line #(.COVER_INDEX(389)) line_389 (
    .clock(line_389_clock),
    .reset(line_389_reset),
    .valid(line_389_valid)
  );
  GEN_w1_line #(.COVER_INDEX(390)) line_390 (
    .clock(line_390_clock),
    .reset(line_390_reset),
    .valid(line_390_valid)
  );
  GEN_w1_line #(.COVER_INDEX(391)) line_391 (
    .clock(line_391_clock),
    .reset(line_391_reset),
    .valid(line_391_valid)
  );
  GEN_w1_line #(.COVER_INDEX(392)) line_392 (
    .clock(line_392_clock),
    .reset(line_392_reset),
    .valid(line_392_valid)
  );
  GEN_w1_line #(.COVER_INDEX(393)) line_393 (
    .clock(line_393_clock),
    .reset(line_393_reset),
    .valid(line_393_valid)
  );
  assign line_380_clock = clock;
  assign line_380_reset = reset;
  assign line_380_valid = newReq ^ line_380_valid_reg;
  assign line_381_clock = clock;
  assign line_381_reset = reset;
  assign line_381_valid = newReq ^ line_381_valid_reg;
  assign line_382_clock = clock;
  assign line_382_reset = reset;
  assign line_382_valid = newReq ^ line_382_valid_reg;
  assign line_383_clock = clock;
  assign line_383_reset = reset;
  assign line_383_valid = newReq ^ line_383_valid_reg;
  assign line_384_clock = clock;
  assign line_384_reset = reset;
  assign line_384_valid = newReq ^ line_384_valid_reg;
  assign line_385_clock = clock;
  assign line_385_reset = reset;
  assign line_385_valid = newReq ^ line_385_valid_reg;
  assign line_386_clock = clock;
  assign line_386_reset = reset;
  assign line_386_valid = _T_4 ^ line_386_valid_reg;
  assign line_387_clock = clock;
  assign line_387_reset = reset;
  assign line_387_valid = _T_4 ^ line_387_valid_reg;
  assign line_388_clock = clock;
  assign line_388_reset = reset;
  assign line_388_valid = _T_5 ^ line_388_valid_reg;
  assign line_389_clock = clock;
  assign line_389_reset = reset;
  assign line_389_valid = _T_5 ^ line_389_valid_reg;
  assign line_390_clock = clock;
  assign line_390_reset = reset;
  assign line_390_valid = _T_6 ^ line_390_valid_reg;
  assign line_391_clock = clock;
  assign line_391_reset = reset;
  assign line_391_valid = wrap ^ line_391_valid_reg;
  assign line_392_clock = clock;
  assign line_392_reset = reset;
  assign line_392_valid = _T_6 ^ line_392_valid_reg;
  assign line_393_clock = clock;
  assign line_393_reset = reset;
  assign line_393_valid = _T_8 ^ line_393_valid_reg;
  assign io_in_ready = state == 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 126:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end else if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      state <= 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
      state <= 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
      state <= 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 113:11]
    end else begin
      state <= _GEN_22;
    end
    if (!(newReq)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
        if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
          shiftReg <= {{1'd0}, _shiftReg_T}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
          shiftReg <= _shiftReg_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
      aSignReg <= aSign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    line_380_valid_reg <= newReq;
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
      qSignReg <= (aSign ^ bSign) & ~divBy0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    line_381_valid_reg <= newReq;
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
      if (bSign) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
        bReg <= _T_3;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    line_382_valid_reg <= newReq;
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
      aValx2Reg <= _aValx2Reg_T; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    line_383_valid_reg <= newReq;
    cnt_value <= _GEN_35[5:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    line_384_valid_reg <= newReq;
    line_385_valid_reg <= newReq;
    line_386_valid_reg <= _T_4;
    line_387_valid_reg <= _T_4;
    line_388_valid_reg <= _T_5;
    line_389_valid_reg <= _T_5;
    line_390_valid_reg <= _T_6;
    line_391_valid_reg <= wrap;
    line_392_valid_reg <= _T_6;
    line_393_valid_reg <= _T_8;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_380_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  qSignReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_381_valid_reg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  bReg = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  line_382_valid_reg = _RAND_7[0:0];
  _RAND_8 = {3{`RANDOM}};
  aValx2Reg = _RAND_8[64:0];
  _RAND_9 = {1{`RANDOM}};
  line_383_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cnt_value = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  line_384_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_385_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_386_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_387_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_388_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_389_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_390_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_391_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_392_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_393_valid_reg = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (newReq) begin
      cover(1'h1);
    end
    //
    if (newReq) begin
      cover(1'h1);
    end
    //
    if (newReq) begin
      cover(1'h1);
    end
    //
    if (newReq) begin
      cover(1'h1);
    end
    //
    if (newReq) begin
      cover(1'h1);
    end
    //
    if (~newReq) begin
      cover(1'h1);
    end
    //
    if (~newReq & _T_4) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & _T_5) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & ~_T_5) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & ~_T_5 & _T_6) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & ~_T_5 & _T_6 & wrap) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & ~_T_5 & ~_T_6) begin
      cover(1'h1);
    end
    //
    if (~newReq & ~_T_4 & ~_T_5 & ~_T_6 & _T_8) begin
      cover(1'h1);
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output [63:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  div_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 43:25]
  wire [64:0] _mul_io_in_bits_0_T_1 = {1'h0,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_0_signBit = io_in_bits_src1[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_0_T_2 = {mul_io_in_bits_0_signBit,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _mul_io_in_bits_0_T_5 = 2'h0 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_6 = 2'h1 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_7 = 2'h2 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_8 = 2'h3 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [64:0] _mul_io_in_bits_0_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_13 = _mul_io_in_bits_0_T_9 | _mul_io_in_bits_0_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_14 = _mul_io_in_bits_0_T_13 | _mul_io_in_bits_0_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_1 = {1'h0,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_1_signBit = io_in_bits_src2[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_1_T_2 = {mul_io_in_bits_1_signBit,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] _mul_io_in_bits_1_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_1_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_13 = _mul_io_in_bits_1_T_9 | _mul_io_in_bits_1_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_14 = _mul_io_in_bits_1_T_13 | _mul_io_in_bits_1_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  div_io_in_bits_0_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_0_T_1 = div_io_in_bits_0_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_0_T_2 = {_div_io_in_bits_0_T_1,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_0_T_4 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_0_T_5 = isDivSign ? _div_io_in_bits_0_T_2 : _div_io_in_bits_0_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire  div_io_in_bits_1_signBit = io_in_bits_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_1_T_1 = div_io_in_bits_1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_1_T_2 = {_div_io_in_bits_1_T_1,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_1_T_4 = {32'h0,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_1_T_5 = isDivSign ? _div_io_in_bits_1_T_2 : _div_io_in_bits_1_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[src/main/scala/nutcore/backend/fu/MDU.scala 178:16]
  wire  io_out_bits_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _io_out_bits_T_1 = io_out_bits_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_T_2 = {_io_out_bits_T_1,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
  wire  isDivReg = _isDivReg_T ? isDiv : isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:21]
  wire  _T = mul_io_out_ready & mul_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  Multiplier mul ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 183:22]
  assign io_out_bits = isW ? _io_out_bits_T_2 : res; // @[src/main/scala/nutcore/backend/fu/MDU.scala 179:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 173:34]
  assign mul_io_in_bits_0 = _mul_io_in_bits_0_T_14 | _mul_io_in_bits_0_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_in_bits_1 = _mul_io_in_bits_1_T_14 | _mul_io_in_bits_1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _div_io_in_bits_0_T_5 : io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _div_io_in_bits_1_T_5 : io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  always @(posedge clock) begin
    isDivReg_REG <= io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg_REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DummyDPICWrapper_1(
  input         clock,
  input         reset,
  input  [63:0] io_bits_privilegeMode, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mcause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_scause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_satp, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mie, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mideleg, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_medeleg // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mcause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_scause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_satp; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mie; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mideleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_medeleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestCSRState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_privilegeMode(dpic_io_privilegeMode),
    .io_mstatus(dpic_io_mstatus),
    .io_sstatus(dpic_io_sstatus),
    .io_mepc(dpic_io_mepc),
    .io_sepc(dpic_io_sepc),
    .io_mtval(dpic_io_mtval),
    .io_stval(dpic_io_stval),
    .io_mtvec(dpic_io_mtvec),
    .io_stvec(dpic_io_stvec),
    .io_mcause(dpic_io_mcause),
    .io_scause(dpic_io_scause),
    .io_satp(dpic_io_satp),
    .io_mip(dpic_io_mip),
    .io_mie(dpic_io_mie),
    .io_mscratch(dpic_io_mscratch),
    .io_sscratch(dpic_io_sscratch),
    .io_mideleg(dpic_io_mideleg),
    .io_medeleg(dpic_io_medeleg),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_privilegeMode = io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mstatus = io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sstatus = io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mepc = io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sepc = io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtval = io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stval = io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtvec = io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stvec = io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mcause = io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_scause = io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_satp = io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mip = io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mie = io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mscratch = io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sscratch = io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mideleg = io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_medeleg = io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DummyDPICWrapper_2(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_interrupt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exception, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_exceptionPC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exceptionInst // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_interrupt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exception; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_interrupt(dpic_io_interrupt),
    .io_exception(dpic_io_exception),
    .io_exceptionPC(dpic_io_exceptionPC),
    .io_exceptionInst(dpic_io_exceptionInst),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_interrupt = io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exception = io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionPC = io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionInst = io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module CSRDiffWrapper(
  input         clock,
  input         reset,
  input  [63:0] io_csrState_privilegeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mtval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_stval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mtvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_stvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mcause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_scause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_satp, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mip, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mie, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mideleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_medeleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input         io_archEvent_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_interrupt, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_exception, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_archEvent_exceptionPC, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_exceptionInst // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftestArchEvent_module_io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] difftest_REG_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg  difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [63:0] difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg  difftestArchEvent_REG_1_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [63:0] difftestArchEvent_REG_1_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  DummyDPICWrapper_1 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_privilegeMode(difftest_module_io_bits_privilegeMode),
    .io_bits_mstatus(difftest_module_io_bits_mstatus),
    .io_bits_sstatus(difftest_module_io_bits_sstatus),
    .io_bits_mepc(difftest_module_io_bits_mepc),
    .io_bits_sepc(difftest_module_io_bits_sepc),
    .io_bits_mtval(difftest_module_io_bits_mtval),
    .io_bits_stval(difftest_module_io_bits_stval),
    .io_bits_mtvec(difftest_module_io_bits_mtvec),
    .io_bits_stvec(difftest_module_io_bits_stvec),
    .io_bits_mcause(difftest_module_io_bits_mcause),
    .io_bits_scause(difftest_module_io_bits_scause),
    .io_bits_satp(difftest_module_io_bits_satp),
    .io_bits_mip(difftest_module_io_bits_mip),
    .io_bits_mie(difftest_module_io_bits_mie),
    .io_bits_mscratch(difftest_module_io_bits_mscratch),
    .io_bits_sscratch(difftest_module_io_bits_sscratch),
    .io_bits_mideleg(difftest_module_io_bits_mideleg),
    .io_bits_medeleg(difftest_module_io_bits_medeleg)
  );
  DummyDPICWrapper_2 difftestArchEvent_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftestArchEvent_module_clock),
    .reset(difftestArchEvent_module_reset),
    .io_valid(difftestArchEvent_module_io_valid),
    .io_bits_valid(difftestArchEvent_module_io_bits_valid),
    .io_bits_interrupt(difftestArchEvent_module_io_bits_interrupt),
    .io_bits_exception(difftestArchEvent_module_io_bits_exception),
    .io_bits_exceptionPC(difftestArchEvent_module_io_bits_exceptionPC),
    .io_bits_exceptionInst(difftestArchEvent_module_io_bits_exceptionInst)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_privilegeMode = difftest_REG_privilegeMode; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mstatus = difftest_REG_mstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sstatus = difftest_REG_sstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mepc = difftest_REG_mepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sepc = difftest_REG_sepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mtval = difftest_REG_mtval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_stval = difftest_REG_stval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mtvec = difftest_REG_mtvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_stvec = difftest_REG_stvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mcause = difftest_REG_mcause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_scause = difftest_REG_scause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_satp = difftest_REG_satp; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mip = difftest_REG_mip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mie = difftest_REG_mie; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mscratch = difftest_REG_mscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sscratch = difftest_REG_sscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mideleg = difftest_REG_mideleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_medeleg = difftest_REG_medeleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftestArchEvent_module_clock = clock;
  assign difftestArchEvent_module_reset = reset;
  assign difftestArchEvent_module_io_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_interrupt = difftestArchEvent_REG_1_interrupt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exception = difftestArchEvent_REG_1_exception; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exceptionPC = difftestArchEvent_REG_1_exceptionPC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exceptionInst = difftestArchEvent_REG_1_exceptionInst; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  always @(posedge clock) begin
    difftest_REG_privilegeMode <= io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mstatus <= io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sstatus <= io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mepc <= io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sepc <= io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mtval <= io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_stval <= io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mtvec <= io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_stvec <= io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mcause <= io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_scause <= io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_satp <= io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mip <= io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mie <= io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mscratch <= io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sscratch <= io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mideleg <= io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_medeleg <= io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftestArchEvent_REG_valid <= io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_interrupt <= io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exception <= io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exceptionPC <= io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exceptionInst <= io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_1_valid <= difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_interrupt <= difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exception <= difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exceptionPC <= difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exceptionInst <= difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_REG_privilegeMode = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  difftest_REG_mstatus = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_sstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  difftest_REG_mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  difftest_REG_sepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  difftest_REG_mtval = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_stval = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  difftest_REG_mtvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  difftest_REG_stvec = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  difftest_REG_mcause = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  difftest_REG_scause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  difftest_REG_satp = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  difftest_REG_mip = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  difftest_REG_mie = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  difftest_REG_mscratch = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  difftest_REG_sscratch = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  difftest_REG_mideleg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  difftest_REG_medeleg = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  difftestArchEvent_REG_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  difftestArchEvent_REG_interrupt = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  difftestArchEvent_REG_exception = _RAND_20[31:0];
  _RAND_21 = {2{`RANDOM}};
  difftestArchEvent_REG_exceptionPC = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  difftestArchEvent_REG_exceptionInst = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  difftestArchEvent_REG_1_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  difftestArchEvent_REG_1_interrupt = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exception = _RAND_25[31:0];
  _RAND_26 = {2{`RANDOM}};
  difftestArchEvent_REG_1_exceptionPC = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exceptionInst = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_12, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_13, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_15, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_3, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_9, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_11, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_crossBoundaryFault, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_instrValid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_illegalJump_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_illegalJump_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_dmemExceptionAddr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_xretIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_xretIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_xretIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_imemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_dmemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_sum, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_mxr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_loadPF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_storePF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_laf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_saf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wenFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isPerfRead, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isExit, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_vmEnable, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_rfWenReal, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         set_lr,
  output        lr_0,
  input         meip_0,
  output [63:0] lrAddr_0,
  output [63:0] satp_0,
  input         mtip_0,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [11:0] intrVecIDU_0,
  input  [63:0] set_lr_addr,
  input         msip_0,
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
`endif // RANDOMIZE_REG_INIT
  wire  CSRDiffWrapper_clock; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire  CSRDiffWrapper_reset; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire  CSRDiffWrapper_io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  reg [1:0] priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
  reg [63:0] mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
  reg [63:0] mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
  reg [63:0] mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
  reg [63:0] mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
  reg [63:0] mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
  reg [63:0] mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
  reg [63:0] mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
  wire [11:0] _mip_T = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:22]
  wire [63:0] _GEN_142 = {{52'd0}, _mip_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire [63:0] _mip_T_1 = _GEN_142 | mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire  mip_s_u = _mip_T_1[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_s = _mip_T_1[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_h = _mip_T_1[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_m = _mip_T_1[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_u = _mip_T_1[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_s = _mip_T_1[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_h = _mip_T_1[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_m = _mip_T_1[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_u = _mip_T_1[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_s = _mip_T_1[9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_h = _mip_T_1[10]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_m = _mip_T_1[11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  reg [63:0] mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  reg [63:0] medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
  reg [63:0] mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
  reg [63:0] mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
  reg [63:0] stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 379:32]
  reg [63:0] satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
  wire [3:0] satpStruct_mode = satp[63:60]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 384:33]
  wire  _vmEnable_T_1 = priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:38]
  wire  vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  reg [63:0] sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
  reg [63:0] scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
  reg [63:0] stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
  reg [63:0] sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
  reg [63:0] scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
  reg  lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
  reg [63:0] lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
  wire  line_394_clock;
  wire  line_394_reset;
  wire  line_394_valid;
  reg  line_394_valid_reg;
  reg [63:0] perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [5:0] lo = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] _T_25 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 507:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdata_T_29 = 12'hf12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_30 = 12'h180 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_59 = _rdata_T_30 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_31 = 12'h140 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_60 = _rdata_T_31 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_88 = _rdata_T_59 | _rdata_T_60; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_32 = 12'h306 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_61 = _rdata_T_32 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_89 = _rdata_T_88 | _rdata_T_61; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_33 = 12'hf11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_34 = 12'h104 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_5 = mie & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_63 = _rdata_T_34 ? _rdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_91 = _rdata_T_89 | _rdata_T_63; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_35 = 12'h144 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _GEN_143 = {{52'd0}, _T_25}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_6 = _GEN_143 & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_64 = _rdata_T_35 ? _rdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_92 = _rdata_T_91 | _rdata_T_64; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_36 = 12'h100 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_7 = mstatus & 64'h80000003000d8122; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_65 = _rdata_T_36 ? _rdata_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_93 = _rdata_T_92 | _rdata_T_65; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_37 = 12'h305 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_66 = _rdata_T_37 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_94 = _rdata_T_93 | _rdata_T_66; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_38 = 12'h300 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_9 = mstatus & 64'h8000000f007ff9aa; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_67 = _rdata_T_38 ? _rdata_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_95 = _rdata_T_94 | _rdata_T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_39 = 12'hf13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_40 = 12'h340 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_69 = _rdata_T_40 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_97 = _rdata_T_95 | _rdata_T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_41 = 12'h142 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_70 = _rdata_T_41 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_98 = _rdata_T_97 | _rdata_T_70; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_42 = 12'h302 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_71 = _rdata_T_42 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_99 = _rdata_T_98 | _rdata_T_71; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_43 = 12'h105 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_72 = _rdata_T_43 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_100 = _rdata_T_99 | _rdata_T_72; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_44 = 12'h141 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_73 = _rdata_T_44 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_101 = _rdata_T_100 | _rdata_T_73; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_45 = 12'h342 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_74 = _rdata_T_45 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_102 = _rdata_T_101 | _rdata_T_74; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_46 = 12'h304 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_75 = _rdata_T_46 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_103 = _rdata_T_102 | _rdata_T_75; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_47 = 12'hb01 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_76 = _rdata_T_47 ? perfCnts_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_104 = _rdata_T_103 | _rdata_T_76; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_48 = 12'h143 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_77 = _rdata_T_48 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_105 = _rdata_T_104 | _rdata_T_77; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_49 = 12'h301 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_78 = _rdata_T_49 ? 64'h8000000000141105 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_106 = _rdata_T_105 | _rdata_T_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_50 = 12'hb00 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_79 = _rdata_T_50 ? perfCnts_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_107 = _rdata_T_106 | _rdata_T_79; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_51 = 12'h344 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_80 = _rdata_T_51 ? _GEN_143 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_108 = _rdata_T_107 | _rdata_T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_52 = 12'hb02 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_81 = _rdata_T_52 ? perfCnts_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_109 = _rdata_T_108 | _rdata_T_81; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_53 = 12'h303 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_82 = _rdata_T_53 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_110 = _rdata_T_109 | _rdata_T_82; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_54 = 12'hf14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_55 = 12'h341 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_84 = _rdata_T_55 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_112 = _rdata_T_110 | _rdata_T_84; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_56 = 12'h343 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_85 = _rdata_T_56 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_85; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_57 = 12'h106 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_86 = _rdata_T_57 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 512:30]
  wire [63:0] _wdata_T_1 = ~io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:33]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:30]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 515:30]
  wire [63:0] _wdata_T_4 = ~csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:33]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:30]
  wire  _wdata_T_6 = 7'h1 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_7 = 7'h2 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_8 = 7'h3 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_9 = 7'h5 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_10 = 7'h6 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_11 = 7'h7 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_in_bits_src1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 522:69]
  wire [7:0] wen_lo = {io_cfIn_exceptionVec_7,io_cfIn_exceptionVec_6,io_cfIn_exceptionVec_5,io_cfIn_exceptionVec_4,1'h0,
    io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire [15:0] _wen_T = {io_cfIn_exceptionVec_15,1'h0,io_cfIn_exceptionVec_13,io_cfIn_exceptionVec_12,4'h0,wen_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire  _wen_T_2 = ~(|_wen_T); // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:23]
  wire  _wen_T_4 = io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:64]
  wire  wen = io_in_valid & ~(|_wen_T) & io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:56]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 526:39]
  wire  isCSRRS = io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 531:40]
  wire  isCSRRC = io_in_bits_func == 7'h3 | io_in_bits_func == 7'h7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 532:40]
  wire  noWriteSideEffect = (isCSRRS | isCSRRC) & io_cfIn_instr[19:15] == 5'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 533:48]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~noWriteSideEffect; // @[src/main/scala/nutcore/backend/fu/CSR.scala 535:58]
  wire  _tvm_T_1 = priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:57]
  wire  tvm = mstatusStruct_tvm & priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:39]
  wire  _io_sfence_vma_invalid_T = priviledgeMode == 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:43]
  wire  _isIllegalTVM_T_1 = addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:42]
  wire  isIllegalTVM = tvm & wen & addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:34]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite | isIllegalTVM; // @[src/main/scala/nutcore/backend/fu/CSR.scala 544:57]
  wire  _canWriteCSR_T = ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:28]
  wire  _canWriteCSR_T_1 = wen & ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:25]
  wire  canWriteCSR = wen & ~isIllegalAccess & (addr != 12'h180 | satpLegalMode); // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:45]
  wire  _T_48 = canWriteCSR & _isIllegalTVM_T_1; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_395_clock;
  wire  line_395_reset;
  wire  line_395_valid;
  reg  line_395_valid_reg;
  wire [63:0] _satp_T = wdata & 64'h8ffff000000fffff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _satp_T_2 = satp & 64'h70000ffffff00000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _satp_T_3 = _satp_T | _satp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_50 = canWriteCSR & addr == 12'h140; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_396_clock;
  wire  line_396_reset;
  wire  line_396_valid;
  reg  line_396_valid_reg;
  wire  _T_52 = canWriteCSR & addr == 12'h306; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_397_clock;
  wire  line_397_reset;
  wire  line_397_valid;
  reg  line_397_valid_reg;
  wire  _T_54 = canWriteCSR & addr == 12'h104; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_398_clock;
  wire  line_398_reset;
  wire  line_398_valid;
  reg  line_398_valid_reg;
  wire [63:0] _mie_T = wdata & sieMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_1 = ~sieMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _mie_T_2 = mie & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_56 = canWriteCSR & addr == 12'h100; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_399_clock;
  wire  line_399_reset;
  wire  line_399_valid;
  reg  line_399_valid_reg;
  wire [63:0] _mstatus_T = wdata & 64'hc0122; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_2 = mstatus & 64'hfffffffffff3fedd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_3 = _mstatus_T | _mstatus_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_mpp = _mstatus_T_3[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_3[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix = mstatus_mstatusOld_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_3[62:13],mstatus_mppFix,_mstatus_T_3[10:0]}
    ; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_63 = canWriteCSR & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_58 = canWriteCSR & addr == 12'h305; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_400_clock;
  wire  line_400_reset;
  wire  line_400_valid;
  reg  line_400_valid_reg;
  wire [63:0] _mtvec_T = wdata & 64'hfffffffffffffffc; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mtvec_T_2 = mtvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtvec_T_3 = _mtvec_T | _mtvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_60 = canWriteCSR & addr == 12'h300; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_401_clock;
  wire  line_401_reset;
  wire  line_401_valid;
  reg  line_401_valid_reg;
  wire [63:0] _mstatus_T_4 = wdata & 64'h80000000007e19aa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_6 = mstatus & 64'h7fffffffff81e655; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_7 = _mstatus_T_4 | _mstatus_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_1_mpp = _mstatus_T_7[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_1_fs = _mstatus_T_7[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix_1 = mstatus_mstatusOld_1_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_1_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew_1 = {mstatus_mstatusOld_1_fs == 2'h3,_mstatus_T_7[62:13],mstatus_mppFix_1,_mstatus_T_7[
    10:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_65 = canWriteCSR & addr == 12'h300 ? mstatus_mstatusNew_1 : _GEN_63; // @[src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_62 = canWriteCSR & addr == 12'h340; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_402_clock;
  wire  line_402_reset;
  wire  line_402_valid;
  reg  line_402_valid_reg;
  wire  _T_64 = canWriteCSR & addr == 12'h142; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_403_clock;
  wire  line_403_reset;
  wire  line_403_valid;
  reg  line_403_valid_reg;
  wire [63:0] _GEN_67 = canWriteCSR & addr == 12'h142 ? wdata : scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_65 = addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_66 = canWriteCSR & addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_404_clock;
  wire  line_404_reset;
  wire  line_404_valid;
  reg  line_404_valid_reg;
  wire [63:0] _medeleg_T = wdata & 64'hb3ff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'hffffffffffff4c00; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_68 = canWriteCSR & addr == 12'h105; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_405_clock;
  wire  line_405_reset;
  wire  line_405_valid;
  reg  line_405_valid_reg;
  wire [63:0] _stvec_T_2 = stvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _stvec_T_3 = _mtvec_T | _stvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_70 = canWriteCSR & addr == 12'h141; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_406_clock;
  wire  line_406_reset;
  wire  line_406_valid;
  reg  line_406_valid_reg;
  wire [63:0] _sepc_T = wdata & 64'hfffffffffffffffe; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _sepc_T_2 = sepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _sepc_T_3 = _sepc_T | _sepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_70 = canWriteCSR & addr == 12'h141 ? _sepc_T_3 : sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_72 = canWriteCSR & addr == 12'h342; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_407_clock;
  wire  line_407_reset;
  wire  line_407_valid;
  reg  line_407_valid_reg;
  wire [63:0] _GEN_71 = canWriteCSR & addr == 12'h342 ? wdata : mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_74 = canWriteCSR & addr == 12'h304; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_408_clock;
  wire  line_408_reset;
  wire  line_408_valid;
  reg  line_408_valid_reg;
  wire [63:0] _mie_T_4 = wdata & 64'haaa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_6 = mie & 64'hfffffffffffff555; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_7 = _mie_T_4 | _mie_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_76 = canWriteCSR & addr == 12'hb01; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_409_clock;
  wire  line_409_reset;
  wire  line_409_valid;
  reg  line_409_valid_reg;
  wire  _T_78 = canWriteCSR & addr == 12'h143; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_410_clock;
  wire  line_410_reset;
  wire  line_410_valid;
  reg  line_410_valid_reg;
  wire [63:0] _GEN_74 = canWriteCSR & addr == 12'h143 ? wdata : stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_79 = addr == 12'hb00; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_80 = canWriteCSR & addr == 12'hb00; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_411_clock;
  wire  line_411_reset;
  wire  line_411_valid;
  reg  line_411_valid_reg;
  wire  _T_81 = addr == 12'hb02; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_82 = canWriteCSR & addr == 12'hb02; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_412_clock;
  wire  line_412_reset;
  wire  line_412_valid;
  reg  line_412_valid_reg;
  wire  _T_84 = canWriteCSR & addr == 12'h303; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_413_clock;
  wire  line_413_reset;
  wire  line_413_valid;
  reg  line_413_valid_reg;
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'hfffffffffffffddd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_86 = canWriteCSR & addr == 12'h341; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_414_clock;
  wire  line_414_reset;
  wire  line_414_valid;
  reg  line_414_valid_reg;
  wire [63:0] _mepc_T_2 = mepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mepc_T_3 = _sepc_T | _mepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_78 = canWriteCSR & addr == 12'h341 ? _mepc_T_3 : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_88 = canWriteCSR & addr == 12'h343; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_415_clock;
  wire  line_415_reset;
  wire  line_415_valid;
  reg  line_415_valid_reg;
  wire [63:0] _GEN_79 = canWriteCSR & addr == 12'h343 ? wdata : mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_90 = canWriteCSR & addr == 12'h106; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_416_clock;
  wire  line_416_reset;
  wire  line_416_valid;
  reg  line_416_valid_reg;
  wire  _isIllegalAddr_illegalAddr_T_1 = _rdata_T_29 ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_3 = _rdata_T_30 ? 1'h0 : _isIllegalAddr_illegalAddr_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_5 = _rdata_T_31 ? 1'h0 : _isIllegalAddr_illegalAddr_T_3; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_7 = _rdata_T_32 ? 1'h0 : _isIllegalAddr_illegalAddr_T_5; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_9 = _rdata_T_33 ? 1'h0 : _isIllegalAddr_illegalAddr_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_11 = _rdata_T_34 ? 1'h0 : _isIllegalAddr_illegalAddr_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_13 = _rdata_T_35 ? 1'h0 : _isIllegalAddr_illegalAddr_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_15 = _rdata_T_36 ? 1'h0 : _isIllegalAddr_illegalAddr_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_17 = _rdata_T_37 ? 1'h0 : _isIllegalAddr_illegalAddr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_19 = _rdata_T_38 ? 1'h0 : _isIllegalAddr_illegalAddr_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_21 = _rdata_T_39 ? 1'h0 : _isIllegalAddr_illegalAddr_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_23 = _rdata_T_40 ? 1'h0 : _isIllegalAddr_illegalAddr_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_25 = _rdata_T_41 ? 1'h0 : _isIllegalAddr_illegalAddr_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_27 = _rdata_T_42 ? 1'h0 : _isIllegalAddr_illegalAddr_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_29 = _rdata_T_43 ? 1'h0 : _isIllegalAddr_illegalAddr_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_31 = _rdata_T_44 ? 1'h0 : _isIllegalAddr_illegalAddr_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_33 = _rdata_T_45 ? 1'h0 : _isIllegalAddr_illegalAddr_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_35 = _rdata_T_46 ? 1'h0 : _isIllegalAddr_illegalAddr_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_37 = _rdata_T_47 ? 1'h0 : _isIllegalAddr_illegalAddr_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_39 = _rdata_T_48 ? 1'h0 : _isIllegalAddr_illegalAddr_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_41 = _rdata_T_49 ? 1'h0 : _isIllegalAddr_illegalAddr_T_39; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_43 = _rdata_T_50 ? 1'h0 : _isIllegalAddr_illegalAddr_T_41; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_45 = _rdata_T_51 ? 1'h0 : _isIllegalAddr_illegalAddr_T_43; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_47 = _rdata_T_52 ? 1'h0 : _isIllegalAddr_illegalAddr_T_45; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_49 = _rdata_T_53 ? 1'h0 : _isIllegalAddr_illegalAddr_T_47; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_51 = _rdata_T_54 ? 1'h0 : _isIllegalAddr_illegalAddr_T_49; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_53 = _rdata_T_55 ? 1'h0 : _isIllegalAddr_illegalAddr_T_51; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_55 = _rdata_T_56 ? 1'h0 : _isIllegalAddr_illegalAddr_T_53; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  isIllegalAddr = _rdata_T_57 ? 1'h0 : _isIllegalAddr_illegalAddr_T_55; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  resetSatp = _isIllegalTVM_T_1 & wen & _canWriteCSR_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 552:42]
  wire  _io_isExit_T = addr == 12'h344; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:38]
  wire  _io_isExit_T_1 = addr == 12'h144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:56]
  wire  _io_isExit_T_9 = _canWriteCSR_T_1 | ~wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:30]
  wire  _io_isExit_T_10 = io_out_valid & (addr == 12'h344 | addr == 12'h144) & _wen_T_4 & _io_isExit_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:93]
  wire  _T_95 = _canWriteCSR_T_1 & _io_isExit_T; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_417_clock;
  wire  line_417_reset;
  wire  line_417_valid;
  reg  line_417_valid_reg;
  wire [63:0] _mipReg_T = wdata & 64'h77f; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mipReg_T_2 = mipReg & 64'hfffffffffffff880; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_3 = _mipReg_T | _mipReg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_97 = _canWriteCSR_T_1 & _io_isExit_T_1; // @[src/main/scala/utils/RegMap.scala 50:56]
  wire  line_418_clock;
  wire  line_418_reset;
  wire  line_418_valid;
  reg  line_418_valid_reg;
  wire [63:0] _mipReg_T_6 = mipReg & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_7 = _mie_T | _mipReg_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _isEbreak_T_1 = io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:90]
  wire  isEcall = addr == 12'h0 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 569:88]
  wire  isMret = _T_65 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 570:88]
  wire  isSret = addr == 12'h102 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 571:88]
  wire  isUret = addr == 12'h2 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 572:88]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:63]
  wire  hasInstrAccessFault = io_cfIn_exceptionVec_1 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 633:67]
  wire  hasLoadPageFault = io_dmemMMU_loadPF | io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 634:43]
  wire  hasStorePageFault = io_dmemMMU_storePF | io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:45]
  wire  hasLoadAccessFault = io_dmemMMU_laf | io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 636:42]
  wire  hasStoreAccessFault = io_dmemMMU_saf | io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 637:43]
  wire [38:0] _imemExceptionAddr_T_1 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 644:42]
  wire  imemExceptionAddr_signBit = _imemExceptionAddr_T_1[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_2 = imemExceptionAddr_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_3 = {_imemExceptionAddr_T_2,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_6 = {25'h0,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_7 = vmEnable ? _imemExceptionAddr_T_3 : _imemExceptionAddr_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 644:12]
  wire  imemExceptionAddr_signBit_1 = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_8 = imemExceptionAddr_signBit_1 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_9 = {_imemExceptionAddr_T_8,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_10 = {25'h0,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_11 = vmEnable ? _imemExceptionAddr_T_9 : _imemExceptionAddr_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 645:12]
  wire [63:0] _imemExceptionAddr_T_12 = io_cfIn_crossBoundaryFault ? _imemExceptionAddr_T_7 : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:10]
  wire [63:0] imemExceptionAddr = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_12; // @[src/main/scala/nutcore/backend/fu/CSR.scala 641:29]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:31]
  wire [11:0] _ideleg_T = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:41]
  wire [63:0] _GEN_144 = {{52'd0}, _ideleg_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
  wire [63:0] ideleg = mideleg & _GEN_144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
  wire  _intrVecEnable_0_T_2 = priviledgeMode < 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:125]
  wire  _intrVecEnable_0_T_4 = priviledgeMode == 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 676:53]
  wire  _intrVecEnable_0_T_7 = priviledgeMode == 2'h3 & mstatusStruct_ie_m | _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 676:87]
  wire  intrVecEnable_0 = ideleg[0] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_1 = ideleg[1] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_2 = ideleg[2] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_3 = ideleg[3] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_4 = ideleg[4] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_5 = ideleg[5] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_6 = ideleg[6] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_7 = ideleg[7] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_8 = ideleg[8] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_9 = ideleg[9] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_10 = ideleg[10] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_11 = ideleg[11] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _ideleg_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:27]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:65]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:65]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:49]
  wire [5:0] intrVecIDU_lo = {intrVec[5],1'h0,intrVec[3],1'h0,intrVec[1],1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:100]
  wire [11:0] intrVecIDU = {intrVec[11],1'h0,intrVec[9],1'h0,intrVec[7],1'h0,intrVecIDU_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:100]
  wire [2:0] _intrNO_T = io_cfIn_intrVec_5 ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_1 = io_cfIn_intrVec_9 ? 4'h9 : {{1'd0}, _intrNO_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_2 = io_cfIn_intrVec_1 ? 4'h1 : _intrNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_3 = io_cfIn_intrVec_7 ? 4'h7 : _intrNO_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_4 = io_cfIn_intrVec_11 ? 4'hb : _intrNO_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _intrNO_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [5:0] _raiseIntr_T = {io_cfIn_intrVec_5,io_cfIn_intrVec_9,io_cfIn_intrVec_1,io_cfIn_intrVec_7,io_cfIn_intrVec_11,
    io_cfIn_intrVec_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:69]
  wire  raiseIntr = |_raiseIntr_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:76]
  wire  _illegalMret_T = io_in_valid & isMret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:33]
  wire  illegalMret = io_in_valid & isMret & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:43]
  wire  _illegalSret_T = io_in_valid & isSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 691:33]
  wire  illegalSret = io_in_valid & isSret & _intrVecEnable_0_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 691:43]
  wire  illegalSModeSret = _illegalSret_T & _tvm_T_1 & mstatusStruct_tsr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:76]
  wire  isIllegalPrivOp = illegalMret | illegalSret | illegalSModeSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 693:52]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:46]
  wire  csrExceptionVec_11 = _intrVecEnable_0_T_4 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 699:70]
  wire  csrExceptionVec_9 = _tvm_T_1 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 700:70]
  wire  csrExceptionVec_8 = _io_sfence_vma_invalid_T & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen | isIllegalPrivOp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:79]
  wire [7:0] raiseExceptionVec_lo = {hasStoreAccessFault,1'h0,hasLoadAccessFault,1'h0,csrExceptionVec_3,
    csrExceptionVec_2,hasInstrAccessFault,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:43]
  wire [15:0] _raiseExceptionVec_T = {hasStorePageFault,1'h0,hasLoadPageFault,1'h0,csrExceptionVec_11,1'h0,
    csrExceptionVec_9,csrExceptionVec_8,raiseExceptionVec_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:43]
  wire [15:0] raiseExceptionVec = _raiseExceptionVec_T | _wen_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:50]
  wire  raiseException = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 710:42]
  wire [2:0] _exceptionNO_T_1 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [2:0] _exceptionNO_T_3 = raiseExceptionVec[7] ? 3'h7 : _exceptionNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_5 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _exceptionNO_T_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_7 = raiseExceptionVec[15] ? 4'hf : _exceptionNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_9 = raiseExceptionVec[4] ? 4'h4 : _exceptionNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_11 = raiseExceptionVec[6] ? 4'h6 : _exceptionNO_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_13 = raiseExceptionVec[8] ? 4'h8 : _exceptionNO_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_15 = raiseExceptionVec[9] ? 4'h9 : _exceptionNO_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_17 = raiseExceptionVec[11] ? 4'hb : _exceptionNO_T_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_19 = raiseExceptionVec[0] ? 4'h0 : _exceptionNO_T_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_21 = raiseExceptionVec[2] ? 4'h2 : _exceptionNO_T_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_23 = raiseExceptionVec[1] ? 4'h1 : _exceptionNO_T_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_25 = raiseExceptionVec[12] ? 4'hc : _exceptionNO_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _exceptionNO_T_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:28]
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:53]
  wire [63:0] _GEN_145 = {{60'd0}, _causeNO_T_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:48]
  wire [63:0] causeNO = _causeNO_T | _GEN_145; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:48]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:58]
  wire [63:0] _redirectTarget_T_3 = _imemExceptionAddr_T_9 + 64'h4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:31]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 758:18]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 760:21]
  wire  delegS = _delegS_T_1[0] & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 760:36]
  wire [63:0] trapTarget = delegS ? stvec : mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 766:20]
  wire  _T_181 = io_in_valid & isUret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:15]
  wire  _T_179 = _illegalSret_T & ~illegalSret & ~illegalSModeSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:41]
  wire  _T_173 = _illegalMret_T & ~illegalMret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:25]
  wire [63:0] _GEN_109 = _illegalSret_T & ~illegalSret & ~illegalSModeSret ? sepc : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63 826:15]
  wire [63:0] retTarget = io_in_valid & isUret ? 64'h0 : _GEN_109; // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26 837:15]
  wire [63:0] _redirectTarget_T_4 = raiseExceptionIntr ? trapTarget : retTarget; // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:8]
  wire [63:0] redirectTarget = resetSatp ? _redirectTarget_T_3 : _redirectTarget_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 720:27]
  reg [63:0] redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
  wire  line_419_clock;
  wire  line_419_reset;
  wire  line_419_valid;
  reg  line_419_valid_reg;
  wire  addrNotLegal_signBit = redirectTargetReg[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,redirectTargetReg[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _addrNotLegal_T_3 = redirectTargetReg != _addrNotLegal_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 735:23]
  wire  _addrNotLegal_T_5 = |redirectTargetReg[63:39]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 736:44]
  wire  addrNotLegal = vmEnable ? _addrNotLegal_T_3 : _addrNotLegal_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 734:25]
  reg  hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
  reg  isIllegalXRET_REG; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
  wire  isIllegalXRET = isIllegalXRET_REG & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:50]
  wire  line_420_clock;
  wire  line_420_reset;
  wire  line_420_valid;
  reg  line_420_valid_reg;
  wire  line_421_clock;
  wire  line_421_reset;
  wire  line_421_valid;
  reg  line_421_valid_reg;
  wire  _T_162 = io_xretIsIllegal_ready & io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_422_clock;
  wire  line_422_reset;
  wire  line_422_valid;
  reg  line_422_valid_reg;
  wire  _GEN_84 = _T_162 ? 1'h0 : hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 742:38 743:20 738:31]
  wire  _GEN_85 = isIllegalXRET | _GEN_84; // @[src/main/scala/nutcore/backend/fu/CSR.scala 740:24 741:20]
  wire  isPageFault = hasInstrPageFault | hasLoadPageFault | hasStorePageFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 761:59]
  wire  isAddrMisAligned = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 762:48]
  wire  isAccessFault = hasInstrAccessFault | hasLoadAccessFault | hasStoreAccessFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 763:65]
  wire  line_423_clock;
  wire  line_423_reset;
  wire  line_423_valid;
  reg  line_423_valid_reg;
  wire  line_424_clock;
  wire  line_424_reset;
  wire  line_424_valid;
  reg  line_424_valid_reg;
  wire  line_425_clock;
  wire  line_425_reset;
  wire  line_425_valid;
  reg  line_425_valid_reg;
  wire  line_426_clock;
  wire  line_426_reset;
  wire  line_426_valid;
  reg  line_426_valid_reg;
  wire [63:0] _GEN_86 = delegS ? io_dmemExceptionAddr : _GEN_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 771:21 772:15]
  wire [63:0] _GEN_87 = delegS ? _GEN_79 : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 771:21 774:15]
  wire  line_427_clock;
  wire  line_427_reset;
  wire  line_427_valid;
  reg  line_427_valid_reg;
  wire  line_428_clock;
  wire  line_428_reset;
  wire  line_428_valid;
  reg  line_428_valid_reg;
  wire [63:0] tval = hasInstrPageFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 779:21]
  wire  line_429_clock;
  wire  line_429_reset;
  wire  line_429_valid;
  reg  line_429_valid_reg;
  wire  line_430_clock;
  wire  line_430_reset;
  wire  line_430_valid;
  reg  line_430_valid_reg;
  wire [63:0] _GEN_88 = delegS ? tval : _GEN_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 780:21 781:15]
  wire [63:0] _GEN_89 = delegS ? _GEN_79 : tval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 780:21 783:15]
  wire  line_431_clock;
  wire  line_431_reset;
  wire  line_431_valid;
  reg  line_431_valid_reg;
  wire  line_432_clock;
  wire  line_432_reset;
  wire  line_432_valid;
  reg  line_432_valid_reg;
  wire [63:0] tval_1 = hasInstrAccessFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 788:21]
  wire  line_433_clock;
  wire  line_433_reset;
  wire  line_433_valid;
  reg  line_433_valid_reg;
  wire  line_434_clock;
  wire  line_434_reset;
  wire  line_434_valid;
  reg  line_434_valid_reg;
  wire [63:0] _GEN_90 = delegS ? tval_1 : _GEN_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 789:21 790:15]
  wire [63:0] _GEN_91 = delegS ? _GEN_79 : tval_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 789:21 792:15]
  wire [63:0] _GEN_92 = isAccessFault ? _GEN_90 : _GEN_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:83]
  wire [63:0] _GEN_93 = isAccessFault ? _GEN_91 : _GEN_79; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:83]
  wire [63:0] _GEN_94 = isPageFault ? _GEN_88 : _GEN_92; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:77]
  wire [63:0] _GEN_95 = isPageFault ? _GEN_89 : _GEN_93; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:77]
  wire [63:0] _GEN_96 = isAddrMisAligned ? _GEN_86 : _GEN_94; // @[src/main/scala/nutcore/backend/fu/CSR.scala 770:60]
  wire [63:0] _GEN_97 = isAddrMisAligned ? _GEN_87 : _GEN_95; // @[src/main/scala/nutcore/backend/fu/CSR.scala 770:60]
  wire [63:0] _GEN_98 = io_instrValid ? _GEN_96 : _GEN_74; // @[src/main/scala/nutcore/backend/fu/CSR.scala 769:24]
  wire [63:0] _GEN_99 = io_instrValid ? _GEN_97 : _GEN_79; // @[src/main/scala/nutcore/backend/fu/CSR.scala 769:24]
  wire  line_435_clock;
  wire  line_435_reset;
  wire  line_435_valid;
  reg  line_435_valid_reg;
  wire  _T_174 = mstatusStruct_mpp != 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 803:26]
  wire  line_436_clock;
  wire  line_436_reset;
  wire  line_436_valid;
  reg  line_436_valid_reg;
  wire  mstatusNew_mprv = mstatusStruct_mpp != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 803:37 804:23 799:30]
  wire [5:0] mstatus_lo_lo = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [14:0] mstatus_lo = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,
    mstatus_lo_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [6:0] mstatus_hi_lo = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_mprv,
    mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [63:0] _mstatus_T_8 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [1:0] _GEN_101 = _illegalMret_T & ~illegalMret ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42 802:20 262:31]
  wire [63:0] _GEN_102 = _illegalMret_T & ~illegalMret ? _mstatus_T_8 : _GEN_65; // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42 808:13]
  wire  line_437_clock;
  wire  line_437_reset;
  wire  line_437_valid;
  reg  line_437_valid_reg;
  wire [1:0] _priviledgeMode_T = {1'h0,mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 818:26]
  wire [1:0] _GEN_146 = {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 819:26]
  wire  _T_180 = _GEN_146 != 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 819:26]
  wire  line_438_clock;
  wire  line_438_reset;
  wire  line_438_valid;
  reg  line_438_valid_reg;
  wire  mstatusNew_1_mprv = _GEN_146 != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 819:37 820:23 815:30]
  wire [5:0] mstatus_lo_lo_1 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [14:0] mstatus_lo_1 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [6:0] mstatus_hi_lo_1 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_1_mprv
    ,mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [63:0] _mstatus_T_9 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo_1,mstatus_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire  line_439_clock;
  wire  line_439_reset;
  wire  line_439_valid;
  reg  line_439_valid_reg;
  wire [5:0] mstatus_lo_lo_2 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [14:0] mstatus_lo_2 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m
    ,mstatusStruct_pie_h,mstatus_lo_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [6:0] mstatus_hi_lo_2 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,
    mstatusStruct_mprv,mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [63:0] _mstatus_T_10 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire  tvalZeroWen = ~(isPageFault | isAddrMisAligned | isAccessFault) | raiseIntr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 840:73]
  wire  line_440_clock;
  wire  line_440_reset;
  wire  line_440_valid;
  reg  line_440_valid_reg;
  wire  line_441_clock;
  wire  line_441_reset;
  wire  line_441_valid;
  reg  line_441_valid_reg;
  wire  line_442_clock;
  wire  line_442_reset;
  wire  line_442_valid;
  reg  line_442_valid_reg;
  wire  line_443_clock;
  wire  line_443_reset;
  wire  line_443_valid;
  reg  line_443_valid_reg;
  wire  line_444_clock;
  wire  line_444_reset;
  wire  line_444_valid;
  reg  line_444_valid_reg;
  wire [1:0] _GEN_117 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 848:22 843:30]
  wire  mstatusNew_3_pie_s = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 849:24 843:30]
  wire  mstatusNew_3_ie_s = delegS ? 1'h0 : mstatusStruct_ie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 850:23 843:30]
  wire [1:0] mstatusNew_3_mpp = delegS ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 860:22]
  wire  mstatusNew_3_pie_m = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 861:24]
  wire  mstatusNew_3_ie_m = delegS & mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 862:23]
  wire [5:0] mstatus_lo_lo_3 = {mstatusNew_3_pie_s,mstatusStruct_pie_u,mstatusNew_3_ie_m,mstatusStruct_ie_h,
    mstatusNew_3_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire  mstatusNew_3_spp = _GEN_117[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:30]
  wire [14:0] mstatus_lo_3 = {mstatusStruct_fs,mstatusNew_3_mpp,mstatusStruct_hpp,mstatusNew_3_spp,mstatusNew_3_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire [63:0] _mstatus_T_11 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire  perfCntCondDisable_0 = wen & _T_79 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1010:42]
  wire  _T_182 = ~perfCntCondDisable_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:92]
  wire  _WIRE = 1'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1001:{33,33}]
  wire  line_445_clock;
  wire  line_445_reset;
  wire  line_445_valid;
  reg  line_445_valid_reg;
  wire [63:0] _perfCnts_0_T_5 = perfCnts_0 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:105]
  wire  perfCntCondDisable_2 = wen & _T_81 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1010:42]
  wire  _T_187 = perfCntCondMinstret & ~perfCntCondDisable_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:89]
  wire  line_446_clock;
  wire  line_446_reset;
  wire  line_446_valid;
  reg  line_446_valid_reg;
  wire [63:0] _perfCnts_2_T_5 = perfCnts_2 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:105]
  wire  line_447_clock;
  wire  line_447_reset;
  wire  line_447_valid;
  reg  line_447_valid_reg;
  wire [63:0] _perfCnts_2_T_7 = perfCnts_2 + 64'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:86]
  wire  line_448_clock;
  wire  line_448_reset;
  wire  line_448_valid;
  reg  line_448_valid_reg;
  wire  line_449_clock;
  wire  line_449_reset;
  wire  line_449_valid;
  reg  line_449_valid_reg;
  wire [3:0] _T_198 = raiseIntr & io_instrValid ? intrNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1087:43]
  wire [3:0] _T_200 = raiseException & io_instrValid ? exceptionNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1088:43]
  CSRDiffWrapper CSRDiffWrapper ( // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
    .clock(CSRDiffWrapper_clock),
    .reset(CSRDiffWrapper_reset),
    .io_csrState_privilegeMode(CSRDiffWrapper_io_csrState_privilegeMode),
    .io_csrState_mstatus(CSRDiffWrapper_io_csrState_mstatus),
    .io_csrState_sstatus(CSRDiffWrapper_io_csrState_sstatus),
    .io_csrState_mepc(CSRDiffWrapper_io_csrState_mepc),
    .io_csrState_sepc(CSRDiffWrapper_io_csrState_sepc),
    .io_csrState_mtval(CSRDiffWrapper_io_csrState_mtval),
    .io_csrState_stval(CSRDiffWrapper_io_csrState_stval),
    .io_csrState_mtvec(CSRDiffWrapper_io_csrState_mtvec),
    .io_csrState_stvec(CSRDiffWrapper_io_csrState_stvec),
    .io_csrState_mcause(CSRDiffWrapper_io_csrState_mcause),
    .io_csrState_scause(CSRDiffWrapper_io_csrState_scause),
    .io_csrState_satp(CSRDiffWrapper_io_csrState_satp),
    .io_csrState_mip(CSRDiffWrapper_io_csrState_mip),
    .io_csrState_mie(CSRDiffWrapper_io_csrState_mie),
    .io_csrState_mscratch(CSRDiffWrapper_io_csrState_mscratch),
    .io_csrState_sscratch(CSRDiffWrapper_io_csrState_sscratch),
    .io_csrState_mideleg(CSRDiffWrapper_io_csrState_mideleg),
    .io_csrState_medeleg(CSRDiffWrapper_io_csrState_medeleg),
    .io_archEvent_valid(CSRDiffWrapper_io_archEvent_valid),
    .io_archEvent_interrupt(CSRDiffWrapper_io_archEvent_interrupt),
    .io_archEvent_exception(CSRDiffWrapper_io_archEvent_exception),
    .io_archEvent_exceptionPC(CSRDiffWrapper_io_archEvent_exceptionPC),
    .io_archEvent_exceptionInst(CSRDiffWrapper_io_archEvent_exceptionInst)
  );
  GEN_w1_line #(.COVER_INDEX(394)) line_394 (
    .clock(line_394_clock),
    .reset(line_394_reset),
    .valid(line_394_valid)
  );
  GEN_w1_line #(.COVER_INDEX(395)) line_395 (
    .clock(line_395_clock),
    .reset(line_395_reset),
    .valid(line_395_valid)
  );
  GEN_w1_line #(.COVER_INDEX(396)) line_396 (
    .clock(line_396_clock),
    .reset(line_396_reset),
    .valid(line_396_valid)
  );
  GEN_w1_line #(.COVER_INDEX(397)) line_397 (
    .clock(line_397_clock),
    .reset(line_397_reset),
    .valid(line_397_valid)
  );
  GEN_w1_line #(.COVER_INDEX(398)) line_398 (
    .clock(line_398_clock),
    .reset(line_398_reset),
    .valid(line_398_valid)
  );
  GEN_w1_line #(.COVER_INDEX(399)) line_399 (
    .clock(line_399_clock),
    .reset(line_399_reset),
    .valid(line_399_valid)
  );
  GEN_w1_line #(.COVER_INDEX(400)) line_400 (
    .clock(line_400_clock),
    .reset(line_400_reset),
    .valid(line_400_valid)
  );
  GEN_w1_line #(.COVER_INDEX(401)) line_401 (
    .clock(line_401_clock),
    .reset(line_401_reset),
    .valid(line_401_valid)
  );
  GEN_w1_line #(.COVER_INDEX(402)) line_402 (
    .clock(line_402_clock),
    .reset(line_402_reset),
    .valid(line_402_valid)
  );
  GEN_w1_line #(.COVER_INDEX(403)) line_403 (
    .clock(line_403_clock),
    .reset(line_403_reset),
    .valid(line_403_valid)
  );
  GEN_w1_line #(.COVER_INDEX(404)) line_404 (
    .clock(line_404_clock),
    .reset(line_404_reset),
    .valid(line_404_valid)
  );
  GEN_w1_line #(.COVER_INDEX(405)) line_405 (
    .clock(line_405_clock),
    .reset(line_405_reset),
    .valid(line_405_valid)
  );
  GEN_w1_line #(.COVER_INDEX(406)) line_406 (
    .clock(line_406_clock),
    .reset(line_406_reset),
    .valid(line_406_valid)
  );
  GEN_w1_line #(.COVER_INDEX(407)) line_407 (
    .clock(line_407_clock),
    .reset(line_407_reset),
    .valid(line_407_valid)
  );
  GEN_w1_line #(.COVER_INDEX(408)) line_408 (
    .clock(line_408_clock),
    .reset(line_408_reset),
    .valid(line_408_valid)
  );
  GEN_w1_line #(.COVER_INDEX(409)) line_409 (
    .clock(line_409_clock),
    .reset(line_409_reset),
    .valid(line_409_valid)
  );
  GEN_w1_line #(.COVER_INDEX(410)) line_410 (
    .clock(line_410_clock),
    .reset(line_410_reset),
    .valid(line_410_valid)
  );
  GEN_w1_line #(.COVER_INDEX(411)) line_411 (
    .clock(line_411_clock),
    .reset(line_411_reset),
    .valid(line_411_valid)
  );
  GEN_w1_line #(.COVER_INDEX(412)) line_412 (
    .clock(line_412_clock),
    .reset(line_412_reset),
    .valid(line_412_valid)
  );
  GEN_w1_line #(.COVER_INDEX(413)) line_413 (
    .clock(line_413_clock),
    .reset(line_413_reset),
    .valid(line_413_valid)
  );
  GEN_w1_line #(.COVER_INDEX(414)) line_414 (
    .clock(line_414_clock),
    .reset(line_414_reset),
    .valid(line_414_valid)
  );
  GEN_w1_line #(.COVER_INDEX(415)) line_415 (
    .clock(line_415_clock),
    .reset(line_415_reset),
    .valid(line_415_valid)
  );
  GEN_w1_line #(.COVER_INDEX(416)) line_416 (
    .clock(line_416_clock),
    .reset(line_416_reset),
    .valid(line_416_valid)
  );
  GEN_w1_line #(.COVER_INDEX(417)) line_417 (
    .clock(line_417_clock),
    .reset(line_417_reset),
    .valid(line_417_valid)
  );
  GEN_w1_line #(.COVER_INDEX(418)) line_418 (
    .clock(line_418_clock),
    .reset(line_418_reset),
    .valid(line_418_valid)
  );
  GEN_w1_line #(.COVER_INDEX(419)) line_419 (
    .clock(line_419_clock),
    .reset(line_419_reset),
    .valid(line_419_valid)
  );
  GEN_w1_line #(.COVER_INDEX(420)) line_420 (
    .clock(line_420_clock),
    .reset(line_420_reset),
    .valid(line_420_valid)
  );
  GEN_w1_line #(.COVER_INDEX(421)) line_421 (
    .clock(line_421_clock),
    .reset(line_421_reset),
    .valid(line_421_valid)
  );
  GEN_w1_line #(.COVER_INDEX(422)) line_422 (
    .clock(line_422_clock),
    .reset(line_422_reset),
    .valid(line_422_valid)
  );
  GEN_w1_line #(.COVER_INDEX(423)) line_423 (
    .clock(line_423_clock),
    .reset(line_423_reset),
    .valid(line_423_valid)
  );
  GEN_w1_line #(.COVER_INDEX(424)) line_424 (
    .clock(line_424_clock),
    .reset(line_424_reset),
    .valid(line_424_valid)
  );
  GEN_w1_line #(.COVER_INDEX(425)) line_425 (
    .clock(line_425_clock),
    .reset(line_425_reset),
    .valid(line_425_valid)
  );
  GEN_w1_line #(.COVER_INDEX(426)) line_426 (
    .clock(line_426_clock),
    .reset(line_426_reset),
    .valid(line_426_valid)
  );
  GEN_w1_line #(.COVER_INDEX(427)) line_427 (
    .clock(line_427_clock),
    .reset(line_427_reset),
    .valid(line_427_valid)
  );
  GEN_w1_line #(.COVER_INDEX(428)) line_428 (
    .clock(line_428_clock),
    .reset(line_428_reset),
    .valid(line_428_valid)
  );
  GEN_w1_line #(.COVER_INDEX(429)) line_429 (
    .clock(line_429_clock),
    .reset(line_429_reset),
    .valid(line_429_valid)
  );
  GEN_w1_line #(.COVER_INDEX(430)) line_430 (
    .clock(line_430_clock),
    .reset(line_430_reset),
    .valid(line_430_valid)
  );
  GEN_w1_line #(.COVER_INDEX(431)) line_431 (
    .clock(line_431_clock),
    .reset(line_431_reset),
    .valid(line_431_valid)
  );
  GEN_w1_line #(.COVER_INDEX(432)) line_432 (
    .clock(line_432_clock),
    .reset(line_432_reset),
    .valid(line_432_valid)
  );
  GEN_w1_line #(.COVER_INDEX(433)) line_433 (
    .clock(line_433_clock),
    .reset(line_433_reset),
    .valid(line_433_valid)
  );
  GEN_w1_line #(.COVER_INDEX(434)) line_434 (
    .clock(line_434_clock),
    .reset(line_434_reset),
    .valid(line_434_valid)
  );
  GEN_w1_line #(.COVER_INDEX(435)) line_435 (
    .clock(line_435_clock),
    .reset(line_435_reset),
    .valid(line_435_valid)
  );
  GEN_w1_line #(.COVER_INDEX(436)) line_436 (
    .clock(line_436_clock),
    .reset(line_436_reset),
    .valid(line_436_valid)
  );
  GEN_w1_line #(.COVER_INDEX(437)) line_437 (
    .clock(line_437_clock),
    .reset(line_437_reset),
    .valid(line_437_valid)
  );
  GEN_w1_line #(.COVER_INDEX(438)) line_438 (
    .clock(line_438_clock),
    .reset(line_438_reset),
    .valid(line_438_valid)
  );
  GEN_w1_line #(.COVER_INDEX(439)) line_439 (
    .clock(line_439_clock),
    .reset(line_439_reset),
    .valid(line_439_valid)
  );
  GEN_w1_line #(.COVER_INDEX(440)) line_440 (
    .clock(line_440_clock),
    .reset(line_440_reset),
    .valid(line_440_valid)
  );
  GEN_w1_line #(.COVER_INDEX(441)) line_441 (
    .clock(line_441_clock),
    .reset(line_441_reset),
    .valid(line_441_valid)
  );
  GEN_w1_line #(.COVER_INDEX(442)) line_442 (
    .clock(line_442_clock),
    .reset(line_442_reset),
    .valid(line_442_valid)
  );
  GEN_w1_line #(.COVER_INDEX(443)) line_443 (
    .clock(line_443_clock),
    .reset(line_443_reset),
    .valid(line_443_valid)
  );
  GEN_w1_line #(.COVER_INDEX(444)) line_444 (
    .clock(line_444_clock),
    .reset(line_444_reset),
    .valid(line_444_valid)
  );
  GEN_w1_line #(.COVER_INDEX(445)) line_445 (
    .clock(line_445_clock),
    .reset(line_445_reset),
    .valid(line_445_valid)
  );
  GEN_w1_line #(.COVER_INDEX(446)) line_446 (
    .clock(line_446_clock),
    .reset(line_446_reset),
    .valid(line_446_valid)
  );
  GEN_w1_line #(.COVER_INDEX(447)) line_447 (
    .clock(line_447_clock),
    .reset(line_447_reset),
    .valid(line_447_valid)
  );
  GEN_w1_line #(.COVER_INDEX(448)) line_448 (
    .clock(line_448_clock),
    .reset(line_448_reset),
    .valid(line_448_valid)
  );
  GEN_w1_line #(.COVER_INDEX(449)) line_449 (
    .clock(line_449_clock),
    .reset(line_449_reset),
    .valid(line_449_valid)
  );
  assign line_394_clock = clock;
  assign line_394_reset = reset;
  assign line_394_valid = set_lr ^ line_394_valid_reg;
  assign line_395_clock = clock;
  assign line_395_reset = reset;
  assign line_395_valid = _T_48 ^ line_395_valid_reg;
  assign line_396_clock = clock;
  assign line_396_reset = reset;
  assign line_396_valid = _T_50 ^ line_396_valid_reg;
  assign line_397_clock = clock;
  assign line_397_reset = reset;
  assign line_397_valid = _T_52 ^ line_397_valid_reg;
  assign line_398_clock = clock;
  assign line_398_reset = reset;
  assign line_398_valid = _T_54 ^ line_398_valid_reg;
  assign line_399_clock = clock;
  assign line_399_reset = reset;
  assign line_399_valid = _T_56 ^ line_399_valid_reg;
  assign line_400_clock = clock;
  assign line_400_reset = reset;
  assign line_400_valid = _T_58 ^ line_400_valid_reg;
  assign line_401_clock = clock;
  assign line_401_reset = reset;
  assign line_401_valid = _T_60 ^ line_401_valid_reg;
  assign line_402_clock = clock;
  assign line_402_reset = reset;
  assign line_402_valid = _T_62 ^ line_402_valid_reg;
  assign line_403_clock = clock;
  assign line_403_reset = reset;
  assign line_403_valid = _T_64 ^ line_403_valid_reg;
  assign line_404_clock = clock;
  assign line_404_reset = reset;
  assign line_404_valid = _T_66 ^ line_404_valid_reg;
  assign line_405_clock = clock;
  assign line_405_reset = reset;
  assign line_405_valid = _T_68 ^ line_405_valid_reg;
  assign line_406_clock = clock;
  assign line_406_reset = reset;
  assign line_406_valid = _T_70 ^ line_406_valid_reg;
  assign line_407_clock = clock;
  assign line_407_reset = reset;
  assign line_407_valid = _T_72 ^ line_407_valid_reg;
  assign line_408_clock = clock;
  assign line_408_reset = reset;
  assign line_408_valid = _T_74 ^ line_408_valid_reg;
  assign line_409_clock = clock;
  assign line_409_reset = reset;
  assign line_409_valid = _T_76 ^ line_409_valid_reg;
  assign line_410_clock = clock;
  assign line_410_reset = reset;
  assign line_410_valid = _T_78 ^ line_410_valid_reg;
  assign line_411_clock = clock;
  assign line_411_reset = reset;
  assign line_411_valid = _T_80 ^ line_411_valid_reg;
  assign line_412_clock = clock;
  assign line_412_reset = reset;
  assign line_412_valid = _T_82 ^ line_412_valid_reg;
  assign line_413_clock = clock;
  assign line_413_reset = reset;
  assign line_413_valid = _T_84 ^ line_413_valid_reg;
  assign line_414_clock = clock;
  assign line_414_reset = reset;
  assign line_414_valid = _T_86 ^ line_414_valid_reg;
  assign line_415_clock = clock;
  assign line_415_reset = reset;
  assign line_415_valid = _T_88 ^ line_415_valid_reg;
  assign line_416_clock = clock;
  assign line_416_reset = reset;
  assign line_416_valid = _T_90 ^ line_416_valid_reg;
  assign line_417_clock = clock;
  assign line_417_reset = reset;
  assign line_417_valid = _T_95 ^ line_417_valid_reg;
  assign line_418_clock = clock;
  assign line_418_reset = reset;
  assign line_418_valid = _T_97 ^ line_418_valid_reg;
  assign line_419_clock = clock;
  assign line_419_reset = reset;
  assign line_419_valid = io_redirect_valid ^ line_419_valid_reg;
  assign line_420_clock = clock;
  assign line_420_reset = reset;
  assign line_420_valid = isIllegalXRET ^ line_420_valid_reg;
  assign line_421_clock = clock;
  assign line_421_reset = reset;
  assign line_421_valid = isIllegalXRET ^ line_421_valid_reg;
  assign line_422_clock = clock;
  assign line_422_reset = reset;
  assign line_422_valid = _T_162 ^ line_422_valid_reg;
  assign line_423_clock = clock;
  assign line_423_reset = reset;
  assign line_423_valid = io_instrValid ^ line_423_valid_reg;
  assign line_424_clock = clock;
  assign line_424_reset = reset;
  assign line_424_valid = isAddrMisAligned ^ line_424_valid_reg;
  assign line_425_clock = clock;
  assign line_425_reset = reset;
  assign line_425_valid = delegS ^ line_425_valid_reg;
  assign line_426_clock = clock;
  assign line_426_reset = reset;
  assign line_426_valid = delegS ^ line_426_valid_reg;
  assign line_427_clock = clock;
  assign line_427_reset = reset;
  assign line_427_valid = isAddrMisAligned ^ line_427_valid_reg;
  assign line_428_clock = clock;
  assign line_428_reset = reset;
  assign line_428_valid = isPageFault ^ line_428_valid_reg;
  assign line_429_clock = clock;
  assign line_429_reset = reset;
  assign line_429_valid = delegS ^ line_429_valid_reg;
  assign line_430_clock = clock;
  assign line_430_reset = reset;
  assign line_430_valid = delegS ^ line_430_valid_reg;
  assign line_431_clock = clock;
  assign line_431_reset = reset;
  assign line_431_valid = isPageFault ^ line_431_valid_reg;
  assign line_432_clock = clock;
  assign line_432_reset = reset;
  assign line_432_valid = isAccessFault ^ line_432_valid_reg;
  assign line_433_clock = clock;
  assign line_433_reset = reset;
  assign line_433_valid = delegS ^ line_433_valid_reg;
  assign line_434_clock = clock;
  assign line_434_reset = reset;
  assign line_434_valid = delegS ^ line_434_valid_reg;
  assign line_435_clock = clock;
  assign line_435_reset = reset;
  assign line_435_valid = _T_173 ^ line_435_valid_reg;
  assign line_436_clock = clock;
  assign line_436_reset = reset;
  assign line_436_valid = _T_174 ^ line_436_valid_reg;
  assign line_437_clock = clock;
  assign line_437_reset = reset;
  assign line_437_valid = _T_179 ^ line_437_valid_reg;
  assign line_438_clock = clock;
  assign line_438_reset = reset;
  assign line_438_valid = _T_180 ^ line_438_valid_reg;
  assign line_439_clock = clock;
  assign line_439_reset = reset;
  assign line_439_valid = _T_181 ^ line_439_valid_reg;
  assign line_440_clock = clock;
  assign line_440_reset = reset;
  assign line_440_valid = raiseExceptionIntr ^ line_440_valid_reg;
  assign line_441_clock = clock;
  assign line_441_reset = reset;
  assign line_441_valid = delegS ^ line_441_valid_reg;
  assign line_442_clock = clock;
  assign line_442_reset = reset;
  assign line_442_valid = tvalZeroWen ^ line_442_valid_reg;
  assign line_443_clock = clock;
  assign line_443_reset = reset;
  assign line_443_valid = delegS ^ line_443_valid_reg;
  assign line_444_clock = clock;
  assign line_444_reset = reset;
  assign line_444_valid = tvalZeroWen ^ line_444_valid_reg;
  assign line_445_clock = clock;
  assign line_445_reset = reset;
  assign line_445_valid = _T_182 ^ line_445_valid_reg;
  assign line_446_clock = clock;
  assign line_446_reset = reset;
  assign line_446_valid = _T_187 ^ line_446_valid_reg;
  assign line_447_clock = clock;
  assign line_447_reset = reset;
  assign line_447_valid = perfCntCondMultiCommit ^ line_447_valid_reg;
  assign line_448_clock = clock;
  assign line_448_reset = reset;
  assign line_448_valid = perfCntCondDisable_0 ^ line_448_valid_reg;
  assign line_449_clock = clock;
  assign line_449_reset = reset;
  assign line_449_valid = perfCntCondDisable_2 ^ line_449_valid_reg;
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 880:16]
  assign io_out_bits = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_redirect_target = redirectTarget[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:22]
  assign io_redirect_valid = io_in_valid & _isEbreak_T_1 | raiseExceptionIntr | resetSatp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 727:80]
  assign io_xretIsIllegal_valid = hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 745:26]
  assign io_xretIsIllegal_bits = redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 746:25]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 603:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_wenFix = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 710:42]
  assign io_isPerfRead = io_out_valid & addr >= 12'hb00 & addr < 12'hb03; // @[src/main/scala/nutcore/backend/fu/CSR.scala 554:52]
  assign io_isExit = _io_isExit_T_10 & io_rfWenReal & rdata != 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:55]
  assign io_vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  assign io_sfence_vma_invalid = priviledgeMode == 2'h0 | tvm; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:53]
  assign io_wfi_invalid = priviledgeMode != 2'h3 & mstatusStruct_tw; // @[src/main/scala/nutcore/backend/fu/CSR.scala 546:46]
  assign lr_0 = lr;
  assign lrAddr_0 = lrAddr;
  assign satp_0 = satp;
  assign intrVecIDU_0 = intrVecIDU;
  assign CSRDiffWrapper_clock = clock;
  assign CSRDiffWrapper_reset = reset;
  assign CSRDiffWrapper_io_csrState_privilegeMode = {{62'd0}, priviledgeMode}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1066:28]
  assign CSRDiffWrapper_io_csrState_mstatus = mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1067:22]
  assign CSRDiffWrapper_io_csrState_sstatus = mstatus & 64'h80000003000d8122; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1068:33]
  assign CSRDiffWrapper_io_csrState_mepc = mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:19]
  assign CSRDiffWrapper_io_csrState_sepc = sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1070:19]
  assign CSRDiffWrapper_io_csrState_mtval = mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1071:19]
  assign CSRDiffWrapper_io_csrState_stval = stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1072:19]
  assign CSRDiffWrapper_io_csrState_mtvec = mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1073:20]
  assign CSRDiffWrapper_io_csrState_stvec = stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1074:20]
  assign CSRDiffWrapper_io_csrState_mcause = mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1075:21]
  assign CSRDiffWrapper_io_csrState_scause = scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1076:21]
  assign CSRDiffWrapper_io_csrState_satp = satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1077:19]
  assign CSRDiffWrapper_io_csrState_mip = mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1078:18]
  assign CSRDiffWrapper_io_csrState_mie = mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1079:18]
  assign CSRDiffWrapper_io_csrState_mscratch = mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1080:23]
  assign CSRDiffWrapper_io_csrState_sscratch = sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1081:23]
  assign CSRDiffWrapper_io_csrState_mideleg = mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1082:22]
  assign CSRDiffWrapper_io_csrState_medeleg = medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1083:22]
  assign CSRDiffWrapper_io_archEvent_valid = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:58]
  assign CSRDiffWrapper_io_archEvent_interrupt = {{28'd0}, _T_198}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1087:37]
  assign CSRDiffWrapper_io_archEvent_exception = {{28'd0}, _T_200}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1088:37]
  assign CSRDiffWrapper_io_archEvent_exceptionPC = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
  assign CSRDiffWrapper_io_archEvent_exceptionInst = io_cfIn_instr[31:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1090:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
      priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        priviledgeMode <= 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 851:22]
      end else begin
        priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 863:22]
      end
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
      priviledgeMode <= 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 834:20]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      priviledgeMode <= _priviledgeMode_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 818:20]
    end else begin
      priviledgeMode <= _GEN_101;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
      mtvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end else if (canWriteCSR & addr == 12'h305) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mtvec <= _mtvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
      mcounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end else if (canWriteCSR & addr == 12'h306) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mcounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
      mcause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mcause <= _GEN_71;
      end else begin
        mcause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 858:14]
      end
    end else begin
      mcause <= _GEN_71;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
      mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mtval <= _GEN_99;
      end else if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 864:26]
        mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 865:15]
      end else begin
        mtval <= _GEN_99;
      end
    end else begin
      mtval <= _GEN_99;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
      mepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mepc <= _GEN_78;
      end else if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
        mepc <= io_illegalJump_bits;
      end else begin
        mepc <= _imemExceptionAddr_T_11;
      end
    end else begin
      mepc <= _GEN_78;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
      mie <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end else if (canWriteCSR & addr == 12'h304) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (canWriteCSR & addr == 12'h104) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
      mipReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end else if (_canWriteCSR_T_1 & _io_isExit_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_canWriteCSR_T_1 & _io_isExit_T) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
      mstatus <= 64'ha00001800; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      mstatus <= _mstatus_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:13]
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
      mstatus <= _mstatus_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:13]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      mstatus <= _mstatus_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:13]
    end else begin
      mstatus <= _GEN_102;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
      medeleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end else if (canWriteCSR & addr == 12'h302) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      medeleg <= _medeleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
      mideleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end else if (canWriteCSR & addr == 12'h303) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mideleg <= _mideleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
      mscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end else if (canWriteCSR & addr == 12'h340) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
      stvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end else if (canWriteCSR & addr == 12'h105) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      stvec <= _stvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
      satp <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end else if (canWriteCSR & _isIllegalTVM_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      satp <= _satp_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
      sepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
          sepc <= io_illegalJump_bits;
        end else begin
          sepc <= _imemExceptionAddr_T_11;
        end
      end else begin
        sepc <= _GEN_70;
      end
    end else begin
      sepc <= _GEN_70;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
      scause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        scause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 846:14]
      end else begin
        scause <= _GEN_67;
      end
    end else begin
      scause <= _GEN_67;
    end
    if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:26]
          stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 853:15]
        end else begin
          stval <= _GEN_98;
        end
      end else begin
        stval <= _GEN_98;
      end
    end else begin
      stval <= _GEN_98;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
      sscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end else if (canWriteCSR & addr == 12'h140) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      sscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
      scounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end else if (canWriteCSR & addr == 12'h106) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      scounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 825:8]
    end else if (_illegalMret_T & ~illegalMret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 809:8]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lr <= set_lr_val; // @[src/main/scala/nutcore/backend/fu/CSR.scala 416:8]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
      lrAddr <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lrAddr <= set_lr_addr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 417:12]
    end
    line_394_valid_reg <= set_lr;
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (~perfCntCondDisable_0) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:96]
      perfCnts_0 <= _perfCnts_0_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:100]
    end else if (canWriteCSR & addr == 12'hb00) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (canWriteCSR & addr == 12'hb01) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:35]
      perfCnts_2 <= _perfCnts_2_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:60]
    end else if (perfCntCondMinstret & ~perfCntCondDisable_2) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:96]
      perfCnts_2 <= _perfCnts_2_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:100]
    end else if (canWriteCSR & addr == 12'hb02) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    line_395_valid_reg <= _T_48;
    line_396_valid_reg <= _T_50;
    line_397_valid_reg <= _T_52;
    line_398_valid_reg <= _T_54;
    line_399_valid_reg <= _T_56;
    line_400_valid_reg <= _T_58;
    line_401_valid_reg <= _T_60;
    line_402_valid_reg <= _T_62;
    line_403_valid_reg <= _T_64;
    line_404_valid_reg <= _T_66;
    line_405_valid_reg <= _T_68;
    line_406_valid_reg <= _T_70;
    line_407_valid_reg <= _T_72;
    line_408_valid_reg <= _T_74;
    line_409_valid_reg <= _T_76;
    line_410_valid_reg <= _T_78;
    line_411_valid_reg <= _T_80;
    line_412_valid_reg <= _T_82;
    line_413_valid_reg <= _T_84;
    line_414_valid_reg <= _T_86;
    line_415_valid_reg <= _T_88;
    line_416_valid_reg <= _T_90;
    line_417_valid_reg <= _T_95;
    line_418_valid_reg <= _T_97;
    if (io_redirect_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
      if (resetSatp) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 720:27]
        redirectTargetReg <= _redirectTarget_T_3;
      end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:8]
        if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 766:20]
          redirectTargetReg <= stvec;
        end else begin
          redirectTargetReg <= mtvec;
        end
      end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
        redirectTargetReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 837:15]
      end else begin
        redirectTargetReg <= _GEN_109;
      end
    end
    line_419_valid_reg <= io_redirect_valid;
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
      hasIllegalXRET <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
    end else begin
      hasIllegalXRET <= _GEN_85;
    end
    isIllegalXRET_REG <= io_redirect_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
    line_420_valid_reg <= isIllegalXRET;
    line_421_valid_reg <= isIllegalXRET;
    line_422_valid_reg <= _T_162;
    line_423_valid_reg <= io_instrValid;
    line_424_valid_reg <= isAddrMisAligned;
    line_425_valid_reg <= delegS;
    line_426_valid_reg <= delegS;
    line_427_valid_reg <= isAddrMisAligned;
    line_428_valid_reg <= isPageFault;
    line_429_valid_reg <= delegS;
    line_430_valid_reg <= delegS;
    line_431_valid_reg <= isPageFault;
    line_432_valid_reg <= isAccessFault;
    line_433_valid_reg <= delegS;
    line_434_valid_reg <= delegS;
    line_435_valid_reg <= _T_173;
    line_436_valid_reg <= _T_174;
    line_437_valid_reg <= _T_179;
    line_438_valid_reg <= _T_180;
    line_439_valid_reg <= _T_181;
    line_440_valid_reg <= raiseExceptionIntr;
    line_441_valid_reg <= delegS;
    line_442_valid_reg <= tvalZeroWen;
    line_443_valid_reg <= delegS;
    line_444_valid_reg <= tvalZeroWen;
    line_445_valid_reg <= _T_182;
    line_446_valid_reg <= _T_187;
    line_447_valid_reg <= perfCntCondMultiCommit;
    line_448_valid_reg <= perfCntCondDisable_0;
    line_449_valid_reg <= perfCntCondDisable_2;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priviledgeMode = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcounteren = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtval = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mepc = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mipReg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  stvec = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  satp = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  sepc = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  scause = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  stval = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  sscratch = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  scounteren = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  lr = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  lrAddr = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  line_394_valid_reg = _RAND_21[0:0];
  _RAND_22 = {2{`RANDOM}};
  perfCnts_0 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  perfCnts_1 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  perfCnts_2 = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  line_395_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_396_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_397_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_398_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_399_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_400_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_401_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_402_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_403_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_404_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_405_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_406_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_407_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_408_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_409_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_410_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_411_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_412_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_413_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_414_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_415_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_416_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_417_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_418_valid_reg = _RAND_48[0:0];
  _RAND_49 = {2{`RANDOM}};
  redirectTargetReg = _RAND_49[63:0];
  _RAND_50 = {1{`RANDOM}};
  line_419_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  hasIllegalXRET = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  isIllegalXRET_REG = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_420_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_421_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_422_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_423_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_424_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_425_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_426_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_427_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_428_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_429_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_430_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_431_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_432_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_433_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_434_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_435_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_436_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_437_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_438_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_439_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_440_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_441_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_442_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_443_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_444_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_445_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_446_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_447_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_448_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_449_valid_reg = _RAND_82[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (set_lr) begin
      cover(1'h1);
    end
    //
    if (_T_48) begin
      cover(1'h1);
    end
    //
    if (_T_50) begin
      cover(1'h1);
    end
    //
    if (_T_52) begin
      cover(1'h1);
    end
    //
    if (_T_54) begin
      cover(1'h1);
    end
    //
    if (_T_56) begin
      cover(1'h1);
    end
    //
    if (_T_58) begin
      cover(1'h1);
    end
    //
    if (_T_60) begin
      cover(1'h1);
    end
    //
    if (_T_62) begin
      cover(1'h1);
    end
    //
    if (_T_64) begin
      cover(1'h1);
    end
    //
    if (_T_66) begin
      cover(1'h1);
    end
    //
    if (_T_68) begin
      cover(1'h1);
    end
    //
    if (_T_70) begin
      cover(1'h1);
    end
    //
    if (_T_72) begin
      cover(1'h1);
    end
    //
    if (_T_74) begin
      cover(1'h1);
    end
    //
    if (_T_76) begin
      cover(1'h1);
    end
    //
    if (_T_78) begin
      cover(1'h1);
    end
    //
    if (_T_80) begin
      cover(1'h1);
    end
    //
    if (_T_82) begin
      cover(1'h1);
    end
    //
    if (_T_84) begin
      cover(1'h1);
    end
    //
    if (_T_86) begin
      cover(1'h1);
    end
    //
    if (_T_88) begin
      cover(1'h1);
    end
    //
    if (_T_90) begin
      cover(1'h1);
    end
    //
    if (_T_95) begin
      cover(1'h1);
    end
    //
    if (_T_97) begin
      cover(1'h1);
    end
    //
    if (io_redirect_valid) begin
      cover(1'h1);
    end
    //
    if (isIllegalXRET) begin
      cover(1'h1);
    end
    //
    if (~isIllegalXRET) begin
      cover(1'h1);
    end
    //
    if (~isIllegalXRET & _T_162) begin
      cover(1'h1);
    end
    //
    if (io_instrValid) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & isAddrMisAligned) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & isAddrMisAligned & delegS) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & isAddrMisAligned & ~delegS) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & isPageFault) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & isPageFault & delegS) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & isPageFault & ~delegS) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & ~isPageFault) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & ~isPageFault & isAccessFault) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & ~isPageFault & isAccessFault & delegS) begin
      cover(1'h1);
    end
    //
    if (io_instrValid & ~isAddrMisAligned & ~isPageFault & isAccessFault & ~delegS) begin
      cover(1'h1);
    end
    //
    if (_T_173) begin
      cover(1'h1);
    end
    //
    if (_T_173 & _T_174) begin
      cover(1'h1);
    end
    //
    if (_T_179) begin
      cover(1'h1);
    end
    //
    if (_T_179 & _T_180) begin
      cover(1'h1);
    end
    //
    if (_T_181) begin
      cover(1'h1);
    end
    //
    if (raiseExceptionIntr) begin
      cover(1'h1);
    end
    //
    if (raiseExceptionIntr & delegS) begin
      cover(1'h1);
    end
    //
    if (raiseExceptionIntr & delegS & tvalZeroWen) begin
      cover(1'h1);
    end
    //
    if (raiseExceptionIntr & ~delegS) begin
      cover(1'h1);
    end
    //
    if (raiseExceptionIntr & ~delegS & tvalZeroWen) begin
      cover(1'h1);
    end
    //
    if (_T_182) begin
      cover(1'h1);
    end
    //
    if (_T_187) begin
      cover(1'h1);
    end
    //
    if (perfCntCondMultiCommit) begin
      cover(1'h1);
    end
    //
    if (perfCntCondDisable_0) begin
      cover(1'h1);
    end
    //
    if (perfCntCondDisable_2) begin
      cover(1'h1);
    end
  end
endmodule
module MOU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DummyDPICWrapper_3(
  input         clock,
  input         reset,
  input         io_bits_hasTrap, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_cycleCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_instrCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_code, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasTrap; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_instrCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasWFI; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_code; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestTrapEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_hasTrap(dpic_io_hasTrap),
    .io_cycleCnt(dpic_io_cycleCnt),
    .io_instrCnt(dpic_io_instrCnt),
    .io_hasWFI(dpic_io_hasWFI),
    .io_code(dpic_io_code),
    .io_pc(dpic_io_pc),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_hasTrap = io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_cycleCnt = io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instrCnt = io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_hasWFI = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_code = io_bits_code; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module EXUDiffWrapper(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [38:0] io_in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [63:0] io_in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_code; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] cycleCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
  wire [63:0] _cycleCnt_T_1 = cycleCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:24]
  reg [63:0] instrCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
  wire [63:0] _instrCnt_T_1 = instrCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:26]
  wire  nutcoretrap = io_in_bits_ctrl_isNutCoreTrap & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 194:66]
  DummyDPICWrapper_3 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_hasTrap(difftest_module_io_bits_hasTrap),
    .io_bits_cycleCnt(difftest_module_io_bits_cycleCnt),
    .io_bits_instrCnt(difftest_module_io_bits_instrCnt),
    .io_bits_code(difftest_module_io_bits_code),
    .io_bits_pc(difftest_module_io_bits_pc)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_hasTrap = nutcoretrap; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 199:21]
  assign difftest_module_io_bits_cycleCnt = cycleCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 202:21]
  assign difftest_module_io_bits_instrCnt = instrCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 203:21]
  assign difftest_module_io_bits_code = io_in_bits_data_src1[31:0]; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 200:21]
  assign difftest_module_io_bits_pc = {{25'd0}, io_in_bits_cf_pc}; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 201:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
      cycleCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
    end else begin
      cycleCnt <= _cycleCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
      instrCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
    end else if (perfCntCondMinstret) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 189:22]
      instrCnt <= _instrCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cycleCnt = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  instrCnt = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [3:0]  io__in_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [2:0]  io__in_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [6:0]  io__in_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [4:0]  io__in_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__out_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__out_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isExit, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__forward_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__sfence_vma_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__wfi_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12_0,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         falseWire,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_1,
  input         io_extra_msip,
  input         io_in_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_offset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_iVmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_jumpIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isMissPredict; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_actualTarget; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_actualTaken; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_REG_0_fuOpType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [1:0] alu_REG_0_btbType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isRVC; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  lsu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [6:0] lsu_io__in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [31:0] lsu_io__instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbAF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scInflight_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_amoReq_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [55:0] lsu_dtlb_paddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_12_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scIsSuccess_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLrVal_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_DTLBFINISH; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lsuMMIO_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_13_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_setLrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  mdu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [6:0] mdu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  csr_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [6:0] csr_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_instrValid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_illegalJump_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wenFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isPerfRead; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_rfWenReal; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_meip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_lrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_satp_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_mtip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMultiCommit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr_val; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [11:0] csr_intrVecIDU_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_set_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_msip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  mou_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [6:0] mou_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushICache_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushTLB_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  diffMod_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [38:0] diffMod_io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [63:0] diffMod_io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  _fuValids_0_T_2 = ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:84]
  wire [15:0] _fuValids_0_T_4 = {2'h0,1'h0,io__in_bits_cf_exceptionVec_12,4'h0,4'h0,1'h0,io__in_bits_cf_exceptionVec_2,
    io__in_bits_cf_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:125]
  wire  _csr_io_cfIn_exceptionVec_13_T = lsu_io__in_valid & lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:62]
  wire  _csr_io_cfIn_exceptionVec_13_T_2 = io__in_bits_ctrl_fuOpType == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _csr_io_cfIn_exceptionVec_13_T_6 = io__in_bits_ctrl_fuOpType[5] & ~_csr_io_cfIn_exceptionVec_13_T_2 |
    io__in_bits_ctrl_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 64:69]
  wire  _csr_io_cfIn_exceptionVec_13_T_7 = ~_csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/fu/LSU.scala 65:40]
  wire  _T = alu_io_jumpIsIllegal_ready & alu_io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = csr_io_xretIsIllegal_ready & csr_io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_2 = _T | _T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:35]
  wire  line_450_clock;
  wire  line_450_reset;
  wire  line_450_valid;
  reg  line_450_valid_reg;
  wire  line_451_clock;
  wire  line_451_reset;
  wire  line_451_valid;
  reg  line_451_valid_reg;
  wire  line_452_clock;
  wire  line_452_reset;
  wire  line_452_valid;
  reg  line_452_valid_reg;
  wire  _GEN_4 = csr_io_vmEnable | io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 104:48 73:15]
  wire  _GEN_5 = csr_io_vmEnable ? io__in_bits_cf_exceptionVec_1 : 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 73:15 106:50]
  wire  fuValids_1 = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4
    ); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  fuValids_3 = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  _T_3 = io__out_bits_decode_ctrl_rfWen & csr_io_isPerfRead; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:39]
  wire  line_453_clock;
  wire  line_453_reset;
  wire  line_453_valid;
  reg  line_453_valid_reg;
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 53:12 src/main/scala/nutcore/backend/seq/EXU.scala 58:26]
  wire  _hasException_T_1 = lsuTlbPF | lsu_io__dtlbAF | lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 123:50]
  wire  _hasException_T_3 = _hasException_T_1 | lsu_io__storeAddrMisaligned | lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 124:63]
  wire  hasException = _hasException_T_3 | lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 125:30]
  wire [38:0] _io_out_bits_decode_cf_redirect_T_target = csr_io_redirect_valid ? csr_io_redirect_target :
    alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_bits_decode_cf_redirect_T_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_valid_T_1 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_3 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _io_out_valid_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_4 = _io_out_valid_T_3 | csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 146:6]
  wire  _io_forward_wb_rfData_T = alu_io_out_ready & alu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _T_10 = _io_forward_wb_rfData_T & ~isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 163:43]
  wire  _T_12 = _io_forward_wb_rfData_T & isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 164:43]
  wire  _T_13 = lsu_io__out_ready & lsu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_14 = mdu_io_out_ready & mdu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = csr_io_out_ready & csr_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  ALU alu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    .io_iVmEnable(alu_io_iVmEnable),
    .io_jumpIsIllegal_ready(alu_io_jumpIsIllegal_ready),
    .io_jumpIsIllegal_valid(alu_io_jumpIsIllegal_valid),
    .io_jumpIsIllegal_bits(alu_io_jumpIsIllegal_bits),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_actualTaken(alu_REG_0_actualTaken),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC)
  );
  UnpipelinedLSU lsu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsu_io__isMMIO),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__dtlbAF(lsu_io__dtlbAF),
    .io__vaddr(lsu_io__vaddr),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .io__loadAccessFault(lsu_io__loadAccessFault),
    .io__storeAccessFault(lsu_io__storeAccessFault),
    .setLr_0(lsu_setLr_0),
    .lr_0(lsu_lr_0),
    .scInflight_0(lsu_scInflight_0),
    .amoReq_0(lsu_amoReq_0),
    .lr_addr(lsu_lr_addr),
    .dtlb_paddr(lsu_dtlb_paddr),
    ._T_12_0(lsu__T_12_0),
    .scIsSuccess_0(lsu_scIsSuccess_0),
    .setLrVal_0(lsu_setLrVal_0),
    .vmEnable(lsu_vmEnable),
    .DTLBFINISH(lsu_DTLBFINISH),
    .lsuMMIO_0(lsu_lsuMMIO_0),
    ._T_13_1(lsu__T_13_1),
    .setLrAddr_0(lsu_setLrAddr_0)
  );
  MDU mdu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_5(csr_io_cfIn_exceptionVec_5),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_7(csr_io_cfIn_exceptionVec_7),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_exceptionVec_13(csr_io_cfIn_exceptionVec_13),
    .io_cfIn_exceptionVec_15(csr_io_cfIn_exceptionVec_15),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossBoundaryFault(csr_io_cfIn_crossBoundaryFault),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_illegalJump_valid(csr_io_illegalJump_valid),
    .io_illegalJump_bits(csr_io_illegalJump_bits),
    .io_dmemExceptionAddr(csr_io_dmemExceptionAddr),
    .io_xretIsIllegal_ready(csr_io_xretIsIllegal_ready),
    .io_xretIsIllegal_valid(csr_io_xretIsIllegal_valid),
    .io_xretIsIllegal_bits(csr_io_xretIsIllegal_bits),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_laf(csr_io_dmemMMU_laf),
    .io_dmemMMU_saf(csr_io_dmemMMU_saf),
    .io_wenFix(csr_io_wenFix),
    .io_isPerfRead(csr_io_isPerfRead),
    .io_isExit(csr_io_isExit),
    .io_vmEnable(csr_io_vmEnable),
    .io_rfWenReal(csr_io_rfWenReal),
    .io_sfence_vma_invalid(csr_io_sfence_vma_invalid),
    .io_wfi_invalid(csr_io_wfi_invalid),
    .set_lr(csr_set_lr),
    .lr_0(csr_lr_0),
    .meip_0(csr_meip_0),
    .lrAddr_0(csr_lrAddr_0),
    .satp_0(csr_satp_0),
    .mtip_0(csr_mtip_0),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .intrVecIDU_0(csr_intrVecIDU_0),
    .set_lr_addr(csr_set_lr_addr),
    .msip_0(csr_msip_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret)
  );
  MOU mou ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
    .clock(mou_clock),
    .reset(mou_reset),
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  EXUDiffWrapper diffMod ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
    .clock(diffMod_clock),
    .reset(diffMod_reset),
    .io_in_valid(diffMod_io_in_valid),
    .io_in_bits_cf_pc(diffMod_io_in_bits_cf_pc),
    .io_in_bits_ctrl_isNutCoreTrap(diffMod_io_in_bits_ctrl_isNutCoreTrap),
    .io_in_bits_data_src1(diffMod_io_in_bits_data_src1),
    .io_flush(diffMod_io_flush),
    .perfCntCondMinstret(diffMod_perfCntCondMinstret)
  );
  GEN_w1_line #(.COVER_INDEX(450)) line_450 (
    .clock(line_450_clock),
    .reset(line_450_reset),
    .valid(line_450_valid)
  );
  GEN_w1_line #(.COVER_INDEX(451)) line_451 (
    .clock(line_451_clock),
    .reset(line_451_reset),
    .valid(line_451_valid)
  );
  GEN_w1_line #(.COVER_INDEX(452)) line_452 (
    .clock(line_452_clock),
    .reset(line_452_reset),
    .valid(line_452_valid)
  );
  GEN_w1_line #(.COVER_INDEX(453)) line_453 (
    .clock(line_453_clock),
    .reset(line_453_reset),
    .valid(line_453_valid)
  );
  assign line_450_clock = clock;
  assign line_450_reset = reset;
  assign line_450_valid = _T_2 ^ line_450_valid_reg;
  assign line_451_clock = clock;
  assign line_451_reset = reset;
  assign line_451_valid = csr_io_vmEnable ^ line_451_valid_reg;
  assign line_452_clock = clock;
  assign line_452_reset = reset;
  assign line_452_valid = csr_io_vmEnable ^ line_452_valid_reg;
  assign line_453_clock = clock;
  assign line_453_reset = reset;
  assign line_453_valid = _T_3 ^ line_453_valid_reg;
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 154:31]
  assign io__out_valid = io__in_valid & _io_out_valid_T_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 143:31]
  assign io__out_bits_decode_cf_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 131:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 130:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target :
    _io_out_bits_decode_cf_redirect_T_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid :
    _io_out_bits_decode_cf_redirect_T_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 128:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~hasException | ~fuValids_1) & ~(csr_io_wenFix &
    fuValids_3); // @[src/main/scala/nutcore/backend/seq/EXU.scala 126:68]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 127:14]
  assign io__out_bits_isMMIO = io__out_bits_decode_ctrl_rfWen & csr_io_isPerfRead | lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:61 112:24 62:22]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 148:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 149:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 151:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 150:35]
  assign io__out_bits_isExit = csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 134:22]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__forward_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 156:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/EXU.scala 157:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 158:24]
  assign io__forward_wb_rfData = _io_forward_wb_rfData_T ? alu_io_out_bits : lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 159:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 160:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 89:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__sfence_vma_invalid = csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 86:25]
  assign io__wfi_invalid = csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 87:18]
  assign lr = csr_lr_0;
  assign scInflight = lsu_scInflight_0;
  assign REG_valid = alu_REG_0_valid;
  assign REG_pc = alu_REG_0_pc;
  assign REG_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_actualTarget = alu_REG_0_actualTarget;
  assign REG_actualTaken = alu_REG_0_actualTaken;
  assign REG_fuOpType = alu_REG_0_fuOpType;
  assign REG_btbType = alu_REG_0_btbType;
  assign REG_isRVC = alu_REG_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign lrAddr = csr_lrAddr_0;
  assign satp = csr_satp_0;
  assign flushICache = mou_flushICache_0;
  assign flushTLB = mou_flushTLB_0;
  assign intrVecIDU = csr_intrVecIDU_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 85:15]
  assign alu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 53:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/EXU.scala 52:17]
  assign alu_io_iVmEnable = csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 90:20]
  assign alu_io_jumpIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:45]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 51:21]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 52:21]
  assign lsu_io__out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 64:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/EXU.scala 61:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_lr_0 = lr;
  assign lsu_lr_addr = lrAddr;
  assign lsu_dtlb_paddr = paddr;
  assign lsu__T_12_0 = _T_12_0;
  assign lsu_scIsSuccess_0 = scIsSuccess;
  assign lsu_vmEnable = vmEnable;
  assign lsu_DTLBFINISH = tlbFinish;
  assign lsu_lsuMMIO_0 = ismmio;
  assign lsu__T_13_1 = _T_13_1;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4)
    ; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/CSR.scala 207:15]
  assign csr_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 84:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_1 = _T | _T_1 ? _GEN_5 : io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 74:48]
  assign csr_io_cfIn_exceptionVec_5 = lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 76:45]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:49]
  assign csr_io_cfIn_exceptionVec_7 = lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 77:46]
  assign csr_io_cfIn_exceptionVec_12 = _T | _T_1 ? _GEN_4 : io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_13 = lsu_io__in_valid & lsu_io__dtlbPF & _csr_io_cfIn_exceptionVec_13_T_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:79]
  assign csr_io_cfIn_exceptionVec_15 = _csr_io_cfIn_exceptionVec_13_T & _csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 79:80]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_crossBoundaryFault = io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_instrValid = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:36]
  assign csr_io_illegalJump_valid = alu_io_jumpIsIllegal_valid | csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 95:60]
  assign csr_io_illegalJump_bits = alu_io_jumpIsIllegal_valid ? alu_io_jumpIsIllegal_bits : csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 96:36]
  assign csr_io_dmemExceptionAddr = lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:28]
  assign csr_io_xretIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 98:45]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_laf = io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_saf = io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_rfWenReal = io__in_bits_ctrl_rfWen & io__in_bits_ctrl_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 85:45]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_msip_0 = io_extra_msip;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign mou_clock = clock;
  assign mou_reset = reset;
  assign mou_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 118:15]
  assign diffMod_clock = clock;
  assign diffMod_reset = reset;
  assign diffMod_io_in_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 171:25]
  assign diffMod_io_in_bits_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_ctrl_isNutCoreTrap = io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_data_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_flush = io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 173:22]
  assign diffMod_perfCntCondMinstret = io_in_valid;
  always @(posedge clock) begin
    line_450_valid_reg <= _T_2;
    line_451_valid_reg <= csr_io_vmEnable;
    line_452_valid_reg <= csr_io_vmEnable;
    line_453_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_450_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_451_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_452_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_453_valid_reg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & csr_io_vmEnable) begin
      cover(1'h1);
    end
    //
    if (_T_2 & ~csr_io_vmEnable) begin
      cover(1'h1);
    end
    //
    if (_T_3) begin
      cover(1'h1);
    end
  end
endmodule
module DummyDPICWrapper_4(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_skip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_isRVC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_rfwen, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_wpdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_wdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_instr, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_special // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_skip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isRVC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_rfwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_fpwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_vecwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_wpdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_wdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_instr; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [9:0] dpic_io_robIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_lqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_sqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isLoad; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isStore; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_nFused; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_special; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestInstrCommit dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_skip(dpic_io_skip),
    .io_isRVC(dpic_io_isRVC),
    .io_rfwen(dpic_io_rfwen),
    .io_fpwen(dpic_io_fpwen),
    .io_vecwen(dpic_io_vecwen),
    .io_wpdest(dpic_io_wpdest),
    .io_wdest(dpic_io_wdest),
    .io_pc(dpic_io_pc),
    .io_instr(dpic_io_instr),
    .io_robIdx(dpic_io_robIdx),
    .io_lqIdx(dpic_io_lqIdx),
    .io_sqIdx(dpic_io_sqIdx),
    .io_isLoad(dpic_io_isLoad),
    .io_isStore(dpic_io_isStore),
    .io_nFused(dpic_io_nFused),
    .io_special(dpic_io_special),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_skip = io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isRVC = io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_rfwen = io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_fpwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_vecwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wpdest = io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wdest = io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instr = io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_robIdx = 10'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_lqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isLoad = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isStore = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_nFused = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_special = io_bits_special; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DiffInstrCommitWrapper(
  input         clock,
  input         reset,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input         io_skip, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input         io_isRVC, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input         io_rfwen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input  [4:0]  io_wpdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input  [7:0]  io_wdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input  [63:0] io_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input  [31:0] io_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
  input  [7:0]  io_special // @[src/main/scala/nutcore/backend/seq/WBU.scala 64:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_special; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg  difftest_REG_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg  difftest_REG_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg  difftest_REG_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg [4:0] difftest_REG_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg [7:0] difftest_REG_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg [63:0] difftest_REG_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg [31:0] difftest_REG_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  reg [7:0] difftest_REG_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  DummyDPICWrapper_4 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_skip(difftest_module_io_bits_skip),
    .io_bits_isRVC(difftest_module_io_bits_isRVC),
    .io_bits_rfwen(difftest_module_io_bits_rfwen),
    .io_bits_wpdest(difftest_module_io_bits_wpdest),
    .io_bits_wdest(difftest_module_io_bits_wdest),
    .io_bits_pc(difftest_module_io_bits_pc),
    .io_bits_instr(difftest_module_io_bits_instr),
    .io_bits_special(difftest_module_io_bits_special)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_skip = difftest_REG_skip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_isRVC = difftest_REG_isRVC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_rfwen = difftest_REG_rfwen; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_wpdest = difftest_REG_wpdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_wdest = difftest_REG_wdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_pc = difftest_REG_pc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_instr = difftest_REG_instr; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  assign difftest_module_io_bits_special = difftest_REG_special; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 67:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_skip <= io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_isRVC <= io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_rfwen <= io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_wpdest <= io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_wdest <= io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_pc <= io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_instr <= io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
    difftest_REG_special <= io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 67:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_skip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  difftest_REG_isRVC = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  difftest_REG_rfwen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  difftest_REG_wpdest = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  difftest_REG_wdest = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_pc = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  difftest_REG_instr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  difftest_REG_special = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_5(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_address, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_address; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestIntWriteback dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_address(dpic_io_address),
    .io_data(dpic_io_data),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_address = io_bits_address; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DiffIntWbWrapper(
  input         clock,
  input         reset,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 100:18]
  input  [4:0]  io_address, // @[src/main/scala/nutcore/backend/seq/WBU.scala 100:18]
  input  [63:0] io_data // @[src/main/scala/nutcore/backend/seq/WBU.scala 100:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_address; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
  reg [4:0] difftest_REG_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
  reg [63:0] difftest_REG_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
  DummyDPICWrapper_5 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_address(difftest_module_io_bits_address),
    .io_bits_data(difftest_module_io_bits_data)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 102:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 102:16]
  assign difftest_module_io_bits_address = difftest_REG_address; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 102:16]
  assign difftest_module_io_bits_data = difftest_REG_data; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 102:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
    difftest_REG_address <= io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
    difftest_REG_data <= io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 102:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_address = _RAND_1[4:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_data = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [2:0]  io__in_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isExit, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__wb_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [4:0]  io__wb_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [63:0] io__wb_rfData, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [38:0] io__redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        falseWire_0,
  output        io_in_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  DiffInstrCommitWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffInstrCommitWrapper_reset; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffInstrCommitWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffInstrCommitWrapper_io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffInstrCommitWrapper_io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffInstrCommitWrapper_io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire [4:0] DiffInstrCommitWrapper_io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire [7:0] DiffInstrCommitWrapper_io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire [63:0] DiffInstrCommitWrapper_io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire [31:0] DiffInstrCommitWrapper_io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire [7:0] DiffInstrCommitWrapper_io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
  wire  DiffIntWbWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
  wire  DiffIntWbWrapper_reset; // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
  wire  DiffIntWbWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
  wire [4:0] DiffIntWbWrapper_io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
  wire [63:0] DiffIntWbWrapper_io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
  wire  line_454_clock;
  wire  line_454_reset;
  wire  line_454_valid;
  reg  line_454_valid_reg;
  wire  line_455_clock;
  wire  line_455_reset;
  wire  line_455_valid;
  reg  line_455_valid_reg;
  wire [63:0] _GEN_6 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  line_456_clock;
  wire  line_456_reset;
  wire  line_456_valid;
  reg  line_456_valid_reg;
  wire [63:0] _GEN_7 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_6; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  line_457_clock;
  wire  line_457_reset;
  wire  line_457_valid;
  reg  line_457_valid_reg;
  wire [63:0] _GEN_8 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_7; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  line_458_clock;
  wire  line_458_reset;
  wire  line_458_valid;
  reg  line_458_valid_reg;
  wire  signBit = io__in_bits_decode_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _T = signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire  _T_4 = io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 85:51]
  wire [1:0] _T_6 = {io__in_bits_isExit,1'h0}; // @[difftest/src/main/scala/Bundles.scala 81:19]
  wire  falseWire = 1'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 58:{27,27}]
  DiffInstrCommitWrapper DiffInstrCommitWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 78:26]
    .clock(DiffInstrCommitWrapper_clock),
    .reset(DiffInstrCommitWrapper_reset),
    .io_valid(DiffInstrCommitWrapper_io_valid),
    .io_skip(DiffInstrCommitWrapper_io_skip),
    .io_isRVC(DiffInstrCommitWrapper_io_isRVC),
    .io_rfwen(DiffInstrCommitWrapper_io_rfwen),
    .io_wpdest(DiffInstrCommitWrapper_io_wpdest),
    .io_wdest(DiffInstrCommitWrapper_io_wdest),
    .io_pc(DiffInstrCommitWrapper_io_pc),
    .io_instr(DiffInstrCommitWrapper_io_instr),
    .io_special(DiffInstrCommitWrapper_io_special)
  );
  DiffIntWbWrapper DiffIntWbWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 110:26]
    .clock(DiffIntWbWrapper_clock),
    .reset(DiffIntWbWrapper_reset),
    .io_valid(DiffIntWbWrapper_io_valid),
    .io_address(DiffIntWbWrapper_io_address),
    .io_data(DiffIntWbWrapper_io_data)
  );
  GEN_w1_line #(.COVER_INDEX(454)) line_454 (
    .clock(line_454_clock),
    .reset(line_454_reset),
    .valid(line_454_valid)
  );
  GEN_w1_line #(.COVER_INDEX(455)) line_455 (
    .clock(line_455_clock),
    .reset(line_455_reset),
    .valid(line_455_valid)
  );
  GEN_w1_line #(.COVER_INDEX(456)) line_456 (
    .clock(line_456_clock),
    .reset(line_456_reset),
    .valid(line_456_valid)
  );
  GEN_w1_line #(.COVER_INDEX(457)) line_457 (
    .clock(line_457_clock),
    .reset(line_457_reset),
    .valid(line_457_valid)
  );
  GEN_w1_line #(.COVER_INDEX(458)) line_458 (
    .clock(line_458_clock),
    .reset(line_458_reset),
    .valid(line_458_valid)
  );
  assign line_454_clock = clock;
  assign line_454_reset = reset;
  assign line_454_valid = 3'h0 == io__in_bits_decode_ctrl_fuType ^ line_454_valid_reg;
  assign line_455_clock = clock;
  assign line_455_reset = reset;
  assign line_455_valid = 3'h1 == io__in_bits_decode_ctrl_fuType ^ line_455_valid_reg;
  assign line_456_clock = clock;
  assign line_456_reset = reset;
  assign line_456_valid = 3'h2 == io__in_bits_decode_ctrl_fuType ^ line_456_valid_reg;
  assign line_457_clock = clock;
  assign line_457_reset = reset;
  assign line_457_valid = 3'h3 == io__in_bits_decode_ctrl_fuType ^ line_457_valid_reg;
  assign line_458_clock = clock;
  assign line_458_reset = reset;
  assign line_458_valid = 3'h4 == io__in_bits_decode_ctrl_fuType ^ line_458_valid_reg;
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 35:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 36:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_8; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/seq/WBU.scala 41:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 42:60]
  assign falseWire_0 = falseWire;
  assign io_in_valid = io__in_valid;
  assign DiffInstrCommitWrapper_clock = clock;
  assign DiffInstrCommitWrapper_reset = reset;
  assign DiffInstrCommitWrapper_io_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 80:20]
  assign DiffInstrCommitWrapper_io_skip = io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/seq/WBU.scala 83:19]
  assign DiffInstrCommitWrapper_io_isRVC = io__in_bits_decode_cf_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 84:56]
  assign DiffInstrCommitWrapper_io_rfwen = io__wb_rfWen & io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 85:35]
  assign DiffInstrCommitWrapper_io_wpdest = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 87:21]
  assign DiffInstrCommitWrapper_io_wdest = {{3'd0}, io__wb_rfDest}; // @[src/main/scala/nutcore/backend/seq/WBU.scala 86:20]
  assign DiffInstrCommitWrapper_io_pc = {_T,io__in_bits_decode_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  assign DiffInstrCommitWrapper_io_instr = io__in_bits_decode_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:20]
  assign DiffInstrCommitWrapper_io_special = {{6'd0}, _T_6}; // @[difftest/src/main/scala/Bundles.scala 81:13]
  assign DiffIntWbWrapper_clock = clock;
  assign DiffIntWbWrapper_reset = reset;
  assign DiffIntWbWrapper_io_valid = io__wb_rfWen & _T_4; // @[src/main/scala/nutcore/backend/seq/WBU.scala 112:35]
  assign DiffIntWbWrapper_io_address = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 113:22]
  assign DiffIntWbWrapper_io_data = io__wb_rfData; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:19]
  always @(posedge clock) begin
    line_454_valid_reg <= 3'h0 == io__in_bits_decode_ctrl_fuType;
    line_455_valid_reg <= 3'h1 == io__in_bits_decode_ctrl_fuType;
    line_456_valid_reg <= 3'h2 == io__in_bits_decode_ctrl_fuType;
    line_457_valid_reg <= 3'h3 == io__in_bits_decode_ctrl_fuType;
    line_458_valid_reg <= 3'h4 == io__in_bits_decode_ctrl_fuType;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_454_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_455_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_456_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_457_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_458_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (3'h0 == io__in_bits_decode_ctrl_fuType) begin
      cover(1'h1);
    end
    //
    if (3'h1 == io__in_bits_decode_ctrl_fuType) begin
      cover(1'h1);
    end
    //
    if (3'h2 == io__in_bits_decode_ctrl_fuType) begin
      cover(1'h1);
    end
    //
    if (3'h3 == io__in_bits_decode_ctrl_fuType) begin
      cover(1'h1);
    end
    //
    if (3'h4 == io__in_bits_decode_ctrl_fuType) begin
      cover(1'h1);
    end
  end
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output        REG_actualTaken,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_0,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_lr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_meip_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scInflight; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isMissPredict; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_actualTarget; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_actualTaken; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_REG_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_REG_btbType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isRVC; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_amoReq; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_lrAddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [55:0] exu_paddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_satp; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_12_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scIsSuccess; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_mtip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushICache; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_falseWire; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_vmEnable; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushTLB; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [11:0] exu_intrVecIDU; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_tlbFinish; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_ismmio; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_13_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_msip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_falseWire_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  line_459_clock;
  wire  line_459_reset;
  wire  line_459_valid;
  reg  line_459_valid_reg;
  wire  _GEN_8 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  line_460_clock;
  wire  line_460_reset;
  wire  line_460_valid;
  reg  line_460_valid_reg;
  wire  _GEN_9 = isu_io_out_valid & exu_io__in_ready | _GEN_8; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  wire  line_461_clock;
  wire  line_461_reset;
  wire  line_461_valid;
  reg  line_461_valid_reg;
  reg [63:0] exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  line_462_clock;
  wire  line_462_reset;
  wire  line_462_valid;
  reg  line_462_valid_reg;
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _T_4 = exu_io__out_valid; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  line_463_clock;
  wire  line_463_reset;
  wire  line_463_valid;
  reg  line_463_valid_reg;
  wire  line_464_clock;
  wire  line_464_reset;
  wire  line_464_valid;
  reg  line_464_valid_reg;
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  line_465_clock;
  wire  line_465_reset;
  wire  line_465_valid;
  reg  line_465_valid_reg;
  ISU isu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(isu_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(isu_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(isu_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(isu_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossBoundaryFault(exu_io__in_bits_cf_crossBoundaryFault),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_isNutCoreTrap(exu_io__in_bits_ctrl_isNutCoreTrap),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_instr(exu_io__out_bits_decode_cf_instr),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_isMMIO(exu_io__out_bits_isMMIO),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__out_bits_isExit(exu_io__out_bits_isExit),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_laf(exu_io__memMMU_dmem_laf),
    .io__memMMU_dmem_saf(exu_io__memMMU_dmem_saf),
    .io__sfence_vma_invalid(exu_io__sfence_vma_invalid),
    .io__wfi_invalid(exu_io__wfi_invalid),
    .lr(exu_lr),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .scInflight(exu_scInflight),
    .REG_valid(exu_REG_valid),
    .REG_pc(exu_REG_pc),
    .REG_isMissPredict(exu_REG_isMissPredict),
    .REG_actualTarget(exu_REG_actualTarget),
    .REG_actualTaken(exu_REG_actualTaken),
    .REG_fuOpType(exu_REG_fuOpType),
    .REG_btbType(exu_REG_btbType),
    .REG_isRVC(exu_REG_isRVC),
    .amoReq(exu_amoReq),
    .lrAddr(exu_lrAddr),
    .paddr(exu_paddr),
    .satp(exu_satp),
    ._T_12_0(exu__T_12_0),
    .scIsSuccess(exu_scIsSuccess),
    .io_extra_mtip(exu_io_extra_mtip),
    .flushICache(exu_flushICache),
    .falseWire(exu_falseWire),
    .vmEnable(exu_vmEnable),
    .flushTLB(exu_flushTLB),
    .intrVecIDU(exu_intrVecIDU),
    .tlbFinish(exu_tlbFinish),
    .ismmio(exu_ismmio),
    ._T_13_1(exu__T_13_1),
    .io_extra_msip(exu_io_extra_msip),
    .io_in_valid(exu_io_in_valid)
  );
  WBU wbu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_isMMIO(wbu_io__in_bits_isMMIO),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_isExit(wbu_io__in_bits_isExit),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .falseWire_0(wbu_falseWire_0),
    .io_in_valid(wbu_io_in_valid)
  );
  GEN_w1_line #(.COVER_INDEX(459)) line_459 (
    .clock(line_459_clock),
    .reset(line_459_reset),
    .valid(line_459_valid)
  );
  GEN_w1_line #(.COVER_INDEX(460)) line_460 (
    .clock(line_460_clock),
    .reset(line_460_reset),
    .valid(line_460_valid)
  );
  GEN_w1_line #(.COVER_INDEX(461)) line_461 (
    .clock(line_461_clock),
    .reset(line_461_reset),
    .valid(line_461_valid)
  );
  GEN_w1_line #(.COVER_INDEX(462)) line_462 (
    .clock(line_462_clock),
    .reset(line_462_reset),
    .valid(line_462_valid)
  );
  GEN_w1_line #(.COVER_INDEX(463)) line_463 (
    .clock(line_463_clock),
    .reset(line_463_reset),
    .valid(line_463_valid)
  );
  GEN_w1_line #(.COVER_INDEX(464)) line_464 (
    .clock(line_464_clock),
    .reset(line_464_reset),
    .valid(line_464_valid)
  );
  GEN_w1_line #(.COVER_INDEX(465)) line_465 (
    .clock(line_465_clock),
    .reset(line_465_reset),
    .valid(line_465_valid)
  );
  assign line_459_clock = clock;
  assign line_459_reset = reset;
  assign line_459_valid = _T ^ line_459_valid_reg;
  assign line_460_clock = clock;
  assign line_460_reset = reset;
  assign line_460_valid = _T_2 ^ line_460_valid_reg;
  assign line_461_clock = clock;
  assign line_461_reset = reset;
  assign line_461_valid = io_flush[0] ^ line_461_valid_reg;
  assign line_462_clock = clock;
  assign line_462_reset = reset;
  assign line_462_valid = _T_2 ^ line_462_valid_reg;
  assign line_463_clock = clock;
  assign line_463_reset = reset;
  assign line_463_valid = _T_4 ^ line_463_valid_reg;
  assign line_464_clock = clock;
  assign line_464_reset = reset;
  assign line_464_valid = io_flush[1] ^ line_464_valid_reg;
  assign line_465_clock = clock;
  assign line_465_reset = reset;
  assign line_465_valid = _T_4 ^ line_465_valid_reg;
  assign io_in_0_ready = isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 698:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_sfence_vma_invalid = exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:25]
  assign io_wfi_invalid = exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign lr = exu_lr;
  assign scInflight = exu_scInflight;
  assign REG_valid = exu_REG_valid;
  assign REG_pc = exu_REG_pc;
  assign REG_isMissPredict = exu_REG_isMissPredict;
  assign REG_actualTarget = exu_REG_actualTarget;
  assign REG_actualTaken = exu_REG_actualTaken;
  assign REG_fuOpType = exu_REG_fuOpType;
  assign REG_btbType = exu_REG_btbType;
  assign REG_isRVC = exu_REG_isRVC;
  assign amoReq = exu_amoReq;
  assign lrAddr = exu_lrAddr;
  assign satp = exu_satp;
  assign flushICache = exu_flushICache;
  assign flushTLB = exu_flushTLB;
  assign intrVecIDU = exu_intrVecIDU;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_flush = io_flush[0]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 688:27]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossBoundaryFault = exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_isNutCoreTrap = exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 689:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_laf = io_memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_saf = io_memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_paddr = paddr;
  assign exu__T_12_0 = _T_12;
  assign exu_scIsSuccess = scIsSuccess;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_falseWire = wbu_falseWire_0;
  assign exu_vmEnable = vmEnable;
  assign exu_tlbFinish = tlbFinish;
  assign exu_ismmio = ismmio;
  assign exu__T_13_1 = _T_13_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isMMIO = wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isExit = wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_9;
    end
    line_459_valid_reg <= _T;
    line_460_valid_reg <= _T_2;
    line_461_valid_reg <= io_flush[0];
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_instr <= isu_io_out_bits_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pc <= isu_io_out_bits_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_crossBoundaryFault <= isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_isNutCoreTrap <= isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src1 <= isu_io_out_bits_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src2 <= isu_io_out_bits_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_imm <= isu_io_out_bits_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    line_462_valid_reg <= _T_2;
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _T_4;
    end
    line_463_valid_reg <= _T_4;
    line_464_valid_reg <= io_flush[1];
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_instr <= exu_io__out_bits_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isMMIO <= exu_io__out_bits_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_0 <= exu_io__out_bits_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_1 <= exu_io__out_bits_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_2 <= exu_io__out_bits_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_3 <= exu_io__out_bits_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isExit <= exu_io__out_bits_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    line_465_valid_reg <= _T_4;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_459_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_460_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_461_valid_reg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc = _RAND_5[38:0];
  _RAND_6 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_12 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_crossBoundaryFault = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_isNutCoreTrap = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm = _RAND_25[63:0];
  _RAND_26 = {1{`RANDOM}};
  line_462_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_463_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_464_valid_reg = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc = _RAND_31[38:0];
  _RAND_32 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target = _RAND_32[38:0];
  _RAND_33 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  wbu_io_in_bits_r_isMMIO = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3 = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  wbu_io_in_bits_r_isExit = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_465_valid_reg = _RAND_43[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (io_flush[0]) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (io_flush[1]) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
  end
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  line_466_clock;
  wire  line_466_reset;
  wire  line_466_valid;
  reg  line_466_valid_reg;
  wire  line_467_clock;
  wire  line_467_reset;
  wire  line_467_valid;
  reg  line_467_valid_reg;
  wire  line_468_clock;
  wire  line_468_reset;
  wire  line_468_valid;
  reg  line_468_valid_reg;
  wire  line_469_clock;
  wire  line_469_reset;
  wire  line_469_valid;
  reg  line_469_valid_reg;
  wire  line_470_clock;
  wire  line_470_reset;
  wire  line_470_valid;
  reg  line_470_valid_reg;
  wire  line_471_clock;
  wire  line_471_reset;
  wire  line_471_valid;
  reg  line_471_valid_reg;
  wire  line_472_clock;
  wire  line_472_reset;
  wire  line_472_valid;
  reg  line_472_valid_reg;
  wire  line_473_clock;
  wire  line_473_reset;
  wire  line_473_valid;
  reg  line_473_valid_reg;
  wire  line_474_clock;
  wire  line_474_reset;
  wire  line_474_valid;
  reg  line_474_valid_reg;
  wire  line_475_clock;
  wire  line_475_reset;
  wire  line_475_valid;
  reg  line_475_valid_reg;
  wire  line_476_clock;
  wire  line_476_reset;
  wire  line_476_valid;
  reg  line_476_valid_reg;
  wire  line_477_clock;
  wire  line_477_reset;
  wire  line_477_valid;
  reg  line_477_valid_reg;
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & wantsLock; // @[src/main/scala/chisel3/util/Arbiter.scala 64:22]
  wire  line_478_clock;
  wire  line_478_reset;
  wire  line_478_valid;
  reg  line_478_valid_reg;
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_479_clock;
  wire  line_479_reset;
  wire  line_479_valid;
  reg  line_479_valid_reg;
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  line_480_clock;
  wire  line_480_reset;
  wire  line_480_valid;
  reg  line_480_valid_reg;
  GEN_w1_line #(.COVER_INDEX(466)) line_466 (
    .clock(line_466_clock),
    .reset(line_466_reset),
    .valid(line_466_valid)
  );
  GEN_w1_line #(.COVER_INDEX(467)) line_467 (
    .clock(line_467_clock),
    .reset(line_467_reset),
    .valid(line_467_valid)
  );
  GEN_w1_line #(.COVER_INDEX(468)) line_468 (
    .clock(line_468_clock),
    .reset(line_468_reset),
    .valid(line_468_valid)
  );
  GEN_w1_line #(.COVER_INDEX(469)) line_469 (
    .clock(line_469_clock),
    .reset(line_469_reset),
    .valid(line_469_valid)
  );
  GEN_w1_line #(.COVER_INDEX(470)) line_470 (
    .clock(line_470_clock),
    .reset(line_470_reset),
    .valid(line_470_valid)
  );
  GEN_w1_line #(.COVER_INDEX(471)) line_471 (
    .clock(line_471_clock),
    .reset(line_471_reset),
    .valid(line_471_valid)
  );
  GEN_w1_line #(.COVER_INDEX(472)) line_472 (
    .clock(line_472_clock),
    .reset(line_472_reset),
    .valid(line_472_valid)
  );
  GEN_w1_line #(.COVER_INDEX(473)) line_473 (
    .clock(line_473_clock),
    .reset(line_473_reset),
    .valid(line_473_valid)
  );
  GEN_w1_line #(.COVER_INDEX(474)) line_474 (
    .clock(line_474_clock),
    .reset(line_474_reset),
    .valid(line_474_valid)
  );
  GEN_w1_line #(.COVER_INDEX(475)) line_475 (
    .clock(line_475_clock),
    .reset(line_475_reset),
    .valid(line_475_valid)
  );
  GEN_w1_line #(.COVER_INDEX(476)) line_476 (
    .clock(line_476_clock),
    .reset(line_476_reset),
    .valid(line_476_valid)
  );
  GEN_w1_line #(.COVER_INDEX(477)) line_477 (
    .clock(line_477_clock),
    .reset(line_477_reset),
    .valid(line_477_valid)
  );
  GEN_w1_line #(.COVER_INDEX(478)) line_478 (
    .clock(line_478_clock),
    .reset(line_478_reset),
    .valid(line_478_valid)
  );
  GEN_w1_line #(.COVER_INDEX(479)) line_479 (
    .clock(line_479_clock),
    .reset(line_479_reset),
    .valid(line_479_valid)
  );
  GEN_w1_line #(.COVER_INDEX(480)) line_480 (
    .clock(line_480_clock),
    .reset(line_480_reset),
    .valid(line_480_valid)
  );
  assign line_466_clock = clock;
  assign line_466_reset = reset;
  assign line_466_valid = ~io_chosen ^ line_466_valid_reg;
  assign line_467_clock = clock;
  assign line_467_reset = reset;
  assign line_467_valid = io_chosen ^ line_467_valid_reg;
  assign line_468_clock = clock;
  assign line_468_reset = reset;
  assign line_468_valid = ~io_chosen ^ line_468_valid_reg;
  assign line_469_clock = clock;
  assign line_469_reset = reset;
  assign line_469_valid = io_chosen ^ line_469_valid_reg;
  assign line_470_clock = clock;
  assign line_470_reset = reset;
  assign line_470_valid = ~io_chosen ^ line_470_valid_reg;
  assign line_471_clock = clock;
  assign line_471_reset = reset;
  assign line_471_valid = io_chosen ^ line_471_valid_reg;
  assign line_472_clock = clock;
  assign line_472_reset = reset;
  assign line_472_valid = ~io_chosen ^ line_472_valid_reg;
  assign line_473_clock = clock;
  assign line_473_reset = reset;
  assign line_473_valid = io_chosen ^ line_473_valid_reg;
  assign line_474_clock = clock;
  assign line_474_reset = reset;
  assign line_474_valid = ~io_chosen ^ line_474_valid_reg;
  assign line_475_clock = clock;
  assign line_475_reset = reset;
  assign line_475_valid = io_chosen ^ line_475_valid_reg;
  assign line_476_clock = clock;
  assign line_476_reset = reset;
  assign line_476_valid = ~io_chosen ^ line_476_valid_reg;
  assign line_477_clock = clock;
  assign line_477_reset = reset;
  assign line_477_valid = io_chosen ^ line_477_valid_reg;
  assign line_478_clock = clock;
  assign line_478_reset = reset;
  assign line_478_valid = _T_1 ^ line_478_valid_reg;
  assign line_479_clock = clock;
  assign line_479_reset = reset;
  assign line_479_valid = locked ^ line_479_valid_reg;
  assign line_480_clock = clock;
  assign line_480_reset = reset;
  assign line_480_valid = io_in_0_valid ^ line_480_valid_reg;
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    line_466_valid_reg <= ~io_chosen;
    line_467_valid_reg <= io_chosen;
    line_468_valid_reg <= ~io_chosen;
    line_469_valid_reg <= io_chosen;
    line_470_valid_reg <= ~io_chosen;
    line_471_valid_reg <= io_chosen;
    line_472_valid_reg <= ~io_chosen;
    line_473_valid_reg <= io_chosen;
    line_474_valid_reg <= ~io_chosen;
    line_475_valid_reg <= io_chosen;
    line_476_valid_reg <= ~io_chosen;
    line_477_valid_reg <= io_chosen;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    line_478_valid_reg <= _T_1;
    line_479_valid_reg <= locked;
    line_480_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_466_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_467_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_468_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_469_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_470_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_471_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_472_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_473_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_474_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_475_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_476_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_477_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lockCount_value = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  lockIdx = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_478_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_479_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_480_valid_reg = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (locked) begin
      cover(1'h1);
    end
    //
    if (io_in_0_valid) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:29]
  wire  _T_12 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_481_clock;
  wire  line_481_reset;
  wire  line_481_valid;
  reg  line_481_valid_reg;
  wire  _T_13 = ~(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_482_clock;
  wire  line_482_reset;
  wire  line_482_valid;
  reg  line_482_valid_reg;
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  line_483_clock;
  wire  line_483_reset;
  wire  line_483_valid;
  reg  line_483_valid_reg;
  wire  line_484_clock;
  wire  line_484_reset;
  wire  line_484_valid;
  reg  line_484_valid_reg;
  wire  line_485_clock;
  wire  line_485_reset;
  wire  line_485_valid;
  reg  line_485_valid_reg;
  wire  line_486_clock;
  wire  line_486_reset;
  wire  line_486_valid;
  reg  line_486_valid_reg;
  wire  _T_14 = 2'h0 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_487_clock;
  wire  line_487_reset;
  wire  line_487_valid;
  reg  line_487_valid_reg;
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_488_clock;
  wire  line_488_reset;
  wire  line_488_valid;
  reg  line_488_valid_reg;
  wire  line_489_clock;
  wire  line_489_reset;
  wire  line_489_valid;
  reg  line_489_valid_reg;
  wire  line_490_clock;
  wire  line_490_reset;
  wire  line_490_valid;
  reg  line_490_valid_reg;
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire  _T_23 = _T_21 | _T_22; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:47]
  wire  line_491_clock;
  wire  line_491_reset;
  wire  line_491_valid;
  reg  line_491_valid_reg;
  wire [1:0] _GEN_21 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  line_492_clock;
  wire  line_492_reset;
  wire  line_492_valid;
  reg  line_492_valid_reg;
  wire  _T_24 = 2'h1 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_493_clock;
  wire  line_493_reset;
  wire  line_493_valid;
  reg  line_493_valid_reg;
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire  _T_27 = _T_25 & _T_26; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:48]
  wire  line_494_clock;
  wire  line_494_reset;
  wire  line_494_valid;
  reg  line_494_valid_reg;
  wire  line_495_clock;
  wire  line_495_reset;
  wire  line_495_valid;
  reg  line_495_valid_reg;
  wire  _T_28 = 2'h2 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_496_clock;
  wire  line_496_reset;
  wire  line_496_valid;
  reg  line_496_valid_reg;
  wire  line_497_clock;
  wire  line_497_reset;
  wire  line_497_valid;
  reg  line_497_valid_reg;
  wire [1:0] _GEN_26 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w1_line #(.COVER_INDEX(481)) line_481 (
    .clock(line_481_clock),
    .reset(line_481_reset),
    .valid(line_481_valid)
  );
  GEN_w1_line #(.COVER_INDEX(482)) line_482 (
    .clock(line_482_clock),
    .reset(line_482_reset),
    .valid(line_482_valid)
  );
  GEN_w1_line #(.COVER_INDEX(483)) line_483 (
    .clock(line_483_clock),
    .reset(line_483_reset),
    .valid(line_483_valid)
  );
  GEN_w1_line #(.COVER_INDEX(484)) line_484 (
    .clock(line_484_clock),
    .reset(line_484_reset),
    .valid(line_484_valid)
  );
  GEN_w1_line #(.COVER_INDEX(485)) line_485 (
    .clock(line_485_clock),
    .reset(line_485_reset),
    .valid(line_485_valid)
  );
  GEN_w1_line #(.COVER_INDEX(486)) line_486 (
    .clock(line_486_clock),
    .reset(line_486_reset),
    .valid(line_486_valid)
  );
  GEN_w1_line #(.COVER_INDEX(487)) line_487 (
    .clock(line_487_clock),
    .reset(line_487_reset),
    .valid(line_487_valid)
  );
  GEN_w1_line #(.COVER_INDEX(488)) line_488 (
    .clock(line_488_clock),
    .reset(line_488_reset),
    .valid(line_488_valid)
  );
  GEN_w1_line #(.COVER_INDEX(489)) line_489 (
    .clock(line_489_clock),
    .reset(line_489_reset),
    .valid(line_489_valid)
  );
  GEN_w1_line #(.COVER_INDEX(490)) line_490 (
    .clock(line_490_clock),
    .reset(line_490_reset),
    .valid(line_490_valid)
  );
  GEN_w1_line #(.COVER_INDEX(491)) line_491 (
    .clock(line_491_clock),
    .reset(line_491_reset),
    .valid(line_491_valid)
  );
  GEN_w1_line #(.COVER_INDEX(492)) line_492 (
    .clock(line_492_clock),
    .reset(line_492_reset),
    .valid(line_492_valid)
  );
  GEN_w1_line #(.COVER_INDEX(493)) line_493 (
    .clock(line_493_clock),
    .reset(line_493_reset),
    .valid(line_493_valid)
  );
  GEN_w1_line #(.COVER_INDEX(494)) line_494 (
    .clock(line_494_clock),
    .reset(line_494_reset),
    .valid(line_494_valid)
  );
  GEN_w1_line #(.COVER_INDEX(495)) line_495 (
    .clock(line_495_clock),
    .reset(line_495_reset),
    .valid(line_495_valid)
  );
  GEN_w1_line #(.COVER_INDEX(496)) line_496 (
    .clock(line_496_clock),
    .reset(line_496_reset),
    .valid(line_496_valid)
  );
  GEN_w1_line #(.COVER_INDEX(497)) line_497 (
    .clock(line_497_clock),
    .reset(line_497_reset),
    .valid(line_497_valid)
  );
  assign line_481_clock = clock;
  assign line_481_reset = reset;
  assign line_481_valid = _T_12 ^ line_481_valid_reg;
  assign line_482_clock = clock;
  assign line_482_reset = reset;
  assign line_482_valid = _T_13 ^ line_482_valid_reg;
  assign line_483_clock = clock;
  assign line_483_reset = reset;
  assign line_483_valid = ~inflightSrc ^ line_483_valid_reg;
  assign line_484_clock = clock;
  assign line_484_reset = reset;
  assign line_484_valid = inflightSrc ^ line_484_valid_reg;
  assign line_485_clock = clock;
  assign line_485_reset = reset;
  assign line_485_valid = ~inflightSrc ^ line_485_valid_reg;
  assign line_486_clock = clock;
  assign line_486_reset = reset;
  assign line_486_valid = inflightSrc ^ line_486_valid_reg;
  assign line_487_clock = clock;
  assign line_487_reset = reset;
  assign line_487_valid = _T_14 ^ line_487_valid_reg;
  assign line_488_clock = clock;
  assign line_488_reset = reset;
  assign line_488_valid = _T_15 ^ line_488_valid_reg;
  assign line_489_clock = clock;
  assign line_489_reset = reset;
  assign line_489_valid = _T_4 ^ line_489_valid_reg;
  assign line_490_clock = clock;
  assign line_490_reset = reset;
  assign line_490_valid = _T_4 ^ line_490_valid_reg;
  assign line_491_clock = clock;
  assign line_491_reset = reset;
  assign line_491_valid = _T_23 ^ line_491_valid_reg;
  assign line_492_clock = clock;
  assign line_492_reset = reset;
  assign line_492_valid = _T_14 ^ line_492_valid_reg;
  assign line_493_clock = clock;
  assign line_493_reset = reset;
  assign line_493_valid = _T_24 ^ line_493_valid_reg;
  assign line_494_clock = clock;
  assign line_494_reset = reset;
  assign line_494_valid = _T_27 ^ line_494_valid_reg;
  assign line_495_clock = clock;
  assign line_495_reset = reset;
  assign line_495_valid = _T_24 ^ line_495_valid_reg;
  assign line_496_clock = clock;
  assign line_496_reset = reset;
  assign line_496_valid = _T_28 ^ line_496_valid_reg;
  assign line_497_clock = clock;
  assign line_497_reset = reset;
  assign line_497_valid = _T_25 ^ line_497_valid_reg;
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_21;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_26;
    end
    line_481_valid_reg <= _T_12;
    line_482_valid_reg <= _T_13;
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    line_483_valid_reg <= ~inflightSrc;
    line_484_valid_reg <= inflightSrc;
    line_485_valid_reg <= ~inflightSrc;
    line_486_valid_reg <= inflightSrc;
    line_487_valid_reg <= _T_14;
    line_488_valid_reg <= _T_15;
    line_489_valid_reg <= _T_4;
    line_490_valid_reg <= _T_4;
    line_491_valid_reg <= _T_23;
    line_492_valid_reg <= _T_14;
    line_493_valid_reg <= _T_24;
    line_494_valid_reg <= _T_27;
    line_495_valid_reg <= _T_24;
    line_496_valid_reg <= _T_28;
    line_497_valid_reg <= _T_25;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_481_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_482_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  inflightSrc = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_483_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_484_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_485_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_486_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_487_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_488_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_489_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_490_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_491_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_492_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_493_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_494_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_495_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_496_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_497_valid_reg = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_12 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (~inflightSrc) begin
      cover(1'h1);
    end
    //
    if (inflightSrc) begin
      cover(1'h1);
    end
    //
    if (~inflightSrc) begin
      cover(1'h1);
    end
    //
    if (inflightSrc) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_4) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5 & _T_23) begin
      cover(1'h1);
    end
    //
    if (~_T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24 & _T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28 & _T_25) begin
      cover(1'h1);
    end
  end
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_2_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_2_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_2_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_3_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [1:0]  io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  line_498_clock;
  wire  line_498_reset;
  wire  line_498_valid;
  reg  line_498_valid_reg;
  wire  line_499_clock;
  wire  line_499_reset;
  wire  line_499_valid;
  reg  line_499_valid_reg;
  wire  _GEN_30 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  line_500_clock;
  wire  line_500_reset;
  wire  line_500_valid;
  reg  line_500_valid_reg;
  wire  _GEN_31 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_30; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  line_501_clock;
  wire  line_501_reset;
  wire  line_501_valid;
  reg  line_501_valid_reg;
  wire  line_502_clock;
  wire  line_502_reset;
  wire  line_502_valid;
  reg  line_502_valid_reg;
  wire  line_503_clock;
  wire  line_503_reset;
  wire  line_503_valid;
  reg  line_503_valid_reg;
  wire [31:0] _GEN_34 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_504_clock;
  wire  line_504_reset;
  wire  line_504_valid;
  reg  line_504_valid_reg;
  wire [31:0] _GEN_35 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_34; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_505_clock;
  wire  line_505_reset;
  wire  line_505_valid;
  reg  line_505_valid_reg;
  wire  line_506_clock;
  wire  line_506_reset;
  wire  line_506_valid;
  reg  line_506_valid_reg;
  wire  line_507_clock;
  wire  line_507_reset;
  wire  line_507_valid;
  reg  line_507_valid_reg;
  wire [2:0] _GEN_38 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_508_clock;
  wire  line_508_reset;
  wire  line_508_valid;
  reg  line_508_valid_reg;
  wire [2:0] _GEN_39 = 2'h2 == io_chosen ? 3'h3 : _GEN_38; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_509_clock;
  wire  line_509_reset;
  wire  line_509_valid;
  reg  line_509_valid_reg;
  wire  line_510_clock;
  wire  line_510_reset;
  wire  line_510_valid;
  reg  line_510_valid_reg;
  wire  line_511_clock;
  wire  line_511_reset;
  wire  line_511_valid;
  reg  line_511_valid_reg;
  wire [3:0] _GEN_42 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_512_clock;
  wire  line_512_reset;
  wire  line_512_valid;
  reg  line_512_valid_reg;
  wire [3:0] _GEN_43 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_42; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_513_clock;
  wire  line_513_reset;
  wire  line_513_valid;
  reg  line_513_valid_reg;
  wire  line_514_clock;
  wire  line_514_reset;
  wire  line_514_valid;
  reg  line_514_valid_reg;
  wire  line_515_clock;
  wire  line_515_reset;
  wire  line_515_valid;
  reg  line_515_valid_reg;
  wire [7:0] _GEN_46 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_516_clock;
  wire  line_516_reset;
  wire  line_516_valid;
  reg  line_516_valid_reg;
  wire [7:0] _GEN_47 = 2'h2 == io_chosen ? 8'hff : _GEN_46; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_517_clock;
  wire  line_517_reset;
  wire  line_517_valid;
  reg  line_517_valid_reg;
  wire  line_518_clock;
  wire  line_518_reset;
  wire  line_518_valid;
  reg  line_518_valid_reg;
  wire  line_519_clock;
  wire  line_519_reset;
  wire  line_519_valid;
  reg  line_519_valid_reg;
  wire [63:0] _GEN_50 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_520_clock;
  wire  line_520_reset;
  wire  line_520_valid;
  reg  line_520_valid_reg;
  wire [63:0] _GEN_51 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_50; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire  line_521_clock;
  wire  line_521_reset;
  wire  line_521_valid;
  reg  line_521_valid_reg;
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & wantsLock; // @[src/main/scala/chisel3/util/Arbiter.scala 64:22]
  wire  line_522_clock;
  wire  line_522_reset;
  wire  line_522_valid;
  reg  line_522_valid_reg;
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_523_clock;
  wire  line_523_reset;
  wire  line_523_valid;
  reg  line_523_valid_reg;
  wire [1:0] _GEN_56 = io_in_2_valid ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire [1:0] _GEN_57 = io_in_1_valid ? 2'h1 : _GEN_56; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire [1:0] io_chosen_choice = io_in_0_valid ? 2'h0 : _GEN_57; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire  _T_4 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_6 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_3_ready_T_1 = locked ? lockIdx == 2'h3 : _T_6; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  line_524_clock;
  wire  line_524_reset;
  wire  line_524_valid;
  reg  line_524_valid_reg;
  wire  line_525_clock;
  wire  line_525_reset;
  wire  line_525_valid;
  reg  line_525_valid_reg;
  wire  line_526_clock;
  wire  line_526_reset;
  wire  line_526_valid;
  reg  line_526_valid_reg;
  GEN_w1_line #(.COVER_INDEX(498)) line_498 (
    .clock(line_498_clock),
    .reset(line_498_reset),
    .valid(line_498_valid)
  );
  GEN_w1_line #(.COVER_INDEX(499)) line_499 (
    .clock(line_499_clock),
    .reset(line_499_reset),
    .valid(line_499_valid)
  );
  GEN_w1_line #(.COVER_INDEX(500)) line_500 (
    .clock(line_500_clock),
    .reset(line_500_reset),
    .valid(line_500_valid)
  );
  GEN_w1_line #(.COVER_INDEX(501)) line_501 (
    .clock(line_501_clock),
    .reset(line_501_reset),
    .valid(line_501_valid)
  );
  GEN_w1_line #(.COVER_INDEX(502)) line_502 (
    .clock(line_502_clock),
    .reset(line_502_reset),
    .valid(line_502_valid)
  );
  GEN_w1_line #(.COVER_INDEX(503)) line_503 (
    .clock(line_503_clock),
    .reset(line_503_reset),
    .valid(line_503_valid)
  );
  GEN_w1_line #(.COVER_INDEX(504)) line_504 (
    .clock(line_504_clock),
    .reset(line_504_reset),
    .valid(line_504_valid)
  );
  GEN_w1_line #(.COVER_INDEX(505)) line_505 (
    .clock(line_505_clock),
    .reset(line_505_reset),
    .valid(line_505_valid)
  );
  GEN_w1_line #(.COVER_INDEX(506)) line_506 (
    .clock(line_506_clock),
    .reset(line_506_reset),
    .valid(line_506_valid)
  );
  GEN_w1_line #(.COVER_INDEX(507)) line_507 (
    .clock(line_507_clock),
    .reset(line_507_reset),
    .valid(line_507_valid)
  );
  GEN_w1_line #(.COVER_INDEX(508)) line_508 (
    .clock(line_508_clock),
    .reset(line_508_reset),
    .valid(line_508_valid)
  );
  GEN_w1_line #(.COVER_INDEX(509)) line_509 (
    .clock(line_509_clock),
    .reset(line_509_reset),
    .valid(line_509_valid)
  );
  GEN_w1_line #(.COVER_INDEX(510)) line_510 (
    .clock(line_510_clock),
    .reset(line_510_reset),
    .valid(line_510_valid)
  );
  GEN_w1_line #(.COVER_INDEX(511)) line_511 (
    .clock(line_511_clock),
    .reset(line_511_reset),
    .valid(line_511_valid)
  );
  GEN_w1_line #(.COVER_INDEX(512)) line_512 (
    .clock(line_512_clock),
    .reset(line_512_reset),
    .valid(line_512_valid)
  );
  GEN_w1_line #(.COVER_INDEX(513)) line_513 (
    .clock(line_513_clock),
    .reset(line_513_reset),
    .valid(line_513_valid)
  );
  GEN_w1_line #(.COVER_INDEX(514)) line_514 (
    .clock(line_514_clock),
    .reset(line_514_reset),
    .valid(line_514_valid)
  );
  GEN_w1_line #(.COVER_INDEX(515)) line_515 (
    .clock(line_515_clock),
    .reset(line_515_reset),
    .valid(line_515_valid)
  );
  GEN_w1_line #(.COVER_INDEX(516)) line_516 (
    .clock(line_516_clock),
    .reset(line_516_reset),
    .valid(line_516_valid)
  );
  GEN_w1_line #(.COVER_INDEX(517)) line_517 (
    .clock(line_517_clock),
    .reset(line_517_reset),
    .valid(line_517_valid)
  );
  GEN_w1_line #(.COVER_INDEX(518)) line_518 (
    .clock(line_518_clock),
    .reset(line_518_reset),
    .valid(line_518_valid)
  );
  GEN_w1_line #(.COVER_INDEX(519)) line_519 (
    .clock(line_519_clock),
    .reset(line_519_reset),
    .valid(line_519_valid)
  );
  GEN_w1_line #(.COVER_INDEX(520)) line_520 (
    .clock(line_520_clock),
    .reset(line_520_reset),
    .valid(line_520_valid)
  );
  GEN_w1_line #(.COVER_INDEX(521)) line_521 (
    .clock(line_521_clock),
    .reset(line_521_reset),
    .valid(line_521_valid)
  );
  GEN_w1_line #(.COVER_INDEX(522)) line_522 (
    .clock(line_522_clock),
    .reset(line_522_reset),
    .valid(line_522_valid)
  );
  GEN_w1_line #(.COVER_INDEX(523)) line_523 (
    .clock(line_523_clock),
    .reset(line_523_reset),
    .valid(line_523_valid)
  );
  GEN_w1_line #(.COVER_INDEX(524)) line_524 (
    .clock(line_524_clock),
    .reset(line_524_reset),
    .valid(line_524_valid)
  );
  GEN_w1_line #(.COVER_INDEX(525)) line_525 (
    .clock(line_525_clock),
    .reset(line_525_reset),
    .valid(line_525_valid)
  );
  GEN_w1_line #(.COVER_INDEX(526)) line_526 (
    .clock(line_526_clock),
    .reset(line_526_reset),
    .valid(line_526_valid)
  );
  assign line_498_clock = clock;
  assign line_498_reset = reset;
  assign line_498_valid = 2'h0 == io_chosen ^ line_498_valid_reg;
  assign line_499_clock = clock;
  assign line_499_reset = reset;
  assign line_499_valid = 2'h1 == io_chosen ^ line_499_valid_reg;
  assign line_500_clock = clock;
  assign line_500_reset = reset;
  assign line_500_valid = 2'h2 == io_chosen ^ line_500_valid_reg;
  assign line_501_clock = clock;
  assign line_501_reset = reset;
  assign line_501_valid = 2'h3 == io_chosen ^ line_501_valid_reg;
  assign line_502_clock = clock;
  assign line_502_reset = reset;
  assign line_502_valid = 2'h0 == io_chosen ^ line_502_valid_reg;
  assign line_503_clock = clock;
  assign line_503_reset = reset;
  assign line_503_valid = 2'h1 == io_chosen ^ line_503_valid_reg;
  assign line_504_clock = clock;
  assign line_504_reset = reset;
  assign line_504_valid = 2'h2 == io_chosen ^ line_504_valid_reg;
  assign line_505_clock = clock;
  assign line_505_reset = reset;
  assign line_505_valid = 2'h3 == io_chosen ^ line_505_valid_reg;
  assign line_506_clock = clock;
  assign line_506_reset = reset;
  assign line_506_valid = 2'h0 == io_chosen ^ line_506_valid_reg;
  assign line_507_clock = clock;
  assign line_507_reset = reset;
  assign line_507_valid = 2'h1 == io_chosen ^ line_507_valid_reg;
  assign line_508_clock = clock;
  assign line_508_reset = reset;
  assign line_508_valid = 2'h2 == io_chosen ^ line_508_valid_reg;
  assign line_509_clock = clock;
  assign line_509_reset = reset;
  assign line_509_valid = 2'h3 == io_chosen ^ line_509_valid_reg;
  assign line_510_clock = clock;
  assign line_510_reset = reset;
  assign line_510_valid = 2'h0 == io_chosen ^ line_510_valid_reg;
  assign line_511_clock = clock;
  assign line_511_reset = reset;
  assign line_511_valid = 2'h1 == io_chosen ^ line_511_valid_reg;
  assign line_512_clock = clock;
  assign line_512_reset = reset;
  assign line_512_valid = 2'h2 == io_chosen ^ line_512_valid_reg;
  assign line_513_clock = clock;
  assign line_513_reset = reset;
  assign line_513_valid = 2'h3 == io_chosen ^ line_513_valid_reg;
  assign line_514_clock = clock;
  assign line_514_reset = reset;
  assign line_514_valid = 2'h0 == io_chosen ^ line_514_valid_reg;
  assign line_515_clock = clock;
  assign line_515_reset = reset;
  assign line_515_valid = 2'h1 == io_chosen ^ line_515_valid_reg;
  assign line_516_clock = clock;
  assign line_516_reset = reset;
  assign line_516_valid = 2'h2 == io_chosen ^ line_516_valid_reg;
  assign line_517_clock = clock;
  assign line_517_reset = reset;
  assign line_517_valid = 2'h3 == io_chosen ^ line_517_valid_reg;
  assign line_518_clock = clock;
  assign line_518_reset = reset;
  assign line_518_valid = 2'h0 == io_chosen ^ line_518_valid_reg;
  assign line_519_clock = clock;
  assign line_519_reset = reset;
  assign line_519_valid = 2'h1 == io_chosen ^ line_519_valid_reg;
  assign line_520_clock = clock;
  assign line_520_reset = reset;
  assign line_520_valid = 2'h2 == io_chosen ^ line_520_valid_reg;
  assign line_521_clock = clock;
  assign line_521_reset = reset;
  assign line_521_valid = 2'h3 == io_chosen ^ line_521_valid_reg;
  assign line_522_clock = clock;
  assign line_522_reset = reset;
  assign line_522_valid = _T_1 ^ line_522_valid_reg;
  assign line_523_clock = clock;
  assign line_523_reset = reset;
  assign line_523_valid = locked ^ line_523_valid_reg;
  assign line_524_clock = clock;
  assign line_524_reset = reset;
  assign line_524_valid = io_in_2_valid ^ line_524_valid_reg;
  assign line_525_clock = clock;
  assign line_525_reset = reset;
  assign line_525_valid = io_in_1_valid ^ line_525_valid_reg;
  assign line_526_clock = clock;
  assign line_526_reset = reset;
  assign line_526_valid = io_in_0_valid ^ line_526_valid_reg;
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_3_ready = _io_in_3_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = 2'h3 == io_chosen ? 1'h0 : _GEN_31; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? 32'h0 : _GEN_35; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? 3'h0 : _GEN_39; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? 4'h0 : _GEN_43; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? 8'h0 : _GEN_47; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? 64'h0 : _GEN_51; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    line_498_valid_reg <= 2'h0 == io_chosen;
    line_499_valid_reg <= 2'h1 == io_chosen;
    line_500_valid_reg <= 2'h2 == io_chosen;
    line_501_valid_reg <= 2'h3 == io_chosen;
    line_502_valid_reg <= 2'h0 == io_chosen;
    line_503_valid_reg <= 2'h1 == io_chosen;
    line_504_valid_reg <= 2'h2 == io_chosen;
    line_505_valid_reg <= 2'h3 == io_chosen;
    line_506_valid_reg <= 2'h0 == io_chosen;
    line_507_valid_reg <= 2'h1 == io_chosen;
    line_508_valid_reg <= 2'h2 == io_chosen;
    line_509_valid_reg <= 2'h3 == io_chosen;
    line_510_valid_reg <= 2'h0 == io_chosen;
    line_511_valid_reg <= 2'h1 == io_chosen;
    line_512_valid_reg <= 2'h2 == io_chosen;
    line_513_valid_reg <= 2'h3 == io_chosen;
    line_514_valid_reg <= 2'h0 == io_chosen;
    line_515_valid_reg <= 2'h1 == io_chosen;
    line_516_valid_reg <= 2'h2 == io_chosen;
    line_517_valid_reg <= 2'h3 == io_chosen;
    line_518_valid_reg <= 2'h0 == io_chosen;
    line_519_valid_reg <= 2'h1 == io_chosen;
    line_520_valid_reg <= 2'h2 == io_chosen;
    line_521_valid_reg <= 2'h3 == io_chosen;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    line_522_valid_reg <= _T_1;
    line_523_valid_reg <= locked;
    line_524_valid_reg <= io_in_2_valid;
    line_525_valid_reg <= io_in_1_valid;
    line_526_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_498_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_499_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_500_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_501_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_502_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_503_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_504_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_505_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_506_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_507_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_508_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_509_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_510_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_511_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_512_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_513_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_514_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_515_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_516_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_517_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_518_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_519_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_520_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_521_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lockCount_value = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  lockIdx = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  line_522_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_523_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_524_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_525_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_526_valid_reg = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h0 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h1 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h2 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (2'h3 == io_chosen) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (locked) begin
      cover(1'h1);
    end
    //
    if (io_in_2_valid) begin
      cover(1'h1);
    end
    //
    if (io_in_1_valid) begin
      cover(1'h1);
    end
    //
    if (io_in_0_valid) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_0_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [1:0] inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:29]
  wire  _T_12 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_527_clock;
  wire  line_527_reset;
  wire  line_527_valid;
  reg  line_527_valid_reg;
  wire  _T_13 = ~(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_528_clock;
  wire  line_528_reset;
  wire  line_528_valid;
  reg  line_528_valid_reg;
  reg [1:0] inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  line_529_clock;
  wire  line_529_reset;
  wire  line_529_valid;
  reg  line_529_valid_reg;
  wire  line_530_clock;
  wire  line_530_reset;
  wire  line_530_valid;
  reg  line_530_valid_reg;
  wire  line_531_clock;
  wire  line_531_reset;
  wire  line_531_valid;
  reg  line_531_valid_reg;
  wire  line_532_clock;
  wire  line_532_reset;
  wire  line_532_valid;
  reg  line_532_valid_reg;
  wire  line_533_clock;
  wire  line_533_reset;
  wire  line_533_valid;
  reg  line_533_valid_reg;
  wire  line_534_clock;
  wire  line_534_reset;
  wire  line_534_valid;
  reg  line_534_valid_reg;
  wire  line_535_clock;
  wire  line_535_reset;
  wire  line_535_valid;
  reg  line_535_valid_reg;
  wire  line_536_clock;
  wire  line_536_reset;
  wire  line_536_valid;
  reg  line_536_valid_reg;
  wire  _T_14 = 2'h0 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_537_clock;
  wire  line_537_reset;
  wire  line_537_valid;
  reg  line_537_valid_reg;
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_538_clock;
  wire  line_538_reset;
  wire  line_538_valid;
  reg  line_538_valid_reg;
  wire  line_539_clock;
  wire  line_539_reset;
  wire  line_539_valid;
  reg  line_539_valid_reg;
  wire  line_540_clock;
  wire  line_540_reset;
  wire  line_540_valid;
  reg  line_540_valid_reg;
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire  _T_23 = _T_21 | _T_22; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:47]
  wire  line_541_clock;
  wire  line_541_reset;
  wire  line_541_valid;
  reg  line_541_valid_reg;
  wire [1:0] _GEN_29 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  line_542_clock;
  wire  line_542_reset;
  wire  line_542_valid;
  reg  line_542_valid_reg;
  wire  _T_24 = 2'h1 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_543_clock;
  wire  line_543_reset;
  wire  line_543_valid;
  reg  line_543_valid_reg;
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire  _T_27 = _T_25 & _T_26; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:48]
  wire  line_544_clock;
  wire  line_544_reset;
  wire  line_544_valid;
  reg  line_544_valid_reg;
  wire  line_545_clock;
  wire  line_545_reset;
  wire  line_545_valid;
  reg  line_545_valid_reg;
  wire  _T_28 = 2'h2 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_546_clock;
  wire  line_546_reset;
  wire  line_546_valid;
  reg  line_546_valid_reg;
  wire  line_547_clock;
  wire  line_547_reset;
  wire  line_547_valid;
  reg  line_547_valid_reg;
  wire [1:0] _GEN_34 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter_1 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w1_line #(.COVER_INDEX(527)) line_527 (
    .clock(line_527_clock),
    .reset(line_527_reset),
    .valid(line_527_valid)
  );
  GEN_w1_line #(.COVER_INDEX(528)) line_528 (
    .clock(line_528_clock),
    .reset(line_528_reset),
    .valid(line_528_valid)
  );
  GEN_w1_line #(.COVER_INDEX(529)) line_529 (
    .clock(line_529_clock),
    .reset(line_529_reset),
    .valid(line_529_valid)
  );
  GEN_w1_line #(.COVER_INDEX(530)) line_530 (
    .clock(line_530_clock),
    .reset(line_530_reset),
    .valid(line_530_valid)
  );
  GEN_w1_line #(.COVER_INDEX(531)) line_531 (
    .clock(line_531_clock),
    .reset(line_531_reset),
    .valid(line_531_valid)
  );
  GEN_w1_line #(.COVER_INDEX(532)) line_532 (
    .clock(line_532_clock),
    .reset(line_532_reset),
    .valid(line_532_valid)
  );
  GEN_w1_line #(.COVER_INDEX(533)) line_533 (
    .clock(line_533_clock),
    .reset(line_533_reset),
    .valid(line_533_valid)
  );
  GEN_w1_line #(.COVER_INDEX(534)) line_534 (
    .clock(line_534_clock),
    .reset(line_534_reset),
    .valid(line_534_valid)
  );
  GEN_w1_line #(.COVER_INDEX(535)) line_535 (
    .clock(line_535_clock),
    .reset(line_535_reset),
    .valid(line_535_valid)
  );
  GEN_w1_line #(.COVER_INDEX(536)) line_536 (
    .clock(line_536_clock),
    .reset(line_536_reset),
    .valid(line_536_valid)
  );
  GEN_w1_line #(.COVER_INDEX(537)) line_537 (
    .clock(line_537_clock),
    .reset(line_537_reset),
    .valid(line_537_valid)
  );
  GEN_w1_line #(.COVER_INDEX(538)) line_538 (
    .clock(line_538_clock),
    .reset(line_538_reset),
    .valid(line_538_valid)
  );
  GEN_w1_line #(.COVER_INDEX(539)) line_539 (
    .clock(line_539_clock),
    .reset(line_539_reset),
    .valid(line_539_valid)
  );
  GEN_w1_line #(.COVER_INDEX(540)) line_540 (
    .clock(line_540_clock),
    .reset(line_540_reset),
    .valid(line_540_valid)
  );
  GEN_w1_line #(.COVER_INDEX(541)) line_541 (
    .clock(line_541_clock),
    .reset(line_541_reset),
    .valid(line_541_valid)
  );
  GEN_w1_line #(.COVER_INDEX(542)) line_542 (
    .clock(line_542_clock),
    .reset(line_542_reset),
    .valid(line_542_valid)
  );
  GEN_w1_line #(.COVER_INDEX(543)) line_543 (
    .clock(line_543_clock),
    .reset(line_543_reset),
    .valid(line_543_valid)
  );
  GEN_w1_line #(.COVER_INDEX(544)) line_544 (
    .clock(line_544_clock),
    .reset(line_544_reset),
    .valid(line_544_valid)
  );
  GEN_w1_line #(.COVER_INDEX(545)) line_545 (
    .clock(line_545_clock),
    .reset(line_545_reset),
    .valid(line_545_valid)
  );
  GEN_w1_line #(.COVER_INDEX(546)) line_546 (
    .clock(line_546_clock),
    .reset(line_546_reset),
    .valid(line_546_valid)
  );
  GEN_w1_line #(.COVER_INDEX(547)) line_547 (
    .clock(line_547_clock),
    .reset(line_547_reset),
    .valid(line_547_valid)
  );
  assign line_527_clock = clock;
  assign line_527_reset = reset;
  assign line_527_valid = _T_12 ^ line_527_valid_reg;
  assign line_528_clock = clock;
  assign line_528_reset = reset;
  assign line_528_valid = _T_13 ^ line_528_valid_reg;
  assign line_529_clock = clock;
  assign line_529_reset = reset;
  assign line_529_valid = 2'h0 == inflightSrc ^ line_529_valid_reg;
  assign line_530_clock = clock;
  assign line_530_reset = reset;
  assign line_530_valid = 2'h1 == inflightSrc ^ line_530_valid_reg;
  assign line_531_clock = clock;
  assign line_531_reset = reset;
  assign line_531_valid = 2'h2 == inflightSrc ^ line_531_valid_reg;
  assign line_532_clock = clock;
  assign line_532_reset = reset;
  assign line_532_valid = 2'h3 == inflightSrc ^ line_532_valid_reg;
  assign line_533_clock = clock;
  assign line_533_reset = reset;
  assign line_533_valid = 2'h0 == inflightSrc ^ line_533_valid_reg;
  assign line_534_clock = clock;
  assign line_534_reset = reset;
  assign line_534_valid = 2'h1 == inflightSrc ^ line_534_valid_reg;
  assign line_535_clock = clock;
  assign line_535_reset = reset;
  assign line_535_valid = 2'h2 == inflightSrc ^ line_535_valid_reg;
  assign line_536_clock = clock;
  assign line_536_reset = reset;
  assign line_536_valid = 2'h3 == inflightSrc ^ line_536_valid_reg;
  assign line_537_clock = clock;
  assign line_537_reset = reset;
  assign line_537_valid = _T_14 ^ line_537_valid_reg;
  assign line_538_clock = clock;
  assign line_538_reset = reset;
  assign line_538_valid = _T_15 ^ line_538_valid_reg;
  assign line_539_clock = clock;
  assign line_539_reset = reset;
  assign line_539_valid = _T_4 ^ line_539_valid_reg;
  assign line_540_clock = clock;
  assign line_540_reset = reset;
  assign line_540_valid = _T_4 ^ line_540_valid_reg;
  assign line_541_clock = clock;
  assign line_541_reset = reset;
  assign line_541_valid = _T_23 ^ line_541_valid_reg;
  assign line_542_clock = clock;
  assign line_542_reset = reset;
  assign line_542_valid = _T_14 ^ line_542_valid_reg;
  assign line_543_clock = clock;
  assign line_543_reset = reset;
  assign line_543_valid = _T_24 ^ line_543_valid_reg;
  assign line_544_clock = clock;
  assign line_544_reset = reset;
  assign line_544_valid = _T_27 ^ line_544_valid_reg;
  assign line_545_clock = clock;
  assign line_545_reset = reset;
  assign line_545_valid = _T_24 ^ line_545_valid_reg;
  assign line_546_clock = clock;
  assign line_546_reset = reset;
  assign line_546_valid = _T_28 ^ line_546_valid_reg;
  assign line_547_clock = clock;
  assign line_547_reset = reset;
  assign line_547_valid = _T_25 ^ line_547_valid_reg;
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_29;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_34;
    end
    line_527_valid_reg <= _T_12;
    line_528_valid_reg <= _T_13;
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    line_529_valid_reg <= 2'h0 == inflightSrc;
    line_530_valid_reg <= 2'h1 == inflightSrc;
    line_531_valid_reg <= 2'h2 == inflightSrc;
    line_532_valid_reg <= 2'h3 == inflightSrc;
    line_533_valid_reg <= 2'h0 == inflightSrc;
    line_534_valid_reg <= 2'h1 == inflightSrc;
    line_535_valid_reg <= 2'h2 == inflightSrc;
    line_536_valid_reg <= 2'h3 == inflightSrc;
    line_537_valid_reg <= _T_14;
    line_538_valid_reg <= _T_15;
    line_539_valid_reg <= _T_4;
    line_540_valid_reg <= _T_4;
    line_541_valid_reg <= _T_23;
    line_542_valid_reg <= _T_14;
    line_543_valid_reg <= _T_24;
    line_544_valid_reg <= _T_27;
    line_545_valid_reg <= _T_24;
    line_546_valid_reg <= _T_28;
    line_547_valid_reg <= _T_25;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_527_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_528_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  inflightSrc = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  line_529_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_530_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_531_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_532_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_533_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_534_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_535_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_536_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_537_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_538_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_539_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_540_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_541_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_542_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_543_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_544_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_545_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_546_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_547_valid_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_12 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (2'h0 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h1 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h2 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h3 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h0 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h1 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h2 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (2'h3 == inflightSrc) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_4) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5 & _T_23) begin
      cover(1'h1);
    end
    //
    if (~_T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24 & _T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28 & _T_25) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [86:0]  io_in_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [86:0]  io_out_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:20]
  wire  hitExec = hitCheck & ~hitADCheck & hitFlag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:41]
  wire  hitinstrPF = ~hitExec & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 290:52]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  line_548_clock;
  wire  line_548_reset;
  wire  line_548_valid;
  reg  line_548_valid_reg;
  wire  _GEN_42 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
  wire  isFlush = needFlush | io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 314:27]
  wire  _T_1 = io_flush & state != 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 315:17]
  wire  line_549_clock;
  wire  line_549_reset;
  wire  line_549_valid;
  reg  line_549_valid_reg;
  wire  _GEN_43 = io_flush & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26 315:{40,52}]
  wire  _T_3 = _alreadyOutFire_T & needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 316:23]
  wire  line_550_clock;
  wire  line_550_reset;
  wire  line_550_valid;
  reg  line_550_valid_reg;
  wire  _GEN_44 = _alreadyOutFire_T & needFlush ? 1'h0 : _GEN_43; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 316:{37,49}]
  reg  missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  _T_4 = 3'h0 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_551_clock;
  wire  line_551_reset;
  wire  line_551_valid;
  reg  line_551_valid_reg;
  wire  _T_5 = ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 324:13]
  wire  _T_8 = miss & _T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:24]
  wire  line_552_clock;
  wire  line_552_reset;
  wire  line_552_valid;
  reg  line_552_valid_reg;
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  line_553_clock;
  wire  line_553_reset;
  wire  line_553_valid;
  reg  line_553_valid_reg;
  wire  _T_9 = 3'h1 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_554_clock;
  wire  line_554_reset;
  wire  line_554_valid;
  reg  line_554_valid_reg;
  wire  line_555_clock;
  wire  line_555_reset;
  wire  line_555_valid;
  reg  line_555_valid_reg;
  wire  line_556_clock;
  wire  line_556_reset;
  wire  line_556_valid;
  reg  line_556_valid_reg;
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_557_clock;
  wire  line_557_reset;
  wire  line_557_valid;
  reg  line_557_valid_reg;
  wire  line_558_clock;
  wire  line_558_reset;
  wire  line_558_valid;
  reg  line_558_valid_reg;
  wire  line_559_clock;
  wire  line_559_reset;
  wire  line_559_valid;
  reg  line_559_valid_reg;
  wire [2:0] _GEN_55 = raddrCancel ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:29]
  wire  _GEN_56 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire [2:0] _GEN_57 = _T_10 ? 3'h2 : _GEN_55; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38 342:15]
  wire  _GEN_58 = _T_10 ? missPTEAF : _GEN_56; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26 341:38]
  wire  _GEN_60 = isFlush ? 1'h0 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22 340:19]
  wire  line_560_clock;
  wire  line_560_reset;
  wire  line_560_valid;
  reg  line_560_valid_reg;
  wire  _T_11 = 3'h2 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_561_clock;
  wire  line_561_reset;
  wire  line_561_valid;
  reg  line_561_valid_reg;
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_562_clock;
  wire  line_562_reset;
  wire  line_562_valid;
  reg  line_562_valid_reg;
  wire  line_563_clock;
  wire  line_563_reset;
  wire  line_563_valid;
  reg  line_563_valid_reg;
  wire  line_564_clock;
  wire  line_564_reset;
  wire  line_564_valid;
  reg  line_564_valid_reg;
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_18 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:49]
  wire  line_565_clock;
  wire  line_565_reset;
  wire  line_565_valid;
  reg  line_565_valid_reg;
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire  _T_22 = ~missflag_v | ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:28]
  wire  line_566_clock;
  wire  line_566_reset;
  wire  line_566_valid;
  reg  line_566_valid_reg;
  wire  line_567_clock;
  wire  line_567_reset;
  wire  line_567_valid;
  reg  line_567_valid_reg;
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire  line_568_clock;
  wire  line_568_reset;
  wire  line_568_valid;
  reg  line_568_valid_reg;
  wire [2:0] _GEN_62 = is_reserved ? 3'h4 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 372:21]
  wire  _GEN_63 = is_reserved | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 371:32 374:25]
  wire [2:0] _GEN_64 = ~missflag_v | ~missflag_r & missflag_w ? 3'h4 : _GEN_62; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:43]
  wire  _GEN_65 = ~missflag_v | ~missflag_r & missflag_w | _GEN_63; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 358:45]
  wire [55:0] _GEN_66 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire  line_569_clock;
  wire  line_569_reset;
  wire  line_569_valid;
  reg  line_569_valid_reg;
  wire  _T_23 = level != 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:27]
  wire  line_570_clock;
  wire  line_570_reset;
  wire  line_570_valid;
  reg  line_570_valid_reg;
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_157 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_157; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:24]
  wire  permExec = permCheck & ~_T_21 & ~permAD & ~misaligned & missflag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:75]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = 8'h40 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | 64'h40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire  _T_24 = ~permExec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 396:19]
  wire  line_571_clock;
  wire  line_571_reset;
  wire  line_571_valid;
  reg  line_571_valid_reg;
  wire  line_572_clock;
  wire  line_572_reset;
  wire  line_572_valid;
  reg  line_572_valid_reg;
  wire  _GEN_67 = ~permExec | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 396:{30,40}]
  wire  _GEN_69 = ~permExec ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 396:30 304:32 399:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_70 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_71 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire  _GEN_72 = level != 2'h0 ? _GEN_67 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 383:36]
  wire [2:0] _GEN_73 = level != 2'h0 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_74 = level != 2'h0 & _GEN_69; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_75 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_83 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_75; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_91 = isFlush ? 18'h3ffff : _GEN_83; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 302:26]
  wire [17:0] _GEN_100 = _T_12 ? _GEN_91 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_127 = 3'h2 == state ? _GEN_100 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_140 = 3'h1 == state ? 18'h3ffff : _GEN_127; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_140; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_76 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_77 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_64 : _GEN_73; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_78 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_65 : _GEN_72; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_79 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_66 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_80 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_70; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_81 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_71; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_82 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_74; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_84 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_76; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [2:0] _GEN_85 = isFlush ? 3'h0 : _GEN_77; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 353:17]
  wire  _GEN_86 = isFlush ? missIPF : _GEN_78; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 352:24]
  wire [55:0] _GEN_87 = isFlush ? raddr : _GEN_79; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 352:24]
  wire [7:0] _GEN_88 = isFlush ? 8'h0 : _GEN_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 305:32]
  wire [63:0] _GEN_89 = isFlush ? memRespStore : _GEN_81; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 301:25]
  wire  _GEN_90 = isFlush ? 1'h0 : _GEN_82; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 304:32]
  wire [17:0] _GEN_92 = isFlush ? missMaskStore : _GEN_84; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 303:26]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_93 = _T_12 ? _GEN_85 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_94 = _T_12 ? _GEN_60 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
  wire  _GEN_95 = _T_12 ? _GEN_86 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 351:33]
  wire  _GEN_99 = _T_12 & _GEN_90; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_102 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire  line_573_clock;
  wire  line_573_reset;
  wire  line_573_valid;
  reg  line_573_valid_reg;
  wire  _T_25 = 3'h3 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_574_clock;
  wire  line_574_reset;
  wire  line_574_valid;
  reg  line_574_valid_reg;
  wire  line_575_clock;
  wire  line_575_reset;
  wire  line_575_valid;
  reg  line_575_valid_reg;
  wire  line_576_clock;
  wire  line_576_reset;
  wire  line_576_valid;
  reg  line_576_valid_reg;
  wire  line_577_clock;
  wire  line_577_reset;
  wire  line_577_valid;
  reg  line_577_valid_reg;
  wire [2:0] _GEN_103 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire [2:0] _GEN_104 = isFlush ? 3'h0 : _GEN_103; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 420:22 421:15]
  wire  line_578_clock;
  wire  line_578_reset;
  wire  line_578_valid;
  reg  line_578_valid_reg;
  wire  _T_27 = 3'h4 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_579_clock;
  wire  line_579_reset;
  wire  line_579_valid;
  reg  line_579_valid_reg;
  wire  _T_29 = io_isFinish | io_flush | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:53]
  wire  line_580_clock;
  wire  line_580_reset;
  wire  line_580_valid;
  reg  line_580_valid_reg;
  wire [2:0] _GEN_105 = io_isFinish | io_flush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_106 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 428:15 318:24]
  wire  _GEN_107 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_108 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire  line_581_clock;
  wire  line_581_reset;
  wire  line_581_valid;
  reg  line_581_valid_reg;
  wire  _T_30 = 3'h5 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_582_clock;
  wire  line_582_reset;
  wire  line_582_valid;
  reg  line_582_valid_reg;
  wire [2:0] _GEN_109 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_110 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_111 = 3'h4 == state ? _GEN_105 : _GEN_109; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_112 = 3'h4 == state ? _GEN_106 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_113 = 3'h4 == state ? _GEN_107 : _GEN_110; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_114 = 3'h4 == state ? _GEN_108 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_115 = 3'h3 == state ? _GEN_104 : _GEN_111; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_116 = 3'h3 == state ? _GEN_60 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_117 = 3'h3 == state ? missIPF : _GEN_112; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_118 = 3'h3 == state ? missPTEAF : _GEN_113; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_119 = 3'h3 == state ? _GEN_42 : _GEN_114; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_139 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_99; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_139; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _io_mem_req_valid_T_3 = ~isFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:76]
  wire  _T_34 = missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:50]
  wire  _T_35 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  line_583_clock;
  wire  line_583_reset;
  wire  line_583_valid;
  reg  line_583_valid_reg;
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire  out_req_valid = io_in_valid & (hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _instrAF_T_2 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _instrAF_T_5 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _instrAF_T_6 = {_instrAF_T_5,_instrAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _instrAF_T_7 = |_instrAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  hasException = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  GEN_w1_line #(.COVER_INDEX(548)) line_548 (
    .clock(line_548_clock),
    .reset(line_548_reset),
    .valid(line_548_valid)
  );
  GEN_w1_line #(.COVER_INDEX(549)) line_549 (
    .clock(line_549_clock),
    .reset(line_549_reset),
    .valid(line_549_valid)
  );
  GEN_w1_line #(.COVER_INDEX(550)) line_550 (
    .clock(line_550_clock),
    .reset(line_550_reset),
    .valid(line_550_valid)
  );
  GEN_w1_line #(.COVER_INDEX(551)) line_551 (
    .clock(line_551_clock),
    .reset(line_551_reset),
    .valid(line_551_valid)
  );
  GEN_w1_line #(.COVER_INDEX(552)) line_552 (
    .clock(line_552_clock),
    .reset(line_552_reset),
    .valid(line_552_valid)
  );
  GEN_w1_line #(.COVER_INDEX(553)) line_553 (
    .clock(line_553_clock),
    .reset(line_553_reset),
    .valid(line_553_valid)
  );
  GEN_w1_line #(.COVER_INDEX(554)) line_554 (
    .clock(line_554_clock),
    .reset(line_554_reset),
    .valid(line_554_valid)
  );
  GEN_w1_line #(.COVER_INDEX(555)) line_555 (
    .clock(line_555_clock),
    .reset(line_555_reset),
    .valid(line_555_valid)
  );
  GEN_w1_line #(.COVER_INDEX(556)) line_556 (
    .clock(line_556_clock),
    .reset(line_556_reset),
    .valid(line_556_valid)
  );
  GEN_w1_line #(.COVER_INDEX(557)) line_557 (
    .clock(line_557_clock),
    .reset(line_557_reset),
    .valid(line_557_valid)
  );
  GEN_w1_line #(.COVER_INDEX(558)) line_558 (
    .clock(line_558_clock),
    .reset(line_558_reset),
    .valid(line_558_valid)
  );
  GEN_w1_line #(.COVER_INDEX(559)) line_559 (
    .clock(line_559_clock),
    .reset(line_559_reset),
    .valid(line_559_valid)
  );
  GEN_w1_line #(.COVER_INDEX(560)) line_560 (
    .clock(line_560_clock),
    .reset(line_560_reset),
    .valid(line_560_valid)
  );
  GEN_w1_line #(.COVER_INDEX(561)) line_561 (
    .clock(line_561_clock),
    .reset(line_561_reset),
    .valid(line_561_valid)
  );
  GEN_w1_line #(.COVER_INDEX(562)) line_562 (
    .clock(line_562_clock),
    .reset(line_562_reset),
    .valid(line_562_valid)
  );
  GEN_w1_line #(.COVER_INDEX(563)) line_563 (
    .clock(line_563_clock),
    .reset(line_563_reset),
    .valid(line_563_valid)
  );
  GEN_w1_line #(.COVER_INDEX(564)) line_564 (
    .clock(line_564_clock),
    .reset(line_564_reset),
    .valid(line_564_valid)
  );
  GEN_w1_line #(.COVER_INDEX(565)) line_565 (
    .clock(line_565_clock),
    .reset(line_565_reset),
    .valid(line_565_valid)
  );
  GEN_w1_line #(.COVER_INDEX(566)) line_566 (
    .clock(line_566_clock),
    .reset(line_566_reset),
    .valid(line_566_valid)
  );
  GEN_w1_line #(.COVER_INDEX(567)) line_567 (
    .clock(line_567_clock),
    .reset(line_567_reset),
    .valid(line_567_valid)
  );
  GEN_w1_line #(.COVER_INDEX(568)) line_568 (
    .clock(line_568_clock),
    .reset(line_568_reset),
    .valid(line_568_valid)
  );
  GEN_w1_line #(.COVER_INDEX(569)) line_569 (
    .clock(line_569_clock),
    .reset(line_569_reset),
    .valid(line_569_valid)
  );
  GEN_w1_line #(.COVER_INDEX(570)) line_570 (
    .clock(line_570_clock),
    .reset(line_570_reset),
    .valid(line_570_valid)
  );
  GEN_w1_line #(.COVER_INDEX(571)) line_571 (
    .clock(line_571_clock),
    .reset(line_571_reset),
    .valid(line_571_valid)
  );
  GEN_w1_line #(.COVER_INDEX(572)) line_572 (
    .clock(line_572_clock),
    .reset(line_572_reset),
    .valid(line_572_valid)
  );
  GEN_w1_line #(.COVER_INDEX(573)) line_573 (
    .clock(line_573_clock),
    .reset(line_573_reset),
    .valid(line_573_valid)
  );
  GEN_w1_line #(.COVER_INDEX(574)) line_574 (
    .clock(line_574_clock),
    .reset(line_574_reset),
    .valid(line_574_valid)
  );
  GEN_w1_line #(.COVER_INDEX(575)) line_575 (
    .clock(line_575_clock),
    .reset(line_575_reset),
    .valid(line_575_valid)
  );
  GEN_w1_line #(.COVER_INDEX(576)) line_576 (
    .clock(line_576_clock),
    .reset(line_576_reset),
    .valid(line_576_valid)
  );
  GEN_w1_line #(.COVER_INDEX(577)) line_577 (
    .clock(line_577_clock),
    .reset(line_577_reset),
    .valid(line_577_valid)
  );
  GEN_w1_line #(.COVER_INDEX(578)) line_578 (
    .clock(line_578_clock),
    .reset(line_578_reset),
    .valid(line_578_valid)
  );
  GEN_w1_line #(.COVER_INDEX(579)) line_579 (
    .clock(line_579_clock),
    .reset(line_579_reset),
    .valid(line_579_valid)
  );
  GEN_w1_line #(.COVER_INDEX(580)) line_580 (
    .clock(line_580_clock),
    .reset(line_580_reset),
    .valid(line_580_valid)
  );
  GEN_w1_line #(.COVER_INDEX(581)) line_581 (
    .clock(line_581_clock),
    .reset(line_581_reset),
    .valid(line_581_valid)
  );
  GEN_w1_line #(.COVER_INDEX(582)) line_582 (
    .clock(line_582_clock),
    .reset(line_582_reset),
    .valid(line_582_valid)
  );
  GEN_w1_line #(.COVER_INDEX(583)) line_583 (
    .clock(line_583_clock),
    .reset(line_583_reset),
    .valid(line_583_valid)
  );
  assign line_548_clock = clock;
  assign line_548_reset = reset;
  assign line_548_valid = _alreadyOutFire_T ^ line_548_valid_reg;
  assign line_549_clock = clock;
  assign line_549_reset = reset;
  assign line_549_valid = _T_1 ^ line_549_valid_reg;
  assign line_550_clock = clock;
  assign line_550_reset = reset;
  assign line_550_valid = _T_3 ^ line_550_valid_reg;
  assign line_551_clock = clock;
  assign line_551_reset = reset;
  assign line_551_valid = _T_4 ^ line_551_valid_reg;
  assign line_552_clock = clock;
  assign line_552_reset = reset;
  assign line_552_valid = _T_8 ^ line_552_valid_reg;
  assign line_553_clock = clock;
  assign line_553_reset = reset;
  assign line_553_valid = _T_4 ^ line_553_valid_reg;
  assign line_554_clock = clock;
  assign line_554_reset = reset;
  assign line_554_valid = _T_9 ^ line_554_valid_reg;
  assign line_555_clock = clock;
  assign line_555_reset = reset;
  assign line_555_valid = isFlush ^ line_555_valid_reg;
  assign line_556_clock = clock;
  assign line_556_reset = reset;
  assign line_556_valid = isFlush ^ line_556_valid_reg;
  assign line_557_clock = clock;
  assign line_557_reset = reset;
  assign line_557_valid = _T_10 ^ line_557_valid_reg;
  assign line_558_clock = clock;
  assign line_558_reset = reset;
  assign line_558_valid = _T_10 ^ line_558_valid_reg;
  assign line_559_clock = clock;
  assign line_559_reset = reset;
  assign line_559_valid = raddrCancel ^ line_559_valid_reg;
  assign line_560_clock = clock;
  assign line_560_reset = reset;
  assign line_560_valid = _T_9 ^ line_560_valid_reg;
  assign line_561_clock = clock;
  assign line_561_reset = reset;
  assign line_561_valid = _T_11 ^ line_561_valid_reg;
  assign line_562_clock = clock;
  assign line_562_reset = reset;
  assign line_562_valid = _T_12 ^ line_562_valid_reg;
  assign line_563_clock = clock;
  assign line_563_reset = reset;
  assign line_563_valid = isFlush ^ line_563_valid_reg;
  assign line_564_clock = clock;
  assign line_564_reset = reset;
  assign line_564_valid = isFlush ^ line_564_valid_reg;
  assign line_565_clock = clock;
  assign line_565_reset = reset;
  assign line_565_valid = _T_18 ^ line_565_valid_reg;
  assign line_566_clock = clock;
  assign line_566_reset = reset;
  assign line_566_valid = _T_22 ^ line_566_valid_reg;
  assign line_567_clock = clock;
  assign line_567_reset = reset;
  assign line_567_valid = _T_22 ^ line_567_valid_reg;
  assign line_568_clock = clock;
  assign line_568_reset = reset;
  assign line_568_valid = is_reserved ^ line_568_valid_reg;
  assign line_569_clock = clock;
  assign line_569_reset = reset;
  assign line_569_valid = _T_18 ^ line_569_valid_reg;
  assign line_570_clock = clock;
  assign line_570_reset = reset;
  assign line_570_valid = _T_23 ^ line_570_valid_reg;
  assign line_571_clock = clock;
  assign line_571_reset = reset;
  assign line_571_valid = _T_24 ^ line_571_valid_reg;
  assign line_572_clock = clock;
  assign line_572_reset = reset;
  assign line_572_valid = _T_24 ^ line_572_valid_reg;
  assign line_573_clock = clock;
  assign line_573_reset = reset;
  assign line_573_valid = _T_11 ^ line_573_valid_reg;
  assign line_574_clock = clock;
  assign line_574_reset = reset;
  assign line_574_valid = _T_25 ^ line_574_valid_reg;
  assign line_575_clock = clock;
  assign line_575_reset = reset;
  assign line_575_valid = isFlush ^ line_575_valid_reg;
  assign line_576_clock = clock;
  assign line_576_reset = reset;
  assign line_576_valid = isFlush ^ line_576_valid_reg;
  assign line_577_clock = clock;
  assign line_577_reset = reset;
  assign line_577_valid = _T_10 ^ line_577_valid_reg;
  assign line_578_clock = clock;
  assign line_578_reset = reset;
  assign line_578_valid = _T_25 ^ line_578_valid_reg;
  assign line_579_clock = clock;
  assign line_579_reset = reset;
  assign line_579_valid = _T_27 ^ line_579_valid_reg;
  assign line_580_clock = clock;
  assign line_580_reset = reset;
  assign line_580_valid = _T_29 ^ line_580_valid_reg;
  assign line_581_clock = clock;
  assign line_581_reset = reset;
  assign line_581_valid = _T_27 ^ line_581_valid_reg;
  assign line_582_clock = clock;
  assign line_582_reset = reset;
  assign line_582_valid = _T_30 ^ line_582_valid_reg;
  assign line_583_clock = clock;
  assign line_583_reset = reset;
  assign line_583_valid = blockRefill ^ line_583_valid_reg;
  assign io_in_ready = io_out_ready & _T_35 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:75]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_user = io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 500:16]
  assign io_iaf = out_req_valid & (~_instrAF_T_7 | missPTEAF); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 486:30]
  assign io_isFinish = _alreadyOutFire_T | hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:32]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 339:15]
      end else begin
        state <= _GEN_57;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_93;
    end else begin
      state <= _GEN_115;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_102;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_89;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_92;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_87;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_42;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_42;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_42;
    end else begin
      alreadyOutFire <= _GEN_119;
    end
    line_548_valid_reg <= _alreadyOutFire_T;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 332:19]
      end else begin
        needFlush <= _GEN_44;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 340:19]
      end else begin
        needFlush <= _GEN_44;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      needFlush <= _GEN_94;
    end else begin
      needFlush <= _GEN_116;
    end
    line_549_valid_reg <= _T_1;
    line_550_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
      missIPF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          missIPF <= _GEN_95;
        end else begin
          missIPF <= _GEN_117;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(isFlush)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
          missPTEAF <= _GEN_58;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_118;
      end
    end
    line_551_valid_reg <= _T_4;
    line_552_valid_reg <= _T_8;
    line_553_valid_reg <= _T_4;
    line_554_valid_reg <= _T_9;
    line_555_valid_reg <= isFlush;
    line_556_valid_reg <= isFlush;
    line_557_valid_reg <= _T_10;
    line_558_valid_reg <= _T_10;
    line_559_valid_reg <= raddrCancel;
    line_560_valid_reg <= _T_9;
    line_561_valid_reg <= _T_11;
    line_562_valid_reg <= _T_12;
    line_563_valid_reg <= isFlush;
    line_564_valid_reg <= isFlush;
    line_565_valid_reg <= _T_18;
    line_566_valid_reg <= _T_22;
    line_567_valid_reg <= _T_22;
    line_568_valid_reg <= is_reserved;
    line_569_valid_reg <= _T_18;
    line_570_valid_reg <= _T_23;
    line_571_valid_reg <= _T_24;
    line_572_valid_reg <= _T_24;
    line_573_valid_reg <= _T_11;
    line_574_valid_reg <= _T_25;
    line_575_valid_reg <= isFlush;
    line_576_valid_reg <= isFlush;
    line_577_valid_reg <= _T_10;
    line_578_valid_reg <= _T_25;
    line_579_valid_reg <= _T_27;
    line_580_valid_reg <= _T_29;
    line_581_valid_reg <= _T_27;
    line_582_valid_reg <= _T_30;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else begin
      REG <= missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_91;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_88;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= _T_34 & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
    line_583_valid_reg <= blockRefill;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  memRespStore = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  missMaskStore = _RAND_4[17:0];
  _RAND_5 = {2{`RANDOM}};
  raddr = _RAND_5[55:0];
  _RAND_6 = {1{`RANDOM}};
  alreadyOutFire = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_548_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_549_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_550_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  missIPF = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  missPTEAF = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_551_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_552_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_553_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_554_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_555_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_556_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_557_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_558_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_559_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_560_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_561_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_562_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_563_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_564_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_565_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_566_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_567_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_568_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_569_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_570_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_571_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_572_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_573_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_574_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_575_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_576_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_577_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_578_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_579_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_580_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_581_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_582_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_2 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  REG_3 = _RAND_47[26:0];
  _RAND_48 = {1{`RANDOM}};
  REG_4 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  REG_5 = _RAND_49[17:0];
  _RAND_50 = {1{`RANDOM}};
  REG_6 = _RAND_50[7:0];
  _RAND_51 = {2{`RANDOM}};
  REG_7 = _RAND_51[43:0];
  _RAND_52 = {2{`RANDOM}};
  REG_8 = _RAND_52[55:0];
  _RAND_53 = {1{`RANDOM}};
  blockRefill = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_583_valid_reg = _RAND_54[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_alreadyOutFire_T) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_3) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _T_8) begin
      cover(1'h1);
    end
    //
    if (~_T_4) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & isFlush) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & _io_mem_req_valid_T_3) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & _io_mem_req_valid_T_3 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & _io_mem_req_valid_T_3 & ~_T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & _io_mem_req_valid_T_3 & ~_T_10 & raddrCancel) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & isFlush) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18 & _T_22) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18 & ~_T_22) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & _T_18 & ~_T_22 & is_reserved) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & ~_T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & ~_T_18 & _T_23) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & ~_T_18 & _T_23 & _T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _io_mem_req_valid_T_3 & ~_T_18 & _T_23 & ~_T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_25) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_25 & isFlush) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_25 & _io_mem_req_valid_T_3) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_25 & _io_mem_req_valid_T_3 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_25) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_25 & _T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_25 & _T_27 & _T_29) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_25 & ~_T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_25 & ~_T_27 & _T_30) begin
      cover(1'h1);
    end
    //
    if (blockRefill) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLBEmpty(
  input   clock,
  input   reset
);
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  line_584_clock;
  wire  line_584_reset;
  wire  line_584_valid;
  reg  line_584_valid_reg;
  wire  line_585_clock;
  wire  line_585_reset;
  wire  line_585_valid;
  reg  line_585_valid_reg;
  wire  _GEN_8 = resetState ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire  wen = resetState | io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:16]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  wire  line_586_clock;
  wire  line_586_reset;
  wire  line_586_valid;
  reg  line_586_valid_reg;
  wire  line_587_clock;
  wire  line_587_reset;
  wire  line_587_valid;
  reg  line_587_valid_reg;
  wire  line_588_clock;
  wire  line_588_reset;
  wire  line_588_valid;
  reg  line_588_valid_reg;
  wire  line_589_clock;
  wire  line_589_reset;
  wire  line_589_valid;
  reg  line_589_valid_reg;
  wire  line_590_clock;
  wire  line_590_reset;
  wire  line_590_valid;
  reg  line_590_valid_reg;
  GEN_w1_line #(.COVER_INDEX(584)) line_584 (
    .clock(line_584_clock),
    .reset(line_584_reset),
    .valid(line_584_valid)
  );
  GEN_w1_line #(.COVER_INDEX(585)) line_585 (
    .clock(line_585_clock),
    .reset(line_585_reset),
    .valid(line_585_valid)
  );
  GEN_w1_line #(.COVER_INDEX(586)) line_586 (
    .clock(line_586_clock),
    .reset(line_586_reset),
    .valid(line_586_valid)
  );
  GEN_w1_line #(.COVER_INDEX(587)) line_587 (
    .clock(line_587_clock),
    .reset(line_587_reset),
    .valid(line_587_valid)
  );
  GEN_w1_line #(.COVER_INDEX(588)) line_588 (
    .clock(line_588_clock),
    .reset(line_588_reset),
    .valid(line_588_valid)
  );
  GEN_w1_line #(.COVER_INDEX(589)) line_589 (
    .clock(line_589_clock),
    .reset(line_589_reset),
    .valid(line_589_valid)
  );
  GEN_w1_line #(.COVER_INDEX(590)) line_590 (
    .clock(line_590_clock),
    .reset(line_590_reset),
    .valid(line_590_valid)
  );
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign line_584_clock = clock;
  assign line_584_reset = reset;
  assign line_584_valid = resetState ^ line_584_valid_reg;
  assign line_585_clock = clock;
  assign line_585_reset = reset;
  assign line_585_valid = resetState ^ line_585_valid_reg;
  assign line_586_clock = clock;
  assign line_586_reset = reset;
  assign line_586_valid = wen ^ line_586_valid_reg;
  assign line_587_clock = clock;
  assign line_587_reset = reset;
  assign line_587_valid = waymask[0] ^ line_587_valid_reg;
  assign line_588_clock = clock;
  assign line_588_reset = reset;
  assign line_588_valid = waymask[1] ^ line_588_valid_reg;
  assign line_589_clock = clock;
  assign line_589_reset = reset;
  assign line_589_valid = waymask[2] ^ line_589_valid_reg;
  assign line_590_clock = clock;
  assign line_590_reset = reset;
  assign line_590_valid = waymask[3] ^ line_590_valid_reg;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
    line_584_valid_reg <= resetState;
    line_585_valid_reg <= resetState;
    line_586_valid_reg <= wen;
    line_587_valid_reg <= waymask[0];
    line_588_valid_reg <= waymask[1];
    line_589_valid_reg <= waymask[2];
    line_590_valid_reg <= waymask[3];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_584_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_585_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_586_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_587_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_588_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_589_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_590_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (resetState) begin
      cover(1'h1);
    end
    //
    if (resetState) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[0]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[1]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[2]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[3]) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_out_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_out_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbEmpty_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  wire  line_591_clock;
  wire  line_591_reset;
  wire  line_591_valid;
  reg  line_591_valid_reg;
  wire  _reqIsLegalInstr_T_2 = io_in_req_bits_addr >= 39'h40000000 & io_in_req_bits_addr < 39'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _reqIsLegalInstr_T_5 = io_in_req_bits_addr >= 39'h80000000 & io_in_req_bits_addr < 39'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _reqIsLegalInstr_T_6 = {_reqIsLegalInstr_T_5,_reqIsLegalInstr_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _reqIsLegalInstr_T_7 = |_reqIsLegalInstr_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  reqIsLegalInstr = vmEnable | _reqIsLegalInstr_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 119:34]
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
  wire  _lastReqAddr_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _lastReqAddr_T_1 = ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:70]
  wire  _lastReqAddr_T_2 = _lastReqAddr_T & ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:67]
  reg [38:0] lastReqAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
  wire  line_592_clock;
  wire  line_592_reset;
  wire  line_592_valid;
  reg  line_592_valid_reg;
  wire  line_593_clock;
  wire  line_593_reset;
  wire  line_593_valid;
  reg  line_593_valid_reg;
  wire  line_594_clock;
  wire  line_594_reset;
  wire  line_594_valid;
  reg  line_594_valid_reg;
  wire  line_595_clock;
  wire  line_595_reset;
  wire  line_595_valid;
  reg  line_595_valid_reg;
  wire  line_596_clock;
  wire  line_596_reset;
  wire  line_596_valid;
  reg  line_596_valid_reg;
  wire  _T_1 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_4 = _T_1 & io_in_resp_bits_user[38:0] == lastReqAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 127:33]
  wire  line_597_clock;
  wire  line_597_reset;
  wire  line_597_valid;
  reg  line_597_valid_reg;
  wire  _GEN_26 = _T_1 & io_in_resp_bits_user[38:0] == lastReqAddr ? 1'h0 : hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 127:96 128:19 120:28]
  wire  _GEN_27 = _lastReqAddr_T | _GEN_26; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 125:33 126:19]
  reg  hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
  wire  _T_6 = _T_1 | io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 132:25]
  wire  line_598_clock;
  wire  line_598_reset;
  wire  line_598_valid;
  reg  line_598_valid_reg;
  wire  line_599_clock;
  wire  line_599_reset;
  wire  line_599_valid;
  reg  line_599_valid_reg;
  wire  line_600_clock;
  wire  line_600_reset;
  wire  line_600_valid;
  reg  line_600_valid_reg;
  wire  _hasIllegalInflight_T = ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:27]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  line_601_clock;
  wire  line_601_reset;
  wire  line_601_valid;
  reg  line_601_valid_reg;
  wire  _GEN_31 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _T_11 = mdUpdate & vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:37]
  wire  line_602_clock;
  wire  line_602_reset;
  wire  line_602_valid;
  reg  line_602_valid_reg;
  wire  _GEN_32 = mdUpdate & vmEnable | _GEN_31; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  wire  line_603_clock;
  wire  line_603_reset;
  wire  line_603_valid;
  reg  line_603_valid_reg;
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [86:0] tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  line_604_clock;
  wire  line_604_reset;
  wire  line_604_valid;
  reg  line_604_valid_reg;
  wire  _T_12 = ~vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:8]
  wire  line_605_clock;
  wire  line_605_reset;
  wire  line_605_valid;
  reg  line_605_valid_reg;
  wire  _T_14 = io_in_req_valid & _hasIllegalInflight_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 158:29]
  wire  line_606_clock;
  wire  line_606_reset;
  wire  line_606_valid;
  reg  line_606_valid_reg;
  wire  _GEN_40 = io_in_req_valid & _hasIllegalInflight_T ? ~hasInflight : io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:23 158:50 159:25]
  wire  line_607_clock;
  wire  line_607_reset;
  wire  line_607_valid;
  reg  line_607_valid_reg;
  wire  _GEN_41 = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 170:23]
  wire  _GEN_42 = ~vmEnable ? io_in_req_valid & reqIsLegalInstr : tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 156:24 170:23]
  wire  _T_16 = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:46]
  wire  line_608_clock;
  wire  line_608_reset;
  wire  line_608_valid;
  reg  line_608_valid_reg;
  wire  _T_20 = hasIllegalInflight & io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:30]
  wire  line_609_clock;
  wire  line_609_reset;
  wire  line_609_valid;
  reg  line_609_valid_reg;
  reg [86:0] userBits; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
  wire  line_610_clock;
  wire  line_610_reset;
  wire  line_610_valid;
  reg  line_610_valid_reg;
  EmbeddedTLBExec tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_ipf(tlbExec_io_ipf),
    .io_iaf(tlbExec_io_iaf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBEmpty tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
    .clock(tlbEmpty_clock),
    .reset(tlbEmpty_reset)
  );
  EmbeddedTLBMD mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  GEN_w1_line #(.COVER_INDEX(591)) line_591 (
    .clock(line_591_clock),
    .reset(line_591_reset),
    .valid(line_591_valid)
  );
  GEN_w1_line #(.COVER_INDEX(592)) line_592 (
    .clock(line_592_clock),
    .reset(line_592_reset),
    .valid(line_592_valid)
  );
  GEN_w1_line #(.COVER_INDEX(593)) line_593 (
    .clock(line_593_clock),
    .reset(line_593_reset),
    .valid(line_593_valid)
  );
  GEN_w1_line #(.COVER_INDEX(594)) line_594 (
    .clock(line_594_clock),
    .reset(line_594_reset),
    .valid(line_594_valid)
  );
  GEN_w1_line #(.COVER_INDEX(595)) line_595 (
    .clock(line_595_clock),
    .reset(line_595_reset),
    .valid(line_595_valid)
  );
  GEN_w1_line #(.COVER_INDEX(596)) line_596 (
    .clock(line_596_clock),
    .reset(line_596_reset),
    .valid(line_596_valid)
  );
  GEN_w1_line #(.COVER_INDEX(597)) line_597 (
    .clock(line_597_clock),
    .reset(line_597_reset),
    .valid(line_597_valid)
  );
  GEN_w1_line #(.COVER_INDEX(598)) line_598 (
    .clock(line_598_clock),
    .reset(line_598_reset),
    .valid(line_598_valid)
  );
  GEN_w1_line #(.COVER_INDEX(599)) line_599 (
    .clock(line_599_clock),
    .reset(line_599_reset),
    .valid(line_599_valid)
  );
  GEN_w1_line #(.COVER_INDEX(600)) line_600 (
    .clock(line_600_clock),
    .reset(line_600_reset),
    .valid(line_600_valid)
  );
  GEN_w1_line #(.COVER_INDEX(601)) line_601 (
    .clock(line_601_clock),
    .reset(line_601_reset),
    .valid(line_601_valid)
  );
  GEN_w1_line #(.COVER_INDEX(602)) line_602 (
    .clock(line_602_clock),
    .reset(line_602_reset),
    .valid(line_602_valid)
  );
  GEN_w1_line #(.COVER_INDEX(603)) line_603 (
    .clock(line_603_clock),
    .reset(line_603_reset),
    .valid(line_603_valid)
  );
  GEN_w1_line #(.COVER_INDEX(604)) line_604 (
    .clock(line_604_clock),
    .reset(line_604_reset),
    .valid(line_604_valid)
  );
  GEN_w1_line #(.COVER_INDEX(605)) line_605 (
    .clock(line_605_clock),
    .reset(line_605_reset),
    .valid(line_605_valid)
  );
  GEN_w1_line #(.COVER_INDEX(606)) line_606 (
    .clock(line_606_clock),
    .reset(line_606_reset),
    .valid(line_606_valid)
  );
  GEN_w1_line #(.COVER_INDEX(607)) line_607 (
    .clock(line_607_clock),
    .reset(line_607_reset),
    .valid(line_607_valid)
  );
  GEN_w1_line #(.COVER_INDEX(608)) line_608 (
    .clock(line_608_clock),
    .reset(line_608_reset),
    .valid(line_608_valid)
  );
  GEN_w1_line #(.COVER_INDEX(609)) line_609 (
    .clock(line_609_clock),
    .reset(line_609_reset),
    .valid(line_609_valid)
  );
  GEN_w1_line #(.COVER_INDEX(610)) line_610 (
    .clock(line_610_clock),
    .reset(line_610_reset),
    .valid(line_610_valid)
  );
  assign line_591_clock = clock;
  assign line_591_reset = reset;
  assign line_591_valid = mdUpdate ^ line_591_valid_reg;
  assign line_592_clock = clock;
  assign line_592_reset = reset;
  assign line_592_valid = _lastReqAddr_T_2 ^ line_592_valid_reg;
  assign line_593_clock = clock;
  assign line_593_reset = reset;
  assign line_593_valid = io_flush ^ line_593_valid_reg;
  assign line_594_clock = clock;
  assign line_594_reset = reset;
  assign line_594_valid = io_flush ^ line_594_valid_reg;
  assign line_595_clock = clock;
  assign line_595_reset = reset;
  assign line_595_valid = _lastReqAddr_T ^ line_595_valid_reg;
  assign line_596_clock = clock;
  assign line_596_reset = reset;
  assign line_596_valid = _lastReqAddr_T ^ line_596_valid_reg;
  assign line_597_clock = clock;
  assign line_597_reset = reset;
  assign line_597_valid = _T_4 ^ line_597_valid_reg;
  assign line_598_clock = clock;
  assign line_598_reset = reset;
  assign line_598_valid = _T_6 ^ line_598_valid_reg;
  assign line_599_clock = clock;
  assign line_599_reset = reset;
  assign line_599_valid = _T_6 ^ line_599_valid_reg;
  assign line_600_clock = clock;
  assign line_600_reset = reset;
  assign line_600_valid = _lastReqAddr_T_2 ^ line_600_valid_reg;
  assign line_601_clock = clock;
  assign line_601_reset = reset;
  assign line_601_valid = tlbExec_io_isFinish ^ line_601_valid_reg;
  assign line_602_clock = clock;
  assign line_602_reset = reset;
  assign line_602_valid = _T_11 ^ line_602_valid_reg;
  assign line_603_clock = clock;
  assign line_603_reset = reset;
  assign line_603_valid = io_flush ^ line_603_valid_reg;
  assign line_604_clock = clock;
  assign line_604_reset = reset;
  assign line_604_valid = mdUpdate ^ line_604_valid_reg;
  assign line_605_clock = clock;
  assign line_605_reset = reset;
  assign line_605_valid = _T_12 ^ line_605_valid_reg;
  assign line_606_clock = clock;
  assign line_606_reset = reset;
  assign line_606_valid = _T_14 ^ line_606_valid_reg;
  assign line_607_clock = clock;
  assign line_607_reset = reset;
  assign line_607_valid = _T_12 ^ line_607_valid_reg;
  assign line_608_clock = clock;
  assign line_608_reset = reset;
  assign line_608_valid = _T_16 ^ line_608_valid_reg;
  assign line_609_clock = clock;
  assign line_609_reset = reset;
  assign line_609_valid = _T_20 ^ line_609_valid_reg;
  assign line_610_clock = clock;
  assign line_610_reset = reset;
  assign line_610_valid = _lastReqAddr_T_2 ^ line_610_valid_reg;
  assign io_in_req_ready = ~vmEnable ? _GEN_40 : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19]
  assign io_in_resp_valid = hasIllegalInflight & io_iaf | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 202:24]
  assign io_in_resp_bits_rdata = hasIllegalInflight & io_iaf ? 64'h0 : io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 203:29]
  assign io_in_resp_bits_user = hasIllegalInflight & io_iaf ? userBits : io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 206:34]
  assign io_out_req_valid = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 191:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 170:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 167:32 170:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_iaf = vmEnable ? tlbExec_io_iaf : hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 212:16]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_user = tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_41; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 190:28]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_flush = io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:20]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbEmpty_clock = clock;
  assign tlbEmpty_reset = reset;
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    line_591_valid_reg <= mdUpdate;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 123:21]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 124:19]
    end else begin
      hasInflight <= _GEN_27;
    end
    if (_lastReqAddr_T & ~io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
      lastReqAddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    line_592_valid_reg <= _lastReqAddr_T_2;
    line_593_valid_reg <= io_flush;
    line_594_valid_reg <= io_flush;
    line_595_valid_reg <= _lastReqAddr_T;
    line_596_valid_reg <= _lastReqAddr_T;
    line_597_valid_reg <= _T_4;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
    end else if (_T_1 | io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 132:38]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 133:24]
    end else if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 134:44]
      hasIllegalInflight <= ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:24]
    end
    line_598_valid_reg <= _T_6;
    line_599_valid_reg <= _T_6;
    line_600_valid_reg <= _lastReqAddr_T_2;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:20]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:28]
    end else begin
      valid <= _GEN_32;
    end
    line_601_valid_reg <= tlbExec_io_isFinish;
    line_602_valid_reg <= _T_11;
    line_603_valid_reg <= io_flush;
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_user <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    line_604_valid_reg <= mdUpdate;
    line_605_valid_reg <= _T_12;
    line_606_valid_reg <= _T_14;
    line_607_valid_reg <= _T_12;
    line_608_valid_reg <= _T_16;
    line_609_valid_reg <= _T_20;
    if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
      userBits <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    line_610_valid_reg <= _lastReqAddr_T_2;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  line_591_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  hasInflight = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  lastReqAddr = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  line_592_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_593_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_594_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_595_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_596_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_597_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  hasIllegalInflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_598_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_599_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_600_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_601_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_602_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_603_valid_reg = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_21[38:0];
  _RAND_22 = {3{`RANDOM}};
  tlbExec_io_in_bits_r_user = _RAND_22[86:0];
  _RAND_23 = {1{`RANDOM}};
  line_604_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_605_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_606_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_607_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_608_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_609_valid_reg = _RAND_28[0:0];
  _RAND_29 = {3{`RANDOM}};
  userBits = _RAND_29[86:0];
  _RAND_30 = {1{`RANDOM}};
  line_610_valid_reg = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (mdUpdate) begin
      cover(1'h1);
    end
    //
    if (_lastReqAddr_T_2) begin
      cover(1'h1);
    end
    //
    if (io_flush) begin
      cover(1'h1);
    end
    //
    if (~io_flush) begin
      cover(1'h1);
    end
    //
    if (_lastReqAddr_T_1 & _lastReqAddr_T) begin
      cover(1'h1);
    end
    //
    if (_lastReqAddr_T_1 & ~_lastReqAddr_T) begin
      cover(1'h1);
    end
    //
    if (_lastReqAddr_T_1 & ~_lastReqAddr_T & _T_4) begin
      cover(1'h1);
    end
    //
    if (_T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_6 & _lastReqAddr_T_2) begin
      cover(1'h1);
    end
    //
    if (tlbExec_io_isFinish) begin
      cover(1'h1);
    end
    //
    if (_T_11) begin
      cover(1'h1);
    end
    //
    if (io_flush) begin
      cover(1'h1);
    end
    //
    if (mdUpdate) begin
      cover(1'h1);
    end
    //
    if (_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_12 & _T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_16) begin
      cover(1'h1);
    end
    //
    if (_T_20) begin
      cover(1'h1);
    end
    //
    if (_T_20 & _lastReqAddr_T_2) begin
      cover(1'h1);
    end
  end
endmodule
module PTERequestFilter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_u // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  isLegal = |(io_in_req_bits_addr >= 32'h80000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasInflight_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _hasInflight_T_2 = _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:33]
  wire  line_611_clock;
  wire  line_611_reset;
  wire  line_611_valid;
  reg  line_611_valid_reg;
  wire  _T_1 = ~io_out_resp_valid & hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:28]
  wire  line_612_clock;
  wire  line_612_reset;
  wire  line_612_valid;
  reg  line_612_valid_reg;
  wire [7:0] _io_in_resp_bits_rdata_T = {3'h7,io_u,4'hf}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 570:33]
  GEN_w1_line #(.COVER_INDEX(611)) line_611 (
    .clock(line_611_clock),
    .reset(line_611_reset),
    .valid(line_611_valid)
  );
  GEN_w1_line #(.COVER_INDEX(612)) line_612 (
    .clock(line_612_clock),
    .reset(line_612_reset),
    .valid(line_612_valid)
  );
  assign line_611_clock = clock;
  assign line_611_reset = reset;
  assign line_611_valid = _hasInflight_T_2 ^ line_611_valid_reg;
  assign line_612_clock = clock;
  assign line_612_reset = reset;
  assign line_612_valid = _T_1 ^ line_612_valid_reg;
  assign io_in_req_ready = isLegal ? io_out_req_ready : ~hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 562:25]
  assign io_in_resp_valid = ~io_out_resp_valid & hasInflight | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 567:22]
  assign io_in_resp_bits_rdata = ~io_out_resp_valid & hasInflight ? {{56'd0}, _io_in_resp_bits_rdata_T} :
    io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 570:27]
  assign io_out_req_valid = io_in_req_valid & isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 561:39]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end else if (~io_out_resp_valid & hasInflight) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:44]
      hasInflight <= 1'h0;
    end else begin
      hasInflight <= _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:15]
    end
    line_611_valid_reg <= _hasInflight_T_2;
    line_612_valid_reg <= _T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasInflight = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_611_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_612_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_hasInflight_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module Cache_fake(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [95:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  line_613_clock;
  wire  line_613_reset;
  wire  line_613_valid;
  reg  line_613_valid_reg;
  reg  needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  _T_2 = io_flush[0] & state != 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 567:21]
  wire  line_614_clock;
  wire  line_614_reset;
  wire  line_614_valid;
  reg  line_614_valid_reg;
  wire  _GEN_32 = io_flush[0] & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26 567:{44,56}]
  wire  _T_4 = state == 3'h0 & needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 568:26]
  wire  line_615_clock;
  wire  line_615_reset;
  wire  line_615_valid;
  reg  line_615_valid_reg;
  wire  _alreadyOutFire_T = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  line_616_clock;
  wire  line_616_reset;
  wire  line_616_valid;
  reg  line_616_valid_reg;
  wire  _GEN_34 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_5 = 3'h0 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_617_clock;
  wire  line_617_reset;
  wire  line_617_valid;
  reg  line_617_valid_reg;
  wire  _T_9 = _ismmioRec_T & ~io_flush[0]; // @[src/main/scala/nutcore/mem/Cache.scala 575:30]
  wire  line_618_clock;
  wire  line_618_reset;
  wire  line_618_valid;
  reg  line_618_valid_reg;
  wire  line_619_clock;
  wire  line_619_reset;
  wire  line_619_valid;
  reg  line_619_valid_reg;
  wire  _T_10 = 3'h1 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_620_clock;
  wire  line_620_reset;
  wire  line_620_valid;
  reg  line_620_valid_reg;
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_621_clock;
  wire  line_621_reset;
  wire  line_621_valid;
  reg  line_621_valid_reg;
  wire  line_622_clock;
  wire  line_622_reset;
  wire  line_622_valid;
  reg  line_622_valid_reg;
  wire  _T_12 = 3'h2 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_623_clock;
  wire  line_623_reset;
  wire  line_623_valid;
  reg  line_623_valid_reg;
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_624_clock;
  wire  line_624_reset;
  wire  line_624_valid;
  reg  line_624_valid_reg;
  wire [2:0] _GEN_37 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  line_625_clock;
  wire  line_625_reset;
  wire  line_625_valid;
  reg  line_625_valid_reg;
  wire  _T_14 = 3'h3 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_626_clock;
  wire  line_626_reset;
  wire  line_626_valid;
  reg  line_626_valid_reg;
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_627_clock;
  wire  line_627_reset;
  wire  line_627_valid;
  reg  line_627_valid_reg;
  wire [2:0] _GEN_38 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  line_628_clock;
  wire  line_628_reset;
  wire  line_628_valid;
  reg  line_628_valid_reg;
  wire  _T_16 = 3'h4 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_629_clock;
  wire  line_629_reset;
  wire  line_629_valid;
  reg  line_629_valid_reg;
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_18 = _T_17 | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 587:33]
  wire  line_630_clock;
  wire  line_630_reset;
  wire  line_630_valid;
  reg  line_630_valid_reg;
  wire [2:0] _GEN_39 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire  line_631_clock;
  wire  line_631_reset;
  wire  line_631_valid;
  reg  line_631_valid_reg;
  wire  _T_19 = 3'h5 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_632_clock;
  wire  line_632_reset;
  wire  line_632_valid;
  reg  line_632_valid_reg;
  wire  _T_22 = _alreadyOutFire_T | needFlush | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 590:44]
  wire  line_633_clock;
  wire  line_633_reset;
  wire  line_633_valid;
  reg  line_633_valid_reg;
  wire [2:0] _GEN_40 = _alreadyOutFire_T | needFlush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_41 = 3'h5 == state ? _GEN_40 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_42 = 3'h4 == state ? _GEN_39 : _GEN_41; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_43 = 3'h3 == state ? _GEN_38 : _GEN_42; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire  line_634_clock;
  wire  line_634_reset;
  wire  line_634_valid;
  reg  line_634_valid_reg;
  wire  line_635_clock;
  wire  line_635_reset;
  wire  line_635_valid;
  reg  line_635_valid_reg;
  wire  line_636_clock;
  wire  line_636_reset;
  wire  line_636_valid;
  reg  line_636_valid_reg;
  wire  line_637_clock;
  wire  line_637_reset;
  wire  line_637_valid;
  reg  line_637_valid_reg;
  wire  line_638_clock;
  wire  line_638_reset;
  wire  line_638_valid;
  reg  line_638_valid_reg;
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire  line_639_clock;
  wire  line_639_reset;
  wire  line_639_valid;
  reg  line_639_valid_reg;
  wire  line_640_clock;
  wire  line_640_reset;
  wire  line_640_valid;
  reg  line_640_valid_reg;
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire  line_641_clock;
  wire  line_641_reset;
  wire  line_641_valid;
  reg  line_641_valid_reg;
  wire  line_642_clock;
  wire  line_642_reset;
  wire  line_642_valid;
  reg  line_642_valid_reg;
  reg [86:0] memuser; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  wire  line_643_clock;
  wire  line_643_reset;
  wire  line_643_valid;
  reg  line_643_valid_reg;
  GEN_w1_line #(.COVER_INDEX(613)) line_613 (
    .clock(line_613_clock),
    .reset(line_613_reset),
    .valid(line_613_valid)
  );
  GEN_w1_line #(.COVER_INDEX(614)) line_614 (
    .clock(line_614_clock),
    .reset(line_614_reset),
    .valid(line_614_valid)
  );
  GEN_w1_line #(.COVER_INDEX(615)) line_615 (
    .clock(line_615_clock),
    .reset(line_615_reset),
    .valid(line_615_valid)
  );
  GEN_w1_line #(.COVER_INDEX(616)) line_616 (
    .clock(line_616_clock),
    .reset(line_616_reset),
    .valid(line_616_valid)
  );
  GEN_w1_line #(.COVER_INDEX(617)) line_617 (
    .clock(line_617_clock),
    .reset(line_617_reset),
    .valid(line_617_valid)
  );
  GEN_w1_line #(.COVER_INDEX(618)) line_618 (
    .clock(line_618_clock),
    .reset(line_618_reset),
    .valid(line_618_valid)
  );
  GEN_w1_line #(.COVER_INDEX(619)) line_619 (
    .clock(line_619_clock),
    .reset(line_619_reset),
    .valid(line_619_valid)
  );
  GEN_w1_line #(.COVER_INDEX(620)) line_620 (
    .clock(line_620_clock),
    .reset(line_620_reset),
    .valid(line_620_valid)
  );
  GEN_w1_line #(.COVER_INDEX(621)) line_621 (
    .clock(line_621_clock),
    .reset(line_621_reset),
    .valid(line_621_valid)
  );
  GEN_w1_line #(.COVER_INDEX(622)) line_622 (
    .clock(line_622_clock),
    .reset(line_622_reset),
    .valid(line_622_valid)
  );
  GEN_w1_line #(.COVER_INDEX(623)) line_623 (
    .clock(line_623_clock),
    .reset(line_623_reset),
    .valid(line_623_valid)
  );
  GEN_w1_line #(.COVER_INDEX(624)) line_624 (
    .clock(line_624_clock),
    .reset(line_624_reset),
    .valid(line_624_valid)
  );
  GEN_w1_line #(.COVER_INDEX(625)) line_625 (
    .clock(line_625_clock),
    .reset(line_625_reset),
    .valid(line_625_valid)
  );
  GEN_w1_line #(.COVER_INDEX(626)) line_626 (
    .clock(line_626_clock),
    .reset(line_626_reset),
    .valid(line_626_valid)
  );
  GEN_w1_line #(.COVER_INDEX(627)) line_627 (
    .clock(line_627_clock),
    .reset(line_627_reset),
    .valid(line_627_valid)
  );
  GEN_w1_line #(.COVER_INDEX(628)) line_628 (
    .clock(line_628_clock),
    .reset(line_628_reset),
    .valid(line_628_valid)
  );
  GEN_w1_line #(.COVER_INDEX(629)) line_629 (
    .clock(line_629_clock),
    .reset(line_629_reset),
    .valid(line_629_valid)
  );
  GEN_w1_line #(.COVER_INDEX(630)) line_630 (
    .clock(line_630_clock),
    .reset(line_630_reset),
    .valid(line_630_valid)
  );
  GEN_w1_line #(.COVER_INDEX(631)) line_631 (
    .clock(line_631_clock),
    .reset(line_631_reset),
    .valid(line_631_valid)
  );
  GEN_w1_line #(.COVER_INDEX(632)) line_632 (
    .clock(line_632_clock),
    .reset(line_632_reset),
    .valid(line_632_valid)
  );
  GEN_w1_line #(.COVER_INDEX(633)) line_633 (
    .clock(line_633_clock),
    .reset(line_633_reset),
    .valid(line_633_valid)
  );
  GEN_w1_line #(.COVER_INDEX(634)) line_634 (
    .clock(line_634_clock),
    .reset(line_634_reset),
    .valid(line_634_valid)
  );
  GEN_w1_line #(.COVER_INDEX(635)) line_635 (
    .clock(line_635_clock),
    .reset(line_635_reset),
    .valid(line_635_valid)
  );
  GEN_w1_line #(.COVER_INDEX(636)) line_636 (
    .clock(line_636_clock),
    .reset(line_636_reset),
    .valid(line_636_valid)
  );
  GEN_w1_line #(.COVER_INDEX(637)) line_637 (
    .clock(line_637_clock),
    .reset(line_637_reset),
    .valid(line_637_valid)
  );
  GEN_w1_line #(.COVER_INDEX(638)) line_638 (
    .clock(line_638_clock),
    .reset(line_638_reset),
    .valid(line_638_valid)
  );
  GEN_w1_line #(.COVER_INDEX(639)) line_639 (
    .clock(line_639_clock),
    .reset(line_639_reset),
    .valid(line_639_valid)
  );
  GEN_w1_line #(.COVER_INDEX(640)) line_640 (
    .clock(line_640_clock),
    .reset(line_640_reset),
    .valid(line_640_valid)
  );
  GEN_w1_line #(.COVER_INDEX(641)) line_641 (
    .clock(line_641_clock),
    .reset(line_641_reset),
    .valid(line_641_valid)
  );
  GEN_w1_line #(.COVER_INDEX(642)) line_642 (
    .clock(line_642_clock),
    .reset(line_642_reset),
    .valid(line_642_valid)
  );
  GEN_w1_line #(.COVER_INDEX(643)) line_643 (
    .clock(line_643_clock),
    .reset(line_643_reset),
    .valid(line_643_valid)
  );
  assign line_613_clock = clock;
  assign line_613_reset = reset;
  assign line_613_valid = _ismmioRec_T ^ line_613_valid_reg;
  assign line_614_clock = clock;
  assign line_614_reset = reset;
  assign line_614_valid = _T_2 ^ line_614_valid_reg;
  assign line_615_clock = clock;
  assign line_615_reset = reset;
  assign line_615_valid = _T_4 ^ line_615_valid_reg;
  assign line_616_clock = clock;
  assign line_616_reset = reset;
  assign line_616_valid = _alreadyOutFire_T ^ line_616_valid_reg;
  assign line_617_clock = clock;
  assign line_617_reset = reset;
  assign line_617_valid = _T_5 ^ line_617_valid_reg;
  assign line_618_clock = clock;
  assign line_618_reset = reset;
  assign line_618_valid = _T_9 ^ line_618_valid_reg;
  assign line_619_clock = clock;
  assign line_619_reset = reset;
  assign line_619_valid = _T_5 ^ line_619_valid_reg;
  assign line_620_clock = clock;
  assign line_620_reset = reset;
  assign line_620_valid = _T_10 ^ line_620_valid_reg;
  assign line_621_clock = clock;
  assign line_621_reset = reset;
  assign line_621_valid = _T_11 ^ line_621_valid_reg;
  assign line_622_clock = clock;
  assign line_622_reset = reset;
  assign line_622_valid = _T_10 ^ line_622_valid_reg;
  assign line_623_clock = clock;
  assign line_623_reset = reset;
  assign line_623_valid = _T_12 ^ line_623_valid_reg;
  assign line_624_clock = clock;
  assign line_624_reset = reset;
  assign line_624_valid = _T_13 ^ line_624_valid_reg;
  assign line_625_clock = clock;
  assign line_625_reset = reset;
  assign line_625_valid = _T_12 ^ line_625_valid_reg;
  assign line_626_clock = clock;
  assign line_626_reset = reset;
  assign line_626_valid = _T_14 ^ line_626_valid_reg;
  assign line_627_clock = clock;
  assign line_627_reset = reset;
  assign line_627_valid = _T_15 ^ line_627_valid_reg;
  assign line_628_clock = clock;
  assign line_628_reset = reset;
  assign line_628_valid = _T_14 ^ line_628_valid_reg;
  assign line_629_clock = clock;
  assign line_629_reset = reset;
  assign line_629_valid = _T_16 ^ line_629_valid_reg;
  assign line_630_clock = clock;
  assign line_630_reset = reset;
  assign line_630_valid = _T_18 ^ line_630_valid_reg;
  assign line_631_clock = clock;
  assign line_631_reset = reset;
  assign line_631_valid = _T_16 ^ line_631_valid_reg;
  assign line_632_clock = clock;
  assign line_632_reset = reset;
  assign line_632_valid = _T_19 ^ line_632_valid_reg;
  assign line_633_clock = clock;
  assign line_633_reset = reset;
  assign line_633_valid = _T_22 ^ line_633_valid_reg;
  assign line_634_clock = clock;
  assign line_634_reset = reset;
  assign line_634_valid = _ismmioRec_T ^ line_634_valid_reg;
  assign line_635_clock = clock;
  assign line_635_reset = reset;
  assign line_635_valid = _ismmioRec_T ^ line_635_valid_reg;
  assign line_636_clock = clock;
  assign line_636_reset = reset;
  assign line_636_valid = _ismmioRec_T ^ line_636_valid_reg;
  assign line_637_clock = clock;
  assign line_637_reset = reset;
  assign line_637_valid = _ismmioRec_T ^ line_637_valid_reg;
  assign line_638_clock = clock;
  assign line_638_reset = reset;
  assign line_638_valid = _ismmioRec_T ^ line_638_valid_reg;
  assign line_639_clock = clock;
  assign line_639_reset = reset;
  assign line_639_valid = _T_17 ^ line_639_valid_reg;
  assign line_640_clock = clock;
  assign line_640_reset = reset;
  assign line_640_valid = _T_17 ^ line_640_valid_reg;
  assign line_641_clock = clock;
  assign line_641_reset = reset;
  assign line_641_valid = _T_13 ^ line_641_valid_reg;
  assign line_642_clock = clock;
  assign line_642_reset = reset;
  assign line_642_valid = _T_13 ^ line_642_valid_reg;
  assign line_643_clock = clock;
  assign line_643_reset = reset;
  assign line_643_valid = _ismmioRec_T ^ line_643_valid_reg;
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5 & ~needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 601:47]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_in_resp_bits_user = memuser; // @[src/main/scala/nutcore/mem/Cache.scala 612:93]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T & ~io_flush[0]) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_37;
    end else begin
      state <= _GEN_43;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    line_613_valid_reg <= _ismmioRec_T;
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    end else if (state == 3'h0 & needFlush) begin // @[src/main/scala/nutcore/mem/Cache.scala 568:40]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 568:52]
    end else begin
      needFlush <= _GEN_32;
    end
    line_614_valid_reg <= _T_2;
    line_615_valid_reg <= _T_4;
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_34;
    end
    line_616_valid_reg <= _alreadyOutFire_T;
    line_617_valid_reg <= _T_5;
    line_618_valid_reg <= _T_9;
    line_619_valid_reg <= _T_5;
    line_620_valid_reg <= _T_10;
    line_621_valid_reg <= _T_11;
    line_622_valid_reg <= _T_10;
    line_623_valid_reg <= _T_12;
    line_624_valid_reg <= _T_13;
    line_625_valid_reg <= _T_12;
    line_626_valid_reg <= _T_14;
    line_627_valid_reg <= _T_15;
    line_628_valid_reg <= _T_14;
    line_629_valid_reg <= _T_16;
    line_630_valid_reg <= _T_18;
    line_631_valid_reg <= _T_16;
    line_632_valid_reg <= _T_19;
    line_633_valid_reg <= _T_22;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    line_634_valid_reg <= _ismmioRec_T;
    line_635_valid_reg <= _ismmioRec_T;
    line_636_valid_reg <= _ismmioRec_T;
    line_637_valid_reg <= _ismmioRec_T;
    line_638_valid_reg <= _ismmioRec_T;
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    line_639_valid_reg <= _T_17;
    line_640_valid_reg <= _T_17;
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    line_641_valid_reg <= _T_13;
    line_642_valid_reg <= _T_13;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
      memuser <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    line_643_valid_reg <= _ismmioRec_T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_613_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  needFlush = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_614_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_615_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  alreadyOutFire = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_616_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_617_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_618_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_619_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_620_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_621_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_622_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_623_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_624_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_625_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_626_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_627_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_628_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_629_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_630_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_631_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_632_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_633_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  reqaddr = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  line_634_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_635_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_636_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_637_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_638_valid_reg = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  mmiordata = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  line_639_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_640_valid_reg = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  memrdata = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  line_641_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_642_valid_reg = _RAND_36[0:0];
  _RAND_37 = {3{`RANDOM}};
  memuser = _RAND_37[86:0];
  _RAND_38 = {1{`RANDOM}};
  line_643_valid_reg = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_alreadyOutFire_T) begin
      cover(1'h1);
    end
    //
    if (_T_5) begin
      cover(1'h1);
    end
    //
    if (_T_5 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_5) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & _T_10 & _T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & _T_12 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & _T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & _T_14 & _T_15) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & _T_16) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & _T_16 & _T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16 & _T_19) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16 & _T_19 & _T_22) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_T_17) begin
      cover(1'h1);
    end
    //
    if (_T_17) begin
      cover(1'h1);
    end
    //
    if (_T_13) begin
      cover(1'h1);
    end
    //
    if (_T_13) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [2:0]   io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [3:0]   io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [7:0]   io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [2:0]   io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [7:0]   io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_out_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          lr_0,
  input          scInflight_0,
  input          ISAMO,
  input  [63:0]  lr_addr,
  output [55:0]  paddr_0,
  output         scIsSuccess_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_r = hitMeta_flag[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire [7:0] _hitRefillFlag_T_1 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 269:26]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  _hitCheck_T_7 = ~io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:31]
  wire  _hitExec_T_1 = hitCheck & ~hitADCheck; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:26]
  wire  hitLoad = _hitExec_T_1 & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 276:41]
  wire  hitStore = _hitExec_T_1 & hitFlag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:42]
  reg  io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
  reg  io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
  reg  io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
  reg  io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
  wire  _loadPF_T_5 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _loadPF_T_7 = ~hitLoad & _loadPF_T_5 & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:40]
  wire  _loadPF_T_8 = ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:50]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  line_644_clock;
  wire  line_644_reset;
  wire  line_644_valid;
  reg  line_644_valid_reg;
  wire  _GEN_44 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  _T_4 = 3'h0 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_645_clock;
  wire  line_645_reset;
  wire  line_645_valid;
  reg  line_645_valid_reg;
  wire  line_646_clock;
  wire  line_646_reset;
  wire  line_646_valid;
  reg  line_646_valid_reg;
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  line_647_clock;
  wire  line_647_reset;
  wire  line_647_valid;
  reg  line_647_valid_reg;
  wire  _T_9 = 3'h1 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_648_clock;
  wire  line_648_reset;
  wire  line_648_valid;
  reg  line_648_valid_reg;
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_649_clock;
  wire  line_649_reset;
  wire  line_649_valid;
  reg  line_649_valid_reg;
  wire  line_650_clock;
  wire  line_650_reset;
  wire  line_650_valid;
  reg  line_650_valid_reg;
  wire  line_651_clock;
  wire  line_651_reset;
  wire  line_651_valid;
  reg  line_651_valid_reg;
  wire [2:0] _GEN_57 = raddrCancel ? 3'h5 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:59]
  wire  _GEN_58 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire  line_652_clock;
  wire  line_652_reset;
  wire  line_652_valid;
  reg  line_652_valid_reg;
  wire  _T_11 = 3'h2 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_653_clock;
  wire  line_653_reset;
  wire  line_653_valid;
  reg  line_653_valid_reg;
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_654_clock;
  wire  line_654_reset;
  wire  line_654_valid;
  reg  line_654_valid_reg;
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_18 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:49]
  wire  line_655_clock;
  wire  line_655_reset;
  wire  line_655_valid;
  reg  line_655_valid_reg;
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire  _T_22 = ~missflag_v | ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:28]
  wire  line_656_clock;
  wire  line_656_reset;
  wire  line_656_valid;
  reg  line_656_valid_reg;
  wire  _loadPF_T_16 = _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:38]
  wire  _storePF_T_15 = io_in_bits_cmd[0] | ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 361:40]
  wire  line_657_clock;
  wire  line_657_reset;
  wire  line_657_valid;
  reg  line_657_valid_reg;
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire  line_658_clock;
  wire  line_658_reset;
  wire  line_658_valid;
  reg  line_658_valid_reg;
  wire [2:0] _GEN_64 = is_reserved ? 3'h5 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 377:23]
  wire  _GEN_65 = is_reserved ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 371:32 378:24]
  wire  _GEN_66 = is_reserved ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 371:32 379:25]
  wire [2:0] _GEN_67 = ~missflag_v | ~missflag_r & missflag_w ? 3'h5 : _GEN_64; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:73]
  wire  _GEN_68 = ~missflag_v | ~missflag_r & missflag_w ? _loadPF_T_5 & _loadPF_T_8 : _GEN_65; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 360:22]
  wire  _GEN_69 = ~missflag_v | ~missflag_r & missflag_w ? io_in_bits_cmd[0] | ISAMO : _GEN_66; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 361:23]
  wire [55:0] _GEN_70 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire  line_659_clock;
  wire  line_659_reset;
  wire  line_659_valid;
  reg  line_659_valid_reg;
  wire  _T_23 = level != 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:27]
  wire  line_660_clock;
  wire  line_660_reset;
  wire  line_660_valid;
  reg  line_660_valid_reg;
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_172 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_172; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u & _hitCheck_T_7); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a | ~missflag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:36]
  wire  _permExec_T_5 = permCheck & ~_T_21 & ~permAD & ~misaligned; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:60]
  wire  permLoad = _permExec_T_5 & (missflag_r | io_pf_status_mxr & missflag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 390:75]
  wire  permStore = _permExec_T_5 & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 391:76]
  wire [63:0] updateData = {56'h0,io_in_bits_cmd[0],7'h40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 392:31]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = _hitRefillFlag_T_1 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | updateData; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire  _T_34 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 403:46]
  wire  line_661_clock;
  wire  line_661_reset;
  wire  line_661_valid;
  reg  line_661_valid_reg;
  wire  line_662_clock;
  wire  line_662_reset;
  wire  line_662_valid;
  reg  line_662_valid_reg;
  wire [2:0] _GEN_71 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 3'h5 : 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 403:80 404:21 408:21]
  wire  _GEN_72 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit
     & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 403:80 405:22]
  wire  _GEN_73 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[
    0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 403:80 406:23]
  wire  _GEN_74 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 403:80 409:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_75 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_76 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire [2:0] _GEN_77 = level != 2'h0 ? _GEN_71 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_78 = level != 2'h0 ? _GEN_72 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 383:36]
  wire  _GEN_79 = level != 2'h0 ? _GEN_73 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 383:36]
  wire  _GEN_80 = level != 2'h0 & _GEN_74; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_81 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_90 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_81; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_109 = _T_12 ? _GEN_90 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_137 = 3'h2 == state ? _GEN_109 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_152 = 3'h1 == state ? 18'h3ffff : _GEN_137; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_152; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_82 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_83 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_67 : _GEN_77; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_84 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_68 : _GEN_78; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_85 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_69 : _GEN_79; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_86 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_70 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_87 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_75; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_88 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_76; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_89 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_91 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_82; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_101 = _T_12 ? _GEN_83 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_103 = _T_12 ? _GEN_84 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 351:33]
  wire  _GEN_104 = _T_12 ? _GEN_85 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 351:33]
  wire  _GEN_108 = _T_12 & _GEN_89; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_111 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire  line_663_clock;
  wire  line_663_reset;
  wire  line_663_valid;
  reg  line_663_valid_reg;
  wire  _T_35 = 3'h3 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_664_clock;
  wire  line_664_reset;
  wire  line_664_valid;
  reg  line_664_valid_reg;
  wire  line_665_clock;
  wire  line_665_reset;
  wire  line_665_valid;
  reg  line_665_valid_reg;
  wire [2:0] _GEN_112 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire  line_666_clock;
  wire  line_666_reset;
  wire  line_666_valid;
  reg  line_666_valid_reg;
  wire  _T_37 = 3'h4 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_667_clock;
  wire  line_667_reset;
  wire  line_667_valid;
  reg  line_667_valid_reg;
  wire  _T_39 = io_isFinish | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:53]
  wire  line_668_clock;
  wire  line_668_reset;
  wire  line_668_valid;
  reg  line_668_valid_reg;
  wire [2:0] _GEN_114 = io_isFinish | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_116 = io_isFinish | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_117 = io_isFinish | alreadyOutFire ? 1'h0 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire  line_669_clock;
  wire  line_669_reset;
  wire  line_669_valid;
  reg  line_669_valid_reg;
  wire  _T_40 = 3'h5 == state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  line_670_clock;
  wire  line_670_reset;
  wire  line_670_valid;
  reg  line_670_valid_reg;
  wire [2:0] _GEN_118 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_119 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_120 = 3'h4 == state ? _GEN_114 : _GEN_118; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_122 = 3'h4 == state ? _GEN_116 : _GEN_119; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_123 = 3'h4 == state ? _GEN_117 : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_124 = 3'h3 == state ? _GEN_112 : _GEN_120; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_127 = 3'h3 == state ? missPTEAF : _GEN_122; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_128 = 3'h3 == state ? _GEN_44 : _GEN_123; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_131 = 3'h2 == state ? _GEN_103 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_132 = 3'h2 == state ? _GEN_104 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_146 = 3'h1 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_131; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_147 = 3'h1 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_132; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_151 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_108; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  loadPF = 3'h0 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_146; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  storePF = 3'h0 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_147; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_151; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _T_45 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  line_671_clock;
  wire  line_671_reset;
  wire  line_671_valid;
  reg  line_671_valid_reg;
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_59 = ~scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:12]
  wire  _T_65 = ~reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
  wire  line_672_clock;
  wire  line_672_reset;
  wire  line_672_valid;
  reg  line_672_valid_reg;
  wire  _T_66 = ~(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
  wire  line_673_clock;
  wire  line_673_reset;
  wire  line_673_valid;
  reg  line_673_valid_reg;
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire [63:0] _GEN_173 = {{8'd0}, paddr}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:49]
  wire  _scIsSuccess_T_7 = hit | state == 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:81]
  wire  out_req_valid = io_in_valid & _scIsSuccess_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _ldReqAF_T_2 = paddr >= 56'h38000000 & paddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_5 = paddr >= 56'h3c000000 & paddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_8 = paddr >= 56'h40600000 & paddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_11 = paddr >= 56'h50000000 & paddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_14 = paddr >= 56'h40001000 & paddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_17 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_20 = paddr >= 56'h40002000 & paddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_23 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _ldReqAF_T_24 = {_ldReqAF_T_23,_ldReqAF_T_20,_ldReqAF_T_17,_ldReqAF_T_14,_ldReqAF_T_11,_ldReqAF_T_8,
    _ldReqAF_T_5,_ldReqAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _ldReqAF_T_25 = |_ldReqAF_T_24; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  ldReqAF = out_req_valid & ~_ldReqAF_T_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 489:34]
  wire  loadAF = (ldReqAF | missPTEAF) & _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 491:54]
  wire  storeAF = ldReqAF & io_in_bits_cmd[0] | ldReqAF & _loadPF_T_5 & ISAMO | missPTEAF & _storePF_T_15; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 492:79]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _hasException_T_2 = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  hasException = _hasException_T_2 | loadPF | storePF | loadAF | storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 494:72]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  wire  scIsSuccess = _T_59 | lr_0 & lr_addr == _GEN_173 | ~(hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:60]
  GEN_w1_line #(.COVER_INDEX(644)) line_644 (
    .clock(line_644_clock),
    .reset(line_644_reset),
    .valid(line_644_valid)
  );
  GEN_w1_line #(.COVER_INDEX(645)) line_645 (
    .clock(line_645_clock),
    .reset(line_645_reset),
    .valid(line_645_valid)
  );
  GEN_w1_line #(.COVER_INDEX(646)) line_646 (
    .clock(line_646_clock),
    .reset(line_646_reset),
    .valid(line_646_valid)
  );
  GEN_w1_line #(.COVER_INDEX(647)) line_647 (
    .clock(line_647_clock),
    .reset(line_647_reset),
    .valid(line_647_valid)
  );
  GEN_w1_line #(.COVER_INDEX(648)) line_648 (
    .clock(line_648_clock),
    .reset(line_648_reset),
    .valid(line_648_valid)
  );
  GEN_w1_line #(.COVER_INDEX(649)) line_649 (
    .clock(line_649_clock),
    .reset(line_649_reset),
    .valid(line_649_valid)
  );
  GEN_w1_line #(.COVER_INDEX(650)) line_650 (
    .clock(line_650_clock),
    .reset(line_650_reset),
    .valid(line_650_valid)
  );
  GEN_w1_line #(.COVER_INDEX(651)) line_651 (
    .clock(line_651_clock),
    .reset(line_651_reset),
    .valid(line_651_valid)
  );
  GEN_w1_line #(.COVER_INDEX(652)) line_652 (
    .clock(line_652_clock),
    .reset(line_652_reset),
    .valid(line_652_valid)
  );
  GEN_w1_line #(.COVER_INDEX(653)) line_653 (
    .clock(line_653_clock),
    .reset(line_653_reset),
    .valid(line_653_valid)
  );
  GEN_w1_line #(.COVER_INDEX(654)) line_654 (
    .clock(line_654_clock),
    .reset(line_654_reset),
    .valid(line_654_valid)
  );
  GEN_w1_line #(.COVER_INDEX(655)) line_655 (
    .clock(line_655_clock),
    .reset(line_655_reset),
    .valid(line_655_valid)
  );
  GEN_w1_line #(.COVER_INDEX(656)) line_656 (
    .clock(line_656_clock),
    .reset(line_656_reset),
    .valid(line_656_valid)
  );
  GEN_w1_line #(.COVER_INDEX(657)) line_657 (
    .clock(line_657_clock),
    .reset(line_657_reset),
    .valid(line_657_valid)
  );
  GEN_w1_line #(.COVER_INDEX(658)) line_658 (
    .clock(line_658_clock),
    .reset(line_658_reset),
    .valid(line_658_valid)
  );
  GEN_w1_line #(.COVER_INDEX(659)) line_659 (
    .clock(line_659_clock),
    .reset(line_659_reset),
    .valid(line_659_valid)
  );
  GEN_w1_line #(.COVER_INDEX(660)) line_660 (
    .clock(line_660_clock),
    .reset(line_660_reset),
    .valid(line_660_valid)
  );
  GEN_w1_line #(.COVER_INDEX(661)) line_661 (
    .clock(line_661_clock),
    .reset(line_661_reset),
    .valid(line_661_valid)
  );
  GEN_w1_line #(.COVER_INDEX(662)) line_662 (
    .clock(line_662_clock),
    .reset(line_662_reset),
    .valid(line_662_valid)
  );
  GEN_w1_line #(.COVER_INDEX(663)) line_663 (
    .clock(line_663_clock),
    .reset(line_663_reset),
    .valid(line_663_valid)
  );
  GEN_w1_line #(.COVER_INDEX(664)) line_664 (
    .clock(line_664_clock),
    .reset(line_664_reset),
    .valid(line_664_valid)
  );
  GEN_w1_line #(.COVER_INDEX(665)) line_665 (
    .clock(line_665_clock),
    .reset(line_665_reset),
    .valid(line_665_valid)
  );
  GEN_w1_line #(.COVER_INDEX(666)) line_666 (
    .clock(line_666_clock),
    .reset(line_666_reset),
    .valid(line_666_valid)
  );
  GEN_w1_line #(.COVER_INDEX(667)) line_667 (
    .clock(line_667_clock),
    .reset(line_667_reset),
    .valid(line_667_valid)
  );
  GEN_w1_line #(.COVER_INDEX(668)) line_668 (
    .clock(line_668_clock),
    .reset(line_668_reset),
    .valid(line_668_valid)
  );
  GEN_w1_line #(.COVER_INDEX(669)) line_669 (
    .clock(line_669_clock),
    .reset(line_669_reset),
    .valid(line_669_valid)
  );
  GEN_w1_line #(.COVER_INDEX(670)) line_670 (
    .clock(line_670_clock),
    .reset(line_670_reset),
    .valid(line_670_valid)
  );
  GEN_w1_line #(.COVER_INDEX(671)) line_671 (
    .clock(line_671_clock),
    .reset(line_671_reset),
    .valid(line_671_valid)
  );
  GEN_w1_line #(.COVER_INDEX(672)) line_672 (
    .clock(line_672_clock),
    .reset(line_672_reset),
    .valid(line_672_valid)
  );
  GEN_w1_line #(.COVER_INDEX(673)) line_673 (
    .clock(line_673_clock),
    .reset(line_673_reset),
    .valid(line_673_valid)
  );
  assign line_644_clock = clock;
  assign line_644_reset = reset;
  assign line_644_valid = _alreadyOutFire_T ^ line_644_valid_reg;
  assign line_645_clock = clock;
  assign line_645_reset = reset;
  assign line_645_valid = _T_4 ^ line_645_valid_reg;
  assign line_646_clock = clock;
  assign line_646_reset = reset;
  assign line_646_valid = miss ^ line_646_valid_reg;
  assign line_647_clock = clock;
  assign line_647_reset = reset;
  assign line_647_valid = _T_4 ^ line_647_valid_reg;
  assign line_648_clock = clock;
  assign line_648_reset = reset;
  assign line_648_valid = _T_9 ^ line_648_valid_reg;
  assign line_649_clock = clock;
  assign line_649_reset = reset;
  assign line_649_valid = _T_10 ^ line_649_valid_reg;
  assign line_650_clock = clock;
  assign line_650_reset = reset;
  assign line_650_valid = _T_10 ^ line_650_valid_reg;
  assign line_651_clock = clock;
  assign line_651_reset = reset;
  assign line_651_valid = raddrCancel ^ line_651_valid_reg;
  assign line_652_clock = clock;
  assign line_652_reset = reset;
  assign line_652_valid = _T_9 ^ line_652_valid_reg;
  assign line_653_clock = clock;
  assign line_653_reset = reset;
  assign line_653_valid = _T_11 ^ line_653_valid_reg;
  assign line_654_clock = clock;
  assign line_654_reset = reset;
  assign line_654_valid = _T_12 ^ line_654_valid_reg;
  assign line_655_clock = clock;
  assign line_655_reset = reset;
  assign line_655_valid = _T_18 ^ line_655_valid_reg;
  assign line_656_clock = clock;
  assign line_656_reset = reset;
  assign line_656_valid = _T_22 ^ line_656_valid_reg;
  assign line_657_clock = clock;
  assign line_657_reset = reset;
  assign line_657_valid = _T_22 ^ line_657_valid_reg;
  assign line_658_clock = clock;
  assign line_658_reset = reset;
  assign line_658_valid = is_reserved ^ line_658_valid_reg;
  assign line_659_clock = clock;
  assign line_659_reset = reset;
  assign line_659_valid = _T_18 ^ line_659_valid_reg;
  assign line_660_clock = clock;
  assign line_660_reset = reset;
  assign line_660_valid = _T_23 ^ line_660_valid_reg;
  assign line_661_clock = clock;
  assign line_661_reset = reset;
  assign line_661_valid = _T_34 ^ line_661_valid_reg;
  assign line_662_clock = clock;
  assign line_662_reset = reset;
  assign line_662_valid = _T_34 ^ line_662_valid_reg;
  assign line_663_clock = clock;
  assign line_663_reset = reset;
  assign line_663_valid = _T_11 ^ line_663_valid_reg;
  assign line_664_clock = clock;
  assign line_664_reset = reset;
  assign line_664_valid = _T_35 ^ line_664_valid_reg;
  assign line_665_clock = clock;
  assign line_665_reset = reset;
  assign line_665_valid = _T_10 ^ line_665_valid_reg;
  assign line_666_clock = clock;
  assign line_666_reset = reset;
  assign line_666_valid = _T_35 ^ line_666_valid_reg;
  assign line_667_clock = clock;
  assign line_667_reset = reset;
  assign line_667_valid = _T_37 ^ line_667_valid_reg;
  assign line_668_clock = clock;
  assign line_668_reset = reset;
  assign line_668_valid = _T_39 ^ line_668_valid_reg;
  assign line_669_clock = clock;
  assign line_669_reset = reset;
  assign line_669_valid = _T_37 ^ line_669_valid_reg;
  assign line_670_clock = clock;
  assign line_670_reset = reset;
  assign line_670_valid = _T_40 ^ line_670_valid_reg;
  assign line_671_clock = clock;
  assign line_671_reset = reset;
  assign line_671_valid = blockRefill ^ line_671_valid_reg;
  assign line_672_clock = clock;
  assign line_672_reset = reset;
  assign line_672_valid = _T_65 ^ line_672_valid_reg;
  assign line_673_clock = clock;
  assign line_673_reset = reset;
  assign line_673_valid = _T_66 ^ line_673_valid_reg;
  assign io_in_ready = io_out_ready & _T_45 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException & scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:92]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_windex = REG_1; // @[src/main/scala/nutcore/mem/TLB.scala 218:17]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_isFinish = _alreadyOutFire_T | _hasException_T_2 | ~scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:54]
  assign paddr_0 = paddr;
  assign scIsSuccess_0 = scIsSuccess;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
      io_pf_loadPF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= _GEN_103;
    end else begin
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
      io_pf_storePF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= _GEN_104;
    end else begin
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
      io_pf_laf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end else begin
      io_pf_laf_REG <= loadAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
      io_pf_saf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end else begin
      io_pf_saf_REG <= storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 342:15]
      end else begin
        state <= _GEN_57;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_101;
    end else begin
      state <= _GEN_124;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_111;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_88;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_91;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_86;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_44;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_44;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_44;
    end else begin
      alreadyOutFire <= _GEN_128;
    end
    line_644_valid_reg <= _alreadyOutFire_T;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(_T_10)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
          missPTEAF <= _GEN_58;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_127;
      end
    end
    line_645_valid_reg <= _T_4;
    line_646_valid_reg <= miss;
    line_647_valid_reg <= _T_4;
    line_648_valid_reg <= _T_9;
    line_649_valid_reg <= _T_10;
    line_650_valid_reg <= _T_10;
    line_651_valid_reg <= raddrCancel;
    line_652_valid_reg <= _T_9;
    line_653_valid_reg <= _T_11;
    line_654_valid_reg <= _T_12;
    line_655_valid_reg <= _T_18;
    line_656_valid_reg <= _T_22;
    line_657_valid_reg <= _T_22;
    line_658_valid_reg <= is_reserved;
    line_659_valid_reg <= _T_18;
    line_660_valid_reg <= _T_23;
    line_661_valid_reg <= _T_34;
    line_662_valid_reg <= _T_34;
    line_663_valid_reg <= _T_11;
    line_664_valid_reg <= _T_35;
    line_665_valid_reg <= _T_10;
    line_666_valid_reg <= _T_35;
    line_667_valid_reg <= _T_37;
    line_668_valid_reg <= _T_39;
    line_669_valid_reg <= _T_37;
    line_670_valid_reg <= _T_40;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else begin
      REG <= 3'h2 == state & _GEN_108;
    end
    REG_1 <= io_in_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_90;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_87;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= missMetaRefill & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
    line_671_valid_reg <= blockRefill;
    line_672_valid_reg <= _T_65;
    line_673_valid_reg <= _T_66;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed: SC is inflight but TLB receives a read request\n    at EmbeddedTLB.scala:476 assert(!scInflight || !io.in.valid || req.isWrite(), \"SC is inflight but TLB receives a read request\")\n"
            ); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  io_pf_loadPF_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_pf_storePF_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_pf_laf_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_pf_saf_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  level = _RAND_6[1:0];
  _RAND_7 = {2{`RANDOM}};
  memRespStore = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  missMaskStore = _RAND_8[17:0];
  _RAND_9 = {2{`RANDOM}};
  raddr = _RAND_9[55:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_644_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  missPTEAF = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_645_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_646_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_647_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_648_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_649_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_650_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_651_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_652_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_653_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_654_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_655_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_656_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_657_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_658_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_659_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_660_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_661_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_662_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_663_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_664_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_665_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_666_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_667_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_668_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_669_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_670_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG_1 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  REG_2 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  REG_3 = _RAND_42[26:0];
  _RAND_43 = {1{`RANDOM}};
  REG_4 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  REG_5 = _RAND_44[17:0];
  _RAND_45 = {1{`RANDOM}};
  REG_6 = _RAND_45[7:0];
  _RAND_46 = {2{`RANDOM}};
  REG_7 = _RAND_46[43:0];
  _RAND_47 = {2{`RANDOM}};
  REG_8 = _RAND_47[55:0];
  _RAND_48 = {1{`RANDOM}};
  blockRefill = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_671_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_672_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_673_valid_reg = _RAND_51[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_alreadyOutFire_T) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4 & miss) begin
      cover(1'h1);
    end
    //
    if (~_T_4) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & ~_T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_9 & ~_T_10 & raddrCancel) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18 & _T_22) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18 & ~_T_22) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & _T_18 & ~_T_22 & is_reserved) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & ~_T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & ~_T_18 & _T_23) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & ~_T_18 & _T_23 & _T_34) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & _T_11 & _T_12 & ~_T_18 & _T_23 & ~_T_34) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_35) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_35) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & _T_35 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_35) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_35 & _T_37) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_35 & _T_37 & _T_39) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_35 & ~_T_37) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_9 & ~_T_11 & ~_T_35 & ~_T_37 & _T_40) begin
      cover(1'h1);
    end
    //
    if (blockRefill) begin
      cover(1'h1);
    end
    //
    if (_T_65) begin
      cover(1'h1);
    end
    //
    if (_T_65 & _T_66) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
    end
  end
endmodule
module EmbeddedTLBEmpty_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [63:0] io_out_bits_wdata // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_rindex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  reg [3:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_674_clock;
  wire  line_674_reset;
  wire  line_674_valid;
  reg  line_674_valid_reg;
  wire  wrap_wrap = resetSet == 4'hf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  line_675_clock;
  wire  line_675_reset;
  wire  line_675_valid;
  reg  line_675_valid_reg;
  wire  _GEN_9 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire  wen = resetState | io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 65:16]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  wire  line_676_clock;
  wire  line_676_reset;
  wire  line_676_valid;
  reg  line_676_valid_reg;
  wire  line_677_clock;
  wire  line_677_reset;
  wire  line_677_valid;
  reg  line_677_valid_reg;
  wire  line_678_clock;
  wire  line_678_reset;
  wire  line_678_valid;
  reg  line_678_valid_reg;
  wire  line_679_clock;
  wire  line_679_reset;
  wire  line_679_valid;
  reg  line_679_valid_reg;
  wire  line_680_clock;
  wire  line_680_reset;
  wire  line_680_valid;
  reg  line_680_valid_reg;
  GEN_w1_line #(.COVER_INDEX(674)) line_674 (
    .clock(line_674_clock),
    .reset(line_674_reset),
    .valid(line_674_valid)
  );
  GEN_w1_line #(.COVER_INDEX(675)) line_675 (
    .clock(line_675_clock),
    .reset(line_675_reset),
    .valid(line_675_valid)
  );
  GEN_w1_line #(.COVER_INDEX(676)) line_676 (
    .clock(line_676_clock),
    .reset(line_676_reset),
    .valid(line_676_valid)
  );
  GEN_w1_line #(.COVER_INDEX(677)) line_677 (
    .clock(line_677_clock),
    .reset(line_677_reset),
    .valid(line_677_valid)
  );
  GEN_w1_line #(.COVER_INDEX(678)) line_678 (
    .clock(line_678_clock),
    .reset(line_678_reset),
    .valid(line_678_valid)
  );
  GEN_w1_line #(.COVER_INDEX(679)) line_679 (
    .clock(line_679_clock),
    .reset(line_679_reset),
    .valid(line_679_valid)
  );
  GEN_w1_line #(.COVER_INDEX(680)) line_680 (
    .clock(line_680_clock),
    .reset(line_680_reset),
    .valid(line_680_valid)
  );
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign line_674_clock = clock;
  assign line_674_reset = reset;
  assign line_674_valid = resetState ^ line_674_valid_reg;
  assign line_675_clock = clock;
  assign line_675_reset = reset;
  assign line_675_valid = resetFinish ^ line_675_valid_reg;
  assign line_676_clock = clock;
  assign line_676_reset = reset;
  assign line_676_valid = wen ^ line_676_valid_reg;
  assign line_677_clock = clock;
  assign line_677_reset = reset;
  assign line_677_valid = waymask[0] ^ line_677_valid_reg;
  assign line_678_clock = clock;
  assign line_678_reset = reset;
  assign line_678_valid = waymask[1] ^ line_678_valid_reg;
  assign line_679_clock = clock;
  assign line_679_reset = reset;
  assign line_679_valid = waymask[2] ^ line_679_valid_reg;
  assign line_680_clock = clock;
  assign line_680_reset = reset;
  assign line_680_valid = waymask[3] ^ line_680_valid_reg;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_9; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    line_674_valid_reg <= resetState;
    line_675_valid_reg <= resetFinish;
    line_676_valid_reg <= wen;
    line_677_valid_reg <= waymask[0];
    line_678_valid_reg <= waymask[1];
    line_679_valid_reg <= waymask[2];
    line_680_valid_reg <= waymask[3];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  line_674_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_675_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_676_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_677_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_678_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_679_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_680_valid_reg = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (resetState) begin
      cover(1'h1);
    end
    //
    if (resetFinish) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[0]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[1]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[2]) begin
      cover(1'h1);
    end
    //
    if (wen & waymask[3]) begin
      cover(1'h1);
    end
  end
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         lr,
  input         scInflight,
  input         amoReq,
  input  [63:0] lrAddr,
  output [55:0] paddr,
  input  [63:0] CSRSATP,
  output        _T_12_0,
  output        scIsSuccess_0,
  output        vmEnable_0,
  input         MOUFlushTLB,
  output        tlbFinish_0,
  output        _T_13_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_lr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_lr_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [55:0] tlbExec_paddr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbEmpty_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_rindex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  wire  line_681_clock;
  wire  line_681_reset;
  wire  line_681_valid;
  reg  line_681_valid_reg;
  wire  _lastReqAddr_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_682_clock;
  wire  line_682_reset;
  wire  line_682_valid;
  reg  line_682_valid_reg;
  wire  line_683_clock;
  wire  line_683_reset;
  wire  line_683_valid;
  reg  line_683_valid_reg;
  wire  line_684_clock;
  wire  line_684_reset;
  wire  line_684_valid;
  reg  line_684_valid_reg;
  wire  line_685_clock;
  wire  line_685_reset;
  wire  line_685_valid;
  reg  line_685_valid_reg;
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  line_686_clock;
  wire  line_686_reset;
  wire  line_686_valid;
  reg  line_686_valid_reg;
  wire  _GEN_24 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _T_6 = mdUpdate & vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:37]
  wire  line_687_clock;
  wire  line_687_reset;
  wire  line_687_valid;
  reg  line_687_valid_reg;
  wire  _GEN_25 = mdUpdate & vmEnable | _GEN_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [2:0] tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [3:0] tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [7:0] tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [63:0] tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  line_688_clock;
  wire  line_688_reset;
  wire  line_688_valid;
  reg  line_688_valid_reg;
  wire  _T_7 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  line_689_clock;
  wire  line_689_reset;
  wire  line_689_valid;
  reg  line_689_valid_reg;
  wire  _GEN_32 = _T_7 ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_8 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  line_690_clock;
  wire  line_690_reset;
  wire  line_690_valid;
  reg  line_690_valid_reg;
  wire  _GEN_33 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_32; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  line_691_clock;
  wire  line_691_reset;
  wire  line_691_valid;
  reg  line_691_valid_reg;
  wire  _T_9 = ~vmEnable; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:8]
  wire  line_692_clock;
  wire  line_692_reset;
  wire  line_692_valid;
  reg  line_692_valid_reg;
  wire  line_693_clock;
  wire  line_693_reset;
  wire  line_693_valid;
  reg  line_693_valid_reg;
  wire  _alreadyOutFinish_T_1 = tlbExec_io_out_valid & ~tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:76]
  reg  alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
  wire  line_694_clock;
  wire  line_694_reset;
  wire  line_694_valid;
  reg  line_694_valid_reg;
  wire  _GEN_53 = tlbExec_io_out_valid & ~tlbExec_io_out_ready | alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:{37,37,37}]
  wire  _T_10 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_11 = alreadyOutFinish & _T_10; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:27]
  wire  line_695_clock;
  wire  line_695_reset;
  wire  line_695_valid;
  reg  line_695_valid_reg;
  wire  _tlbFinish_T_2 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _tlbFinish_T_3 = tlbExec_io_pf_laf | tlbExec_io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _tlbFinish_T_4 = _tlbFinish_T_2 | _tlbFinish_T_3; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  tlbFinish = tlbExec_io_out_valid & ~alreadyOutFinish | _tlbFinish_T_4 | ~scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 180:95]
  wire  _T_12 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _T_13 = io_csrMMU_laf | io_csrMMU_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  EmbeddedTLBExec_1 tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_isFinish(tlbExec_io_isFinish),
    .lr_0(tlbExec_lr_0),
    .scInflight_0(tlbExec_scInflight_0),
    .ISAMO(tlbExec_ISAMO),
    .lr_addr(tlbExec_lr_addr),
    .paddr_0(tlbExec_paddr_0),
    .scIsSuccess_0(tlbExec_scIsSuccess_0)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
    .clock(tlbEmpty_clock),
    .reset(tlbEmpty_reset),
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  GEN_w1_line #(.COVER_INDEX(681)) line_681 (
    .clock(line_681_clock),
    .reset(line_681_reset),
    .valid(line_681_valid)
  );
  GEN_w1_line #(.COVER_INDEX(682)) line_682 (
    .clock(line_682_clock),
    .reset(line_682_reset),
    .valid(line_682_valid)
  );
  GEN_w1_line #(.COVER_INDEX(683)) line_683 (
    .clock(line_683_clock),
    .reset(line_683_reset),
    .valid(line_683_valid)
  );
  GEN_w1_line #(.COVER_INDEX(684)) line_684 (
    .clock(line_684_clock),
    .reset(line_684_reset),
    .valid(line_684_valid)
  );
  GEN_w1_line #(.COVER_INDEX(685)) line_685 (
    .clock(line_685_clock),
    .reset(line_685_reset),
    .valid(line_685_valid)
  );
  GEN_w1_line #(.COVER_INDEX(686)) line_686 (
    .clock(line_686_clock),
    .reset(line_686_reset),
    .valid(line_686_valid)
  );
  GEN_w1_line #(.COVER_INDEX(687)) line_687 (
    .clock(line_687_clock),
    .reset(line_687_reset),
    .valid(line_687_valid)
  );
  GEN_w1_line #(.COVER_INDEX(688)) line_688 (
    .clock(line_688_clock),
    .reset(line_688_reset),
    .valid(line_688_valid)
  );
  GEN_w1_line #(.COVER_INDEX(689)) line_689 (
    .clock(line_689_clock),
    .reset(line_689_reset),
    .valid(line_689_valid)
  );
  GEN_w1_line #(.COVER_INDEX(690)) line_690 (
    .clock(line_690_clock),
    .reset(line_690_reset),
    .valid(line_690_valid)
  );
  GEN_w1_line #(.COVER_INDEX(691)) line_691 (
    .clock(line_691_clock),
    .reset(line_691_reset),
    .valid(line_691_valid)
  );
  GEN_w1_line #(.COVER_INDEX(692)) line_692 (
    .clock(line_692_clock),
    .reset(line_692_reset),
    .valid(line_692_valid)
  );
  GEN_w1_line #(.COVER_INDEX(693)) line_693 (
    .clock(line_693_clock),
    .reset(line_693_reset),
    .valid(line_693_valid)
  );
  GEN_w1_line #(.COVER_INDEX(694)) line_694 (
    .clock(line_694_clock),
    .reset(line_694_reset),
    .valid(line_694_valid)
  );
  GEN_w1_line #(.COVER_INDEX(695)) line_695 (
    .clock(line_695_clock),
    .reset(line_695_reset),
    .valid(line_695_valid)
  );
  assign line_681_clock = clock;
  assign line_681_reset = reset;
  assign line_681_valid = mdUpdate ^ line_681_valid_reg;
  assign line_682_clock = clock;
  assign line_682_reset = reset;
  assign line_682_valid = _lastReqAddr_T ^ line_682_valid_reg;
  assign line_683_clock = clock;
  assign line_683_reset = reset;
  assign line_683_valid = io_in_resp_valid ^ line_683_valid_reg;
  assign line_684_clock = clock;
  assign line_684_reset = reset;
  assign line_684_valid = io_in_resp_valid ^ line_684_valid_reg;
  assign line_685_clock = clock;
  assign line_685_reset = reset;
  assign line_685_valid = _lastReqAddr_T ^ line_685_valid_reg;
  assign line_686_clock = clock;
  assign line_686_reset = reset;
  assign line_686_valid = tlbExec_io_isFinish ^ line_686_valid_reg;
  assign line_687_clock = clock;
  assign line_687_reset = reset;
  assign line_687_valid = _T_6 ^ line_687_valid_reg;
  assign line_688_clock = clock;
  assign line_688_reset = reset;
  assign line_688_valid = mdUpdate ^ line_688_valid_reg;
  assign line_689_clock = clock;
  assign line_689_reset = reset;
  assign line_689_valid = _T_7 ^ line_689_valid_reg;
  assign line_690_clock = clock;
  assign line_690_reset = reset;
  assign line_690_valid = _T_8 ^ line_690_valid_reg;
  assign line_691_clock = clock;
  assign line_691_reset = reset;
  assign line_691_valid = _T_8 ^ line_691_valid_reg;
  assign line_692_clock = clock;
  assign line_692_reset = reset;
  assign line_692_valid = _T_9 ^ line_692_valid_reg;
  assign line_693_clock = clock;
  assign line_693_reset = reset;
  assign line_693_valid = _T_9 ^ line_693_valid_reg;
  assign line_694_clock = clock;
  assign line_694_reset = reset;
  assign line_694_valid = _alreadyOutFinish_T_1 ^ line_694_valid_reg;
  assign line_695_clock = clock;
  assign line_695_reset = reset;
  assign line_695_valid = _T_11 ^ line_695_valid_reg;
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19 149:23]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 148:24 169:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 169:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 163:26 169:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 164:25 169:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 165:27 169:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 166:27 169:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_csrMMU_loadPF = ~vmEnable ? 1'h0 : tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 150:24 95:17]
  assign io_csrMMU_storePF = ~vmEnable ? 1'h0 : tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 151:25 95:17]
  assign io_csrMMU_laf = ~vmEnable ? 1'h0 : tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 152:21 95:17]
  assign io_csrMMU_saf = ~vmEnable ? 1'h0 : tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 153:21 95:17]
  assign paddr = tlbExec_paddr_0;
  assign _T_12_0 = _T_12;
  assign scIsSuccess_0 = tlbExec_scIsSuccess_0;
  assign vmEnable_0 = vmEnable;
  assign tlbFinish_0 = tlbFinish;
  assign _T_13_1 = _T_13;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_size = tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_cmd = tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wmask = tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wdata = tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 src/main/scala/utils/Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_lr_0 = lr;
  assign tlbExec_scInflight_0 = scInflight;
  assign tlbExec_ISAMO = amoReq;
  assign tlbExec_lr_addr = lrAddr;
  assign tlbEmpty_clock = clock;
  assign tlbEmpty_reset = reset;
  assign tlbEmpty_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 147:29 169:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    line_681_valid_reg <= mdUpdate;
    line_682_valid_reg <= _lastReqAddr_T;
    line_683_valid_reg <= io_in_resp_valid;
    line_684_valid_reg <= io_in_resp_valid;
    line_685_valid_reg <= _lastReqAddr_T;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else begin
      valid <= _GEN_25;
    end
    line_686_valid_reg <= tlbExec_io_isFinish;
    line_687_valid_reg <= _T_6;
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    line_688_valid_reg <= mdUpdate;
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_33;
    end
    line_689_valid_reg <= _T_7;
    line_690_valid_reg <= _T_8;
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_addr <= tlbExec_io_out_bits_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_size <= tlbExec_io_out_bits_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_cmd <= tlbExec_io_out_bits_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wmask <= tlbExec_io_out_bits_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wdata <= tlbExec_io_out_bits_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    line_691_valid_reg <= _T_8;
    line_692_valid_reg <= _T_9;
    line_693_valid_reg <= _T_9;
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
    end else if (alreadyOutFinish & _T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:53]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:72]
    end else begin
      alreadyOutFinish <= _GEN_53;
    end
    line_694_valid_reg <= _alreadyOutFinish_T_1;
    line_695_valid_reg <= _T_11;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  line_681_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_682_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_683_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_684_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_685_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_686_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_687_valid_reg = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_12[38:0];
  _RAND_13 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_size = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_cmd = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_wmask = _RAND_15[7:0];
  _RAND_16 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_wdata = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  line_688_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_689_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_690_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_addr = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_size = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_cmd = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_wmask = _RAND_24[7:0];
  _RAND_25 = {2{`RANDOM}};
  tlbEmpty_io_in_bits_r_wdata = _RAND_25[63:0];
  _RAND_26 = {1{`RANDOM}};
  line_691_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_692_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_693_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  alreadyOutFinish = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_694_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_695_valid_reg = _RAND_31[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (mdUpdate) begin
      cover(1'h1);
    end
    //
    if (_lastReqAddr_T) begin
      cover(1'h1);
    end
    //
    if (io_in_resp_valid) begin
      cover(1'h1);
    end
    //
    if (~io_in_resp_valid) begin
      cover(1'h1);
    end
    //
    if (~io_in_resp_valid & _lastReqAddr_T) begin
      cover(1'h1);
    end
    //
    if (tlbExec_io_isFinish) begin
      cover(1'h1);
    end
    //
    if (_T_6) begin
      cover(1'h1);
    end
    //
    if (mdUpdate) begin
      cover(1'h1);
    end
    //
    if (_T_7) begin
      cover(1'h1);
    end
    //
    if (_T_8) begin
      cover(1'h1);
    end
    //
    if (_T_8) begin
      cover(1'h1);
    end
    //
    if (_T_9) begin
      cover(1'h1);
    end
    //
    if (~_T_9) begin
      cover(1'h1);
    end
    //
    if (_alreadyOutFinish_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_11) begin
      cover(1'h1);
    end
  end
endmodule
module PTERequestFilter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_u // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  isLegal = |(io_in_req_bits_addr >= 32'h80000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasInflight_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _hasInflight_T_2 = _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:33]
  wire  line_696_clock;
  wire  line_696_reset;
  wire  line_696_valid;
  reg  line_696_valid_reg;
  wire  _T_1 = ~io_out_resp_valid & hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:28]
  wire  line_697_clock;
  wire  line_697_reset;
  wire  line_697_valid;
  reg  line_697_valid_reg;
  wire [7:0] _io_in_resp_bits_rdata_T = {3'h7,io_u,4'hf}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 570:33]
  GEN_w1_line #(.COVER_INDEX(696)) line_696 (
    .clock(line_696_clock),
    .reset(line_696_reset),
    .valid(line_696_valid)
  );
  GEN_w1_line #(.COVER_INDEX(697)) line_697 (
    .clock(line_697_clock),
    .reset(line_697_reset),
    .valid(line_697_valid)
  );
  assign line_696_clock = clock;
  assign line_696_reset = reset;
  assign line_696_valid = _hasInflight_T_2 ^ line_696_valid_reg;
  assign line_697_clock = clock;
  assign line_697_reset = reset;
  assign line_697_valid = _T_1 ^ line_697_valid_reg;
  assign io_in_req_ready = isLegal ? io_out_req_ready : ~hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 562:25]
  assign io_in_resp_valid = ~io_out_resp_valid & hasInflight | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 567:22]
  assign io_in_resp_bits_rdata = ~io_out_resp_valid & hasInflight ? {{56'd0}, _io_in_resp_bits_rdata_T} :
    io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 570:27]
  assign io_out_req_valid = io_in_req_valid & isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 561:39]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end else if (~io_out_resp_valid & hasInflight) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:44]
      hasInflight <= 1'h0;
    end else begin
      hasInflight <= _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:15]
    end
    line_696_valid_reg <= _hasInflight_T_2;
    line_697_valid_reg <= _T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasInflight = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_696_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_697_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_hasInflight_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module Cache_fake_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_out_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_out_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        ismmio_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  line_698_clock;
  wire  line_698_reset;
  wire  line_698_valid;
  reg  line_698_valid_reg;
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  line_699_clock;
  wire  line_699_reset;
  wire  line_699_valid;
  reg  line_699_valid_reg;
  wire  _GEN_34 = io_in_resp_valid | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_5 = 3'h0 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_700_clock;
  wire  line_700_reset;
  wire  line_700_valid;
  reg  line_700_valid_reg;
  wire  line_701_clock;
  wire  line_701_reset;
  wire  line_701_valid;
  reg  line_701_valid_reg;
  wire  line_702_clock;
  wire  line_702_reset;
  wire  line_702_valid;
  reg  line_702_valid_reg;
  wire  _T_10 = 3'h1 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_703_clock;
  wire  line_703_reset;
  wire  line_703_valid;
  reg  line_703_valid_reg;
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_704_clock;
  wire  line_704_reset;
  wire  line_704_valid;
  reg  line_704_valid_reg;
  wire  line_705_clock;
  wire  line_705_reset;
  wire  line_705_valid;
  reg  line_705_valid_reg;
  wire  _T_12 = 3'h2 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_706_clock;
  wire  line_706_reset;
  wire  line_706_valid;
  reg  line_706_valid_reg;
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_707_clock;
  wire  line_707_reset;
  wire  line_707_valid;
  reg  line_707_valid_reg;
  wire [2:0] _GEN_37 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  line_708_clock;
  wire  line_708_reset;
  wire  line_708_valid;
  reg  line_708_valid_reg;
  wire  _T_14 = 3'h3 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_709_clock;
  wire  line_709_reset;
  wire  line_709_valid;
  reg  line_709_valid_reg;
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_710_clock;
  wire  line_710_reset;
  wire  line_710_valid;
  reg  line_710_valid_reg;
  wire [2:0] _GEN_38 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  line_711_clock;
  wire  line_711_reset;
  wire  line_711_valid;
  reg  line_711_valid_reg;
  wire  _T_16 = 3'h4 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_712_clock;
  wire  line_712_reset;
  wire  line_712_valid;
  reg  line_712_valid_reg;
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_18 = _T_17 | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 587:33]
  wire  line_713_clock;
  wire  line_713_reset;
  wire  line_713_valid;
  reg  line_713_valid_reg;
  wire [2:0] _GEN_39 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire  line_714_clock;
  wire  line_714_reset;
  wire  line_714_valid;
  reg  line_714_valid_reg;
  wire  _T_19 = 3'h5 == state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire  line_715_clock;
  wire  line_715_reset;
  wire  line_715_valid;
  reg  line_715_valid_reg;
  wire  line_716_clock;
  wire  line_716_reset;
  wire  line_716_valid;
  reg  line_716_valid_reg;
  wire [2:0] _GEN_40 = _GEN_34 ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_41 = 3'h5 == state ? _GEN_40 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_42 = 3'h4 == state ? _GEN_39 : _GEN_41; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_43 = 3'h3 == state ? _GEN_38 : _GEN_42; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire  line_717_clock;
  wire  line_717_reset;
  wire  line_717_valid;
  reg  line_717_valid_reg;
  reg [3:0] cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  wire  line_718_clock;
  wire  line_718_reset;
  wire  line_718_valid;
  reg  line_718_valid_reg;
  reg [2:0] size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  wire  line_719_clock;
  wire  line_719_reset;
  wire  line_719_valid;
  reg  line_719_valid_reg;
  reg [63:0] wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  wire  line_720_clock;
  wire  line_720_reset;
  wire  line_720_valid;
  reg  line_720_valid_reg;
  reg [7:0] wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  wire  line_721_clock;
  wire  line_721_reset;
  wire  line_721_valid;
  reg  line_721_valid_reg;
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire  line_722_clock;
  wire  line_722_reset;
  wire  line_722_valid;
  reg  line_722_valid_reg;
  reg [3:0] mmiocmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  wire  line_723_clock;
  wire  line_723_reset;
  wire  line_723_valid;
  reg  line_723_valid_reg;
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire  line_724_clock;
  wire  line_724_reset;
  wire  line_724_valid;
  reg  line_724_valid_reg;
  reg [3:0] memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  wire  line_725_clock;
  wire  line_725_reset;
  wire  line_725_valid;
  reg  line_725_valid_reg;
  wire  line_726_clock;
  wire  line_726_reset;
  wire  line_726_valid;
  reg  line_726_valid_reg;
  GEN_w1_line #(.COVER_INDEX(698)) line_698 (
    .clock(line_698_clock),
    .reset(line_698_reset),
    .valid(line_698_valid)
  );
  GEN_w1_line #(.COVER_INDEX(699)) line_699 (
    .clock(line_699_clock),
    .reset(line_699_reset),
    .valid(line_699_valid)
  );
  GEN_w1_line #(.COVER_INDEX(700)) line_700 (
    .clock(line_700_clock),
    .reset(line_700_reset),
    .valid(line_700_valid)
  );
  GEN_w1_line #(.COVER_INDEX(701)) line_701 (
    .clock(line_701_clock),
    .reset(line_701_reset),
    .valid(line_701_valid)
  );
  GEN_w1_line #(.COVER_INDEX(702)) line_702 (
    .clock(line_702_clock),
    .reset(line_702_reset),
    .valid(line_702_valid)
  );
  GEN_w1_line #(.COVER_INDEX(703)) line_703 (
    .clock(line_703_clock),
    .reset(line_703_reset),
    .valid(line_703_valid)
  );
  GEN_w1_line #(.COVER_INDEX(704)) line_704 (
    .clock(line_704_clock),
    .reset(line_704_reset),
    .valid(line_704_valid)
  );
  GEN_w1_line #(.COVER_INDEX(705)) line_705 (
    .clock(line_705_clock),
    .reset(line_705_reset),
    .valid(line_705_valid)
  );
  GEN_w1_line #(.COVER_INDEX(706)) line_706 (
    .clock(line_706_clock),
    .reset(line_706_reset),
    .valid(line_706_valid)
  );
  GEN_w1_line #(.COVER_INDEX(707)) line_707 (
    .clock(line_707_clock),
    .reset(line_707_reset),
    .valid(line_707_valid)
  );
  GEN_w1_line #(.COVER_INDEX(708)) line_708 (
    .clock(line_708_clock),
    .reset(line_708_reset),
    .valid(line_708_valid)
  );
  GEN_w1_line #(.COVER_INDEX(709)) line_709 (
    .clock(line_709_clock),
    .reset(line_709_reset),
    .valid(line_709_valid)
  );
  GEN_w1_line #(.COVER_INDEX(710)) line_710 (
    .clock(line_710_clock),
    .reset(line_710_reset),
    .valid(line_710_valid)
  );
  GEN_w1_line #(.COVER_INDEX(711)) line_711 (
    .clock(line_711_clock),
    .reset(line_711_reset),
    .valid(line_711_valid)
  );
  GEN_w1_line #(.COVER_INDEX(712)) line_712 (
    .clock(line_712_clock),
    .reset(line_712_reset),
    .valid(line_712_valid)
  );
  GEN_w1_line #(.COVER_INDEX(713)) line_713 (
    .clock(line_713_clock),
    .reset(line_713_reset),
    .valid(line_713_valid)
  );
  GEN_w1_line #(.COVER_INDEX(714)) line_714 (
    .clock(line_714_clock),
    .reset(line_714_reset),
    .valid(line_714_valid)
  );
  GEN_w1_line #(.COVER_INDEX(715)) line_715 (
    .clock(line_715_clock),
    .reset(line_715_reset),
    .valid(line_715_valid)
  );
  GEN_w1_line #(.COVER_INDEX(716)) line_716 (
    .clock(line_716_clock),
    .reset(line_716_reset),
    .valid(line_716_valid)
  );
  GEN_w1_line #(.COVER_INDEX(717)) line_717 (
    .clock(line_717_clock),
    .reset(line_717_reset),
    .valid(line_717_valid)
  );
  GEN_w1_line #(.COVER_INDEX(718)) line_718 (
    .clock(line_718_clock),
    .reset(line_718_reset),
    .valid(line_718_valid)
  );
  GEN_w1_line #(.COVER_INDEX(719)) line_719 (
    .clock(line_719_clock),
    .reset(line_719_reset),
    .valid(line_719_valid)
  );
  GEN_w1_line #(.COVER_INDEX(720)) line_720 (
    .clock(line_720_clock),
    .reset(line_720_reset),
    .valid(line_720_valid)
  );
  GEN_w1_line #(.COVER_INDEX(721)) line_721 (
    .clock(line_721_clock),
    .reset(line_721_reset),
    .valid(line_721_valid)
  );
  GEN_w1_line #(.COVER_INDEX(722)) line_722 (
    .clock(line_722_clock),
    .reset(line_722_reset),
    .valid(line_722_valid)
  );
  GEN_w1_line #(.COVER_INDEX(723)) line_723 (
    .clock(line_723_clock),
    .reset(line_723_reset),
    .valid(line_723_valid)
  );
  GEN_w1_line #(.COVER_INDEX(724)) line_724 (
    .clock(line_724_clock),
    .reset(line_724_reset),
    .valid(line_724_valid)
  );
  GEN_w1_line #(.COVER_INDEX(725)) line_725 (
    .clock(line_725_clock),
    .reset(line_725_reset),
    .valid(line_725_valid)
  );
  GEN_w1_line #(.COVER_INDEX(726)) line_726 (
    .clock(line_726_clock),
    .reset(line_726_reset),
    .valid(line_726_valid)
  );
  assign line_698_clock = clock;
  assign line_698_reset = reset;
  assign line_698_valid = _ismmioRec_T ^ line_698_valid_reg;
  assign line_699_clock = clock;
  assign line_699_reset = reset;
  assign line_699_valid = io_in_resp_valid ^ line_699_valid_reg;
  assign line_700_clock = clock;
  assign line_700_reset = reset;
  assign line_700_valid = _T_5 ^ line_700_valid_reg;
  assign line_701_clock = clock;
  assign line_701_reset = reset;
  assign line_701_valid = _ismmioRec_T ^ line_701_valid_reg;
  assign line_702_clock = clock;
  assign line_702_reset = reset;
  assign line_702_valid = _T_5 ^ line_702_valid_reg;
  assign line_703_clock = clock;
  assign line_703_reset = reset;
  assign line_703_valid = _T_10 ^ line_703_valid_reg;
  assign line_704_clock = clock;
  assign line_704_reset = reset;
  assign line_704_valid = _T_11 ^ line_704_valid_reg;
  assign line_705_clock = clock;
  assign line_705_reset = reset;
  assign line_705_valid = _T_10 ^ line_705_valid_reg;
  assign line_706_clock = clock;
  assign line_706_reset = reset;
  assign line_706_valid = _T_12 ^ line_706_valid_reg;
  assign line_707_clock = clock;
  assign line_707_reset = reset;
  assign line_707_valid = _T_13 ^ line_707_valid_reg;
  assign line_708_clock = clock;
  assign line_708_reset = reset;
  assign line_708_valid = _T_12 ^ line_708_valid_reg;
  assign line_709_clock = clock;
  assign line_709_reset = reset;
  assign line_709_valid = _T_14 ^ line_709_valid_reg;
  assign line_710_clock = clock;
  assign line_710_reset = reset;
  assign line_710_valid = _T_15 ^ line_710_valid_reg;
  assign line_711_clock = clock;
  assign line_711_reset = reset;
  assign line_711_valid = _T_14 ^ line_711_valid_reg;
  assign line_712_clock = clock;
  assign line_712_reset = reset;
  assign line_712_valid = _T_16 ^ line_712_valid_reg;
  assign line_713_clock = clock;
  assign line_713_reset = reset;
  assign line_713_valid = _T_18 ^ line_713_valid_reg;
  assign line_714_clock = clock;
  assign line_714_reset = reset;
  assign line_714_valid = _T_16 ^ line_714_valid_reg;
  assign line_715_clock = clock;
  assign line_715_reset = reset;
  assign line_715_valid = _T_19 ^ line_715_valid_reg;
  assign line_716_clock = clock;
  assign line_716_reset = reset;
  assign line_716_valid = _GEN_34 ^ line_716_valid_reg;
  assign line_717_clock = clock;
  assign line_717_reset = reset;
  assign line_717_valid = _ismmioRec_T ^ line_717_valid_reg;
  assign line_718_clock = clock;
  assign line_718_reset = reset;
  assign line_718_valid = _ismmioRec_T ^ line_718_valid_reg;
  assign line_719_clock = clock;
  assign line_719_reset = reset;
  assign line_719_valid = _ismmioRec_T ^ line_719_valid_reg;
  assign line_720_clock = clock;
  assign line_720_reset = reset;
  assign line_720_valid = _ismmioRec_T ^ line_720_valid_reg;
  assign line_721_clock = clock;
  assign line_721_reset = reset;
  assign line_721_valid = _ismmioRec_T ^ line_721_valid_reg;
  assign line_722_clock = clock;
  assign line_722_reset = reset;
  assign line_722_valid = _T_17 ^ line_722_valid_reg;
  assign line_723_clock = clock;
  assign line_723_reset = reset;
  assign line_723_valid = _T_17 ^ line_723_valid_reg;
  assign line_724_clock = clock;
  assign line_724_reset = reset;
  assign line_724_valid = _T_13 ^ line_724_valid_reg;
  assign line_725_clock = clock;
  assign line_725_reset = reset;
  assign line_725_valid = _T_13 ^ line_725_valid_reg;
  assign line_726_clock = clock;
  assign line_726_reset = reset;
  assign line_726_valid = _ismmioRec_T ^ line_726_valid_reg;
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5; // @[src/main/scala/nutcore/mem/Cache.scala 601:30]
  assign io_in_resp_bits_cmd = ismmioRec ? mmiocmd : memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 609:29]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_out_mem_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_out_mem_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_out_mem_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mmio_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mmio_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  assign ismmio_0 = ismmio;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_37;
    end else begin
      state <= _GEN_43;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    line_698_valid_reg <= _ismmioRec_T;
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_34;
    end
    line_699_valid_reg <= io_in_resp_valid;
    line_700_valid_reg <= _T_5;
    line_701_valid_reg <= _ismmioRec_T;
    line_702_valid_reg <= _T_5;
    line_703_valid_reg <= _T_10;
    line_704_valid_reg <= _T_11;
    line_705_valid_reg <= _T_10;
    line_706_valid_reg <= _T_12;
    line_707_valid_reg <= _T_13;
    line_708_valid_reg <= _T_12;
    line_709_valid_reg <= _T_14;
    line_710_valid_reg <= _T_15;
    line_711_valid_reg <= _T_14;
    line_712_valid_reg <= _T_16;
    line_713_valid_reg <= _T_18;
    line_714_valid_reg <= _T_16;
    line_715_valid_reg <= _T_19;
    line_716_valid_reg <= _GEN_34;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    line_717_valid_reg <= _ismmioRec_T;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
      cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    line_718_valid_reg <= _ismmioRec_T;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
      size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    line_719_valid_reg <= _ismmioRec_T;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
      wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    line_720_valid_reg <= _ismmioRec_T;
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
      wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    line_721_valid_reg <= _ismmioRec_T;
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    line_722_valid_reg <= _T_17;
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
      mmiocmd <= io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    line_723_valid_reg <= _T_17;
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    line_724_valid_reg <= _T_13;
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
      memcmd <= io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
    line_725_valid_reg <= _T_13;
    line_726_valid_reg <= _ismmioRec_T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_698_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alreadyOutFire = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_699_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_700_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_701_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_702_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_703_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_704_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_705_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_706_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_707_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_708_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_709_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_710_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_711_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_712_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_713_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_714_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_715_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_716_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  reqaddr = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  line_717_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  cmd = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  line_718_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  size = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  line_719_valid_reg = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  wdata = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  line_720_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  wmask = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  line_721_valid_reg = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  mmiordata = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  line_722_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  mmiocmd = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  line_723_valid_reg = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  memrdata = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  line_724_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  memcmd = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  line_725_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_726_valid_reg = _RAND_40[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (io_in_resp_valid) begin
      cover(1'h1);
    end
    //
    if (_T_5) begin
      cover(1'h1);
    end
    //
    if (_T_5 & _ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (~_T_5) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & _T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & _T_10 & _T_11) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & _T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & _T_12 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & _T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & _T_14 & _T_15) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & _T_16) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & _T_16 & _T_18) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16 & _T_19) begin
      cover(1'h1);
    end
    //
    if (~_T_5 & ~_T_10 & ~_T_12 & ~_T_14 & ~_T_16 & _T_19 & _GEN_34) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
    //
    if (_T_17) begin
      cover(1'h1);
    end
    //
    if (_T_17) begin
      cover(1'h1);
    end
    //
    if (_T_13) begin
      cover(1'h1);
    end
    //
    if (_T_13) begin
      cover(1'h1);
    end
    //
    if (_ismmioRec_T) begin
      cover(1'h1);
    end
  end
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_imem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_imem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_imem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_imem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_dmem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_dmem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [2:0]  io_dmem_mem_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_dmem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_dmem_mem_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_dmem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_dmem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_dmem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_frontend_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_extra_meip_0,
  output        isWFI,
  input         io_extra_mtip,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_reset; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_flushVec; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [1:0] frontend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_isWFI; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [11:0] frontend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  backend_clock; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_reset; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_flush; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_laf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_saf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_lr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_meip_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scInflight; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_actualTaken; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_amoReq; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_lrAddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [55:0] backend_paddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_satp; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scIsSuccess; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_mtip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_vmEnable; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [11:0] backend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_tlbFinish; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_ismmio; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_13_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_msip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  mmioXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  dmemXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_2_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_2_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  itlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] itlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_imem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [1:0] io_imem_cache_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  dtlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] dtlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_lr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_amoReq; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_lrAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [55:0] dtlb_paddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_12_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_vmEnable_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_tlbFinish_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_13_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_1_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_dmem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_ismmio_0; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  reg [63:0] dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [1:0] ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  reg [1:0] ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] _ringBufferAllowin_T_1 = ringBufferHead + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire [1:0] _ringBufferAllowin_T_4 = ringBufferHead + 2'h2; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire  ringBufferAllowin = _ringBufferAllowin_T_1 != ringBufferTail & _ringBufferAllowin_T_4 != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 33:124]
  wire  needEnqueue_0 = frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 36:27 37:20]
  wire [1:0] enqueueSize = {{1'd0}, needEnqueue_0}; // @[src/main/scala/utils/PipelineVector.scala 40:44]
  wire  enqueueFire_0 = enqueueSize >= 2'h1; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  enqueueFire_1 = enqueueSize >= 2'h2; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  wen = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_727_clock;
  wire  line_727_reset;
  wire  line_727_valid;
  reg  line_727_valid_reg;
  wire  line_728_clock;
  wire  line_728_reset;
  wire  line_728_valid;
  reg  line_728_valid_reg;
  wire [2:0] _T_1 = {{1'd0}, ringBufferHead}; // @[src/main/scala/utils/PipelineVector.scala 45:45]
  wire [63:0] _dataBuffer_T_cf_instr = needEnqueue_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pnpc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [3:0] _dataBuffer_T_cf_brIdx = needEnqueue_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [2:0] _dataBuffer_T_ctrl_fuType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [6:0] _dataBuffer_T_ctrl_fuOpType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc1 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc2 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfDest = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _dataBuffer_T_data_imm = needEnqueue_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire  _GEN_0 = 2'h0 == _T_1[1:0]; // @[src/main/scala/utils/PipelineVector.scala 45:63]
  wire  line_729_clock;
  wire  line_729_reset;
  wire  line_729_valid;
  reg  line_729_valid_reg;
  wire [63:0] _GEN_901 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_1 = 2'h1 == _T_1[1:0]; // @[src/main/scala/utils/PipelineVector.scala 45:63]
  wire  line_730_clock;
  wire  line_730_reset;
  wire  line_730_valid;
  reg  line_730_valid_reg;
  wire [63:0] _GEN_902 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_2 = 2'h2 == _T_1[1:0]; // @[src/main/scala/utils/PipelineVector.scala 45:63]
  wire  line_731_clock;
  wire  line_731_reset;
  wire  line_731_valid;
  reg  line_731_valid_reg;
  wire [63:0] _GEN_903 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_3 = 2'h3 == _T_1[1:0]; // @[src/main/scala/utils/PipelineVector.scala 45:63]
  wire  line_732_clock;
  wire  line_732_reset;
  wire  line_732_valid;
  reg  line_732_valid_reg;
  wire [63:0] _GEN_904 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_733_clock;
  wire  line_733_reset;
  wire  line_733_valid;
  reg  line_733_valid_reg;
  wire [38:0] _GEN_905 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_734_clock;
  wire  line_734_reset;
  wire  line_734_valid;
  reg  line_734_valid_reg;
  wire [38:0] _GEN_906 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_735_clock;
  wire  line_735_reset;
  wire  line_735_valid;
  reg  line_735_valid_reg;
  wire [38:0] _GEN_907 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_736_clock;
  wire  line_736_reset;
  wire  line_736_valid;
  reg  line_736_valid_reg;
  wire [38:0] _GEN_908 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_737_clock;
  wire  line_737_reset;
  wire  line_737_valid;
  reg  line_737_valid_reg;
  wire [38:0] _GEN_909 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_738_clock;
  wire  line_738_reset;
  wire  line_738_valid;
  reg  line_738_valid_reg;
  wire [38:0] _GEN_910 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_739_clock;
  wire  line_739_reset;
  wire  line_739_valid;
  reg  line_739_valid_reg;
  wire [38:0] _GEN_911 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_740_clock;
  wire  line_740_reset;
  wire  line_740_valid;
  reg  line_740_valid_reg;
  wire [38:0] _GEN_912 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_741_clock;
  wire  line_741_reset;
  wire  line_741_valid;
  reg  line_741_valid_reg;
  wire  line_742_clock;
  wire  line_742_reset;
  wire  line_742_valid;
  reg  line_742_valid_reg;
  wire  line_743_clock;
  wire  line_743_reset;
  wire  line_743_valid;
  reg  line_743_valid_reg;
  wire  line_744_clock;
  wire  line_744_reset;
  wire  line_744_valid;
  reg  line_744_valid_reg;
  wire  line_745_clock;
  wire  line_745_reset;
  wire  line_745_valid;
  reg  line_745_valid_reg;
  wire  line_746_clock;
  wire  line_746_reset;
  wire  line_746_valid;
  reg  line_746_valid_reg;
  wire  line_747_clock;
  wire  line_747_reset;
  wire  line_747_valid;
  reg  line_747_valid_reg;
  wire  line_748_clock;
  wire  line_748_reset;
  wire  line_748_valid;
  reg  line_748_valid_reg;
  wire  line_749_clock;
  wire  line_749_reset;
  wire  line_749_valid;
  reg  line_749_valid_reg;
  wire  line_750_clock;
  wire  line_750_reset;
  wire  line_750_valid;
  reg  line_750_valid_reg;
  wire  line_751_clock;
  wire  line_751_reset;
  wire  line_751_valid;
  reg  line_751_valid_reg;
  wire  line_752_clock;
  wire  line_752_reset;
  wire  line_752_valid;
  reg  line_752_valid_reg;
  wire  line_753_clock;
  wire  line_753_reset;
  wire  line_753_valid;
  reg  line_753_valid_reg;
  wire  line_754_clock;
  wire  line_754_reset;
  wire  line_754_valid;
  reg  line_754_valid_reg;
  wire  line_755_clock;
  wire  line_755_reset;
  wire  line_755_valid;
  reg  line_755_valid_reg;
  wire  line_756_clock;
  wire  line_756_reset;
  wire  line_756_valid;
  reg  line_756_valid_reg;
  wire  line_757_clock;
  wire  line_757_reset;
  wire  line_757_valid;
  reg  line_757_valid_reg;
  wire  _GEN_929 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_758_clock;
  wire  line_758_reset;
  wire  line_758_valid;
  reg  line_758_valid_reg;
  wire  _GEN_930 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_759_clock;
  wire  line_759_reset;
  wire  line_759_valid;
  reg  line_759_valid_reg;
  wire  _GEN_931 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_760_clock;
  wire  line_760_reset;
  wire  line_760_valid;
  reg  line_760_valid_reg;
  wire  _GEN_932 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_761_clock;
  wire  line_761_reset;
  wire  line_761_valid;
  reg  line_761_valid_reg;
  wire  _GEN_933 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_762_clock;
  wire  line_762_reset;
  wire  line_762_valid;
  reg  line_762_valid_reg;
  wire  _GEN_934 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_763_clock;
  wire  line_763_reset;
  wire  line_763_valid;
  reg  line_763_valid_reg;
  wire  _GEN_935 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_764_clock;
  wire  line_764_reset;
  wire  line_764_valid;
  reg  line_764_valid_reg;
  wire  _GEN_936 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_765_clock;
  wire  line_765_reset;
  wire  line_765_valid;
  reg  line_765_valid_reg;
  wire  line_766_clock;
  wire  line_766_reset;
  wire  line_766_valid;
  reg  line_766_valid_reg;
  wire  line_767_clock;
  wire  line_767_reset;
  wire  line_767_valid;
  reg  line_767_valid_reg;
  wire  line_768_clock;
  wire  line_768_reset;
  wire  line_768_valid;
  reg  line_768_valid_reg;
  wire  line_769_clock;
  wire  line_769_reset;
  wire  line_769_valid;
  reg  line_769_valid_reg;
  wire  line_770_clock;
  wire  line_770_reset;
  wire  line_770_valid;
  reg  line_770_valid_reg;
  wire  line_771_clock;
  wire  line_771_reset;
  wire  line_771_valid;
  reg  line_771_valid_reg;
  wire  line_772_clock;
  wire  line_772_reset;
  wire  line_772_valid;
  reg  line_772_valid_reg;
  wire  line_773_clock;
  wire  line_773_reset;
  wire  line_773_valid;
  reg  line_773_valid_reg;
  wire  line_774_clock;
  wire  line_774_reset;
  wire  line_774_valid;
  reg  line_774_valid_reg;
  wire  line_775_clock;
  wire  line_775_reset;
  wire  line_775_valid;
  reg  line_775_valid_reg;
  wire  line_776_clock;
  wire  line_776_reset;
  wire  line_776_valid;
  reg  line_776_valid_reg;
  wire  line_777_clock;
  wire  line_777_reset;
  wire  line_777_valid;
  reg  line_777_valid_reg;
  wire  line_778_clock;
  wire  line_778_reset;
  wire  line_778_valid;
  reg  line_778_valid_reg;
  wire  line_779_clock;
  wire  line_779_reset;
  wire  line_779_valid;
  reg  line_779_valid_reg;
  wire  line_780_clock;
  wire  line_780_reset;
  wire  line_780_valid;
  reg  line_780_valid_reg;
  wire  line_781_clock;
  wire  line_781_reset;
  wire  line_781_valid;
  reg  line_781_valid_reg;
  wire  line_782_clock;
  wire  line_782_reset;
  wire  line_782_valid;
  reg  line_782_valid_reg;
  wire  line_783_clock;
  wire  line_783_reset;
  wire  line_783_valid;
  reg  line_783_valid_reg;
  wire  line_784_clock;
  wire  line_784_reset;
  wire  line_784_valid;
  reg  line_784_valid_reg;
  wire  line_785_clock;
  wire  line_785_reset;
  wire  line_785_valid;
  reg  line_785_valid_reg;
  wire  line_786_clock;
  wire  line_786_reset;
  wire  line_786_valid;
  reg  line_786_valid_reg;
  wire  line_787_clock;
  wire  line_787_reset;
  wire  line_787_valid;
  reg  line_787_valid_reg;
  wire  line_788_clock;
  wire  line_788_reset;
  wire  line_788_valid;
  reg  line_788_valid_reg;
  wire  line_789_clock;
  wire  line_789_reset;
  wire  line_789_valid;
  reg  line_789_valid_reg;
  wire  line_790_clock;
  wire  line_790_reset;
  wire  line_790_valid;
  reg  line_790_valid_reg;
  wire  line_791_clock;
  wire  line_791_reset;
  wire  line_791_valid;
  reg  line_791_valid_reg;
  wire  line_792_clock;
  wire  line_792_reset;
  wire  line_792_valid;
  reg  line_792_valid_reg;
  wire  line_793_clock;
  wire  line_793_reset;
  wire  line_793_valid;
  reg  line_793_valid_reg;
  wire  line_794_clock;
  wire  line_794_reset;
  wire  line_794_valid;
  reg  line_794_valid_reg;
  wire  line_795_clock;
  wire  line_795_reset;
  wire  line_795_valid;
  reg  line_795_valid_reg;
  wire  line_796_clock;
  wire  line_796_reset;
  wire  line_796_valid;
  reg  line_796_valid_reg;
  wire  line_797_clock;
  wire  line_797_reset;
  wire  line_797_valid;
  reg  line_797_valid_reg;
  wire  line_798_clock;
  wire  line_798_reset;
  wire  line_798_valid;
  reg  line_798_valid_reg;
  wire  line_799_clock;
  wire  line_799_reset;
  wire  line_799_valid;
  reg  line_799_valid_reg;
  wire  line_800_clock;
  wire  line_800_reset;
  wire  line_800_valid;
  reg  line_800_valid_reg;
  wire  line_801_clock;
  wire  line_801_reset;
  wire  line_801_valid;
  reg  line_801_valid_reg;
  wire  _GEN_973 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_802_clock;
  wire  line_802_reset;
  wire  line_802_valid;
  reg  line_802_valid_reg;
  wire  _GEN_974 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_803_clock;
  wire  line_803_reset;
  wire  line_803_valid;
  reg  line_803_valid_reg;
  wire  _GEN_975 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_804_clock;
  wire  line_804_reset;
  wire  line_804_valid;
  reg  line_804_valid_reg;
  wire  _GEN_976 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_805_clock;
  wire  line_805_reset;
  wire  line_805_valid;
  reg  line_805_valid_reg;
  wire  line_806_clock;
  wire  line_806_reset;
  wire  line_806_valid;
  reg  line_806_valid_reg;
  wire  line_807_clock;
  wire  line_807_reset;
  wire  line_807_valid;
  reg  line_807_valid_reg;
  wire  line_808_clock;
  wire  line_808_reset;
  wire  line_808_valid;
  reg  line_808_valid_reg;
  wire  line_809_clock;
  wire  line_809_reset;
  wire  line_809_valid;
  reg  line_809_valid_reg;
  wire  line_810_clock;
  wire  line_810_reset;
  wire  line_810_valid;
  reg  line_810_valid_reg;
  wire  line_811_clock;
  wire  line_811_reset;
  wire  line_811_valid;
  reg  line_811_valid_reg;
  wire  line_812_clock;
  wire  line_812_reset;
  wire  line_812_valid;
  reg  line_812_valid_reg;
  wire  line_813_clock;
  wire  line_813_reset;
  wire  line_813_valid;
  reg  line_813_valid_reg;
  wire  line_814_clock;
  wire  line_814_reset;
  wire  line_814_valid;
  reg  line_814_valid_reg;
  wire  line_815_clock;
  wire  line_815_reset;
  wire  line_815_valid;
  reg  line_815_valid_reg;
  wire  line_816_clock;
  wire  line_816_reset;
  wire  line_816_valid;
  reg  line_816_valid_reg;
  wire  line_817_clock;
  wire  line_817_reset;
  wire  line_817_valid;
  reg  line_817_valid_reg;
  wire  line_818_clock;
  wire  line_818_reset;
  wire  line_818_valid;
  reg  line_818_valid_reg;
  wire  line_819_clock;
  wire  line_819_reset;
  wire  line_819_valid;
  reg  line_819_valid_reg;
  wire  line_820_clock;
  wire  line_820_reset;
  wire  line_820_valid;
  reg  line_820_valid_reg;
  wire  line_821_clock;
  wire  line_821_reset;
  wire  line_821_valid;
  reg  line_821_valid_reg;
  wire  _GEN_993 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_822_clock;
  wire  line_822_reset;
  wire  line_822_valid;
  reg  line_822_valid_reg;
  wire  _GEN_994 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_823_clock;
  wire  line_823_reset;
  wire  line_823_valid;
  reg  line_823_valid_reg;
  wire  _GEN_995 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_824_clock;
  wire  line_824_reset;
  wire  line_824_valid;
  reg  line_824_valid_reg;
  wire  _GEN_996 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_825_clock;
  wire  line_825_reset;
  wire  line_825_valid;
  reg  line_825_valid_reg;
  wire  line_826_clock;
  wire  line_826_reset;
  wire  line_826_valid;
  reg  line_826_valid_reg;
  wire  line_827_clock;
  wire  line_827_reset;
  wire  line_827_valid;
  reg  line_827_valid_reg;
  wire  line_828_clock;
  wire  line_828_reset;
  wire  line_828_valid;
  reg  line_828_valid_reg;
  wire  line_829_clock;
  wire  line_829_reset;
  wire  line_829_valid;
  reg  line_829_valid_reg;
  wire  _GEN_1001 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_830_clock;
  wire  line_830_reset;
  wire  line_830_valid;
  reg  line_830_valid_reg;
  wire  _GEN_1002 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_831_clock;
  wire  line_831_reset;
  wire  line_831_valid;
  reg  line_831_valid_reg;
  wire  _GEN_1003 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_832_clock;
  wire  line_832_reset;
  wire  line_832_valid;
  reg  line_832_valid_reg;
  wire  _GEN_1004 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_833_clock;
  wire  line_833_reset;
  wire  line_833_valid;
  reg  line_833_valid_reg;
  wire  line_834_clock;
  wire  line_834_reset;
  wire  line_834_valid;
  reg  line_834_valid_reg;
  wire  line_835_clock;
  wire  line_835_reset;
  wire  line_835_valid;
  reg  line_835_valid_reg;
  wire  line_836_clock;
  wire  line_836_reset;
  wire  line_836_valid;
  reg  line_836_valid_reg;
  wire  line_837_clock;
  wire  line_837_reset;
  wire  line_837_valid;
  reg  line_837_valid_reg;
  wire  _GEN_1009 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_838_clock;
  wire  line_838_reset;
  wire  line_838_valid;
  reg  line_838_valid_reg;
  wire  _GEN_1010 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_839_clock;
  wire  line_839_reset;
  wire  line_839_valid;
  reg  line_839_valid_reg;
  wire  _GEN_1011 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_840_clock;
  wire  line_840_reset;
  wire  line_840_valid;
  reg  line_840_valid_reg;
  wire  _GEN_1012 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_841_clock;
  wire  line_841_reset;
  wire  line_841_valid;
  reg  line_841_valid_reg;
  wire  line_842_clock;
  wire  line_842_reset;
  wire  line_842_valid;
  reg  line_842_valid_reg;
  wire  line_843_clock;
  wire  line_843_reset;
  wire  line_843_valid;
  reg  line_843_valid_reg;
  wire  line_844_clock;
  wire  line_844_reset;
  wire  line_844_valid;
  reg  line_844_valid_reg;
  wire  line_845_clock;
  wire  line_845_reset;
  wire  line_845_valid;
  reg  line_845_valid_reg;
  wire  _GEN_1017 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_846_clock;
  wire  line_846_reset;
  wire  line_846_valid;
  reg  line_846_valid_reg;
  wire  _GEN_1018 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_847_clock;
  wire  line_847_reset;
  wire  line_847_valid;
  reg  line_847_valid_reg;
  wire  _GEN_1019 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_848_clock;
  wire  line_848_reset;
  wire  line_848_valid;
  reg  line_848_valid_reg;
  wire  _GEN_1020 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_849_clock;
  wire  line_849_reset;
  wire  line_849_valid;
  reg  line_849_valid_reg;
  wire  line_850_clock;
  wire  line_850_reset;
  wire  line_850_valid;
  reg  line_850_valid_reg;
  wire  line_851_clock;
  wire  line_851_reset;
  wire  line_851_valid;
  reg  line_851_valid_reg;
  wire  line_852_clock;
  wire  line_852_reset;
  wire  line_852_valid;
  reg  line_852_valid_reg;
  wire  line_853_clock;
  wire  line_853_reset;
  wire  line_853_valid;
  reg  line_853_valid_reg;
  wire  _GEN_1025 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_854_clock;
  wire  line_854_reset;
  wire  line_854_valid;
  reg  line_854_valid_reg;
  wire  _GEN_1026 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_855_clock;
  wire  line_855_reset;
  wire  line_855_valid;
  reg  line_855_valid_reg;
  wire  _GEN_1027 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_856_clock;
  wire  line_856_reset;
  wire  line_856_valid;
  reg  line_856_valid_reg;
  wire  _GEN_1028 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_857_clock;
  wire  line_857_reset;
  wire  line_857_valid;
  reg  line_857_valid_reg;
  wire  line_858_clock;
  wire  line_858_reset;
  wire  line_858_valid;
  reg  line_858_valid_reg;
  wire  line_859_clock;
  wire  line_859_reset;
  wire  line_859_valid;
  reg  line_859_valid_reg;
  wire  line_860_clock;
  wire  line_860_reset;
  wire  line_860_valid;
  reg  line_860_valid_reg;
  wire  line_861_clock;
  wire  line_861_reset;
  wire  line_861_valid;
  reg  line_861_valid_reg;
  wire  _GEN_1033 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 :
    dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_862_clock;
  wire  line_862_reset;
  wire  line_862_valid;
  reg  line_862_valid_reg;
  wire  _GEN_1034 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 :
    dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_863_clock;
  wire  line_863_reset;
  wire  line_863_valid;
  reg  line_863_valid_reg;
  wire  _GEN_1035 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 :
    dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_864_clock;
  wire  line_864_reset;
  wire  line_864_valid;
  reg  line_864_valid_reg;
  wire  _GEN_1036 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 :
    dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_865_clock;
  wire  line_865_reset;
  wire  line_865_valid;
  reg  line_865_valid_reg;
  wire [3:0] _GEN_1037 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_866_clock;
  wire  line_866_reset;
  wire  line_866_valid;
  reg  line_866_valid_reg;
  wire [3:0] _GEN_1038 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_867_clock;
  wire  line_867_reset;
  wire  line_867_valid;
  reg  line_867_valid_reg;
  wire [3:0] _GEN_1039 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_868_clock;
  wire  line_868_reset;
  wire  line_868_valid;
  reg  line_868_valid_reg;
  wire [3:0] _GEN_1040 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_869_clock;
  wire  line_869_reset;
  wire  line_869_valid;
  reg  line_869_valid_reg;
  wire  line_870_clock;
  wire  line_870_reset;
  wire  line_870_valid;
  reg  line_870_valid_reg;
  wire  line_871_clock;
  wire  line_871_reset;
  wire  line_871_valid;
  reg  line_871_valid_reg;
  wire  line_872_clock;
  wire  line_872_reset;
  wire  line_872_valid;
  reg  line_872_valid_reg;
  wire  line_873_clock;
  wire  line_873_reset;
  wire  line_873_valid;
  reg  line_873_valid_reg;
  wire  _GEN_1045 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_874_clock;
  wire  line_874_reset;
  wire  line_874_valid;
  reg  line_874_valid_reg;
  wire  _GEN_1046 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_875_clock;
  wire  line_875_reset;
  wire  line_875_valid;
  reg  line_875_valid_reg;
  wire  _GEN_1047 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_876_clock;
  wire  line_876_reset;
  wire  line_876_valid;
  reg  line_876_valid_reg;
  wire  _GEN_1048 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_877_clock;
  wire  line_877_reset;
  wire  line_877_valid;
  reg  line_877_valid_reg;
  wire  line_878_clock;
  wire  line_878_reset;
  wire  line_878_valid;
  reg  line_878_valid_reg;
  wire  line_879_clock;
  wire  line_879_reset;
  wire  line_879_valid;
  reg  line_879_valid_reg;
  wire  line_880_clock;
  wire  line_880_reset;
  wire  line_880_valid;
  reg  line_880_valid_reg;
  wire  line_881_clock;
  wire  line_881_reset;
  wire  line_881_valid;
  reg  line_881_valid_reg;
  wire  line_882_clock;
  wire  line_882_reset;
  wire  line_882_valid;
  reg  line_882_valid_reg;
  wire  line_883_clock;
  wire  line_883_reset;
  wire  line_883_valid;
  reg  line_883_valid_reg;
  wire  line_884_clock;
  wire  line_884_reset;
  wire  line_884_valid;
  reg  line_884_valid_reg;
  wire  line_885_clock;
  wire  line_885_reset;
  wire  line_885_valid;
  reg  line_885_valid_reg;
  wire  line_886_clock;
  wire  line_886_reset;
  wire  line_886_valid;
  reg  line_886_valid_reg;
  wire  line_887_clock;
  wire  line_887_reset;
  wire  line_887_valid;
  reg  line_887_valid_reg;
  wire  line_888_clock;
  wire  line_888_reset;
  wire  line_888_valid;
  reg  line_888_valid_reg;
  wire  line_889_clock;
  wire  line_889_reset;
  wire  line_889_valid;
  reg  line_889_valid_reg;
  wire  _GEN_1061 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type :
    dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_890_clock;
  wire  line_890_reset;
  wire  line_890_valid;
  reg  line_890_valid_reg;
  wire  _GEN_1062 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type :
    dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_891_clock;
  wire  line_891_reset;
  wire  line_891_valid;
  reg  line_891_valid_reg;
  wire  _GEN_1063 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type :
    dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_892_clock;
  wire  line_892_reset;
  wire  line_892_valid;
  reg  line_892_valid_reg;
  wire  _GEN_1064 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type :
    dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_893_clock;
  wire  line_893_reset;
  wire  line_893_valid;
  reg  line_893_valid_reg;
  wire  _GEN_1065 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type :
    dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_894_clock;
  wire  line_894_reset;
  wire  line_894_valid;
  reg  line_894_valid_reg;
  wire  _GEN_1066 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type :
    dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_895_clock;
  wire  line_895_reset;
  wire  line_895_valid;
  reg  line_895_valid_reg;
  wire  _GEN_1067 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type :
    dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_896_clock;
  wire  line_896_reset;
  wire  line_896_valid;
  reg  line_896_valid_reg;
  wire  _GEN_1068 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type :
    dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_897_clock;
  wire  line_897_reset;
  wire  line_897_valid;
  reg  line_897_valid_reg;
  wire [2:0] _GEN_1069 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_898_clock;
  wire  line_898_reset;
  wire  line_898_valid;
  reg  line_898_valid_reg;
  wire [2:0] _GEN_1070 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_899_clock;
  wire  line_899_reset;
  wire  line_899_valid;
  reg  line_899_valid_reg;
  wire [2:0] _GEN_1071 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_900_clock;
  wire  line_900_reset;
  wire  line_900_valid;
  reg  line_900_valid_reg;
  wire [2:0] _GEN_1072 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_901_clock;
  wire  line_901_reset;
  wire  line_901_valid;
  reg  line_901_valid_reg;
  wire [6:0] _GEN_1073 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_902_clock;
  wire  line_902_reset;
  wire  line_902_valid;
  reg  line_902_valid_reg;
  wire [6:0] _GEN_1074 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_903_clock;
  wire  line_903_reset;
  wire  line_903_valid;
  reg  line_903_valid_reg;
  wire [6:0] _GEN_1075 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_904_clock;
  wire  line_904_reset;
  wire  line_904_valid;
  reg  line_904_valid_reg;
  wire [6:0] _GEN_1076 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_905_clock;
  wire  line_905_reset;
  wire  line_905_valid;
  reg  line_905_valid_reg;
  wire [4:0] _GEN_1077 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_906_clock;
  wire  line_906_reset;
  wire  line_906_valid;
  reg  line_906_valid_reg;
  wire [4:0] _GEN_1078 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_907_clock;
  wire  line_907_reset;
  wire  line_907_valid;
  reg  line_907_valid_reg;
  wire [4:0] _GEN_1079 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_908_clock;
  wire  line_908_reset;
  wire  line_908_valid;
  reg  line_908_valid_reg;
  wire [4:0] _GEN_1080 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_909_clock;
  wire  line_909_reset;
  wire  line_909_valid;
  reg  line_909_valid_reg;
  wire [4:0] _GEN_1081 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_910_clock;
  wire  line_910_reset;
  wire  line_910_valid;
  reg  line_910_valid_reg;
  wire [4:0] _GEN_1082 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_911_clock;
  wire  line_911_reset;
  wire  line_911_valid;
  reg  line_911_valid_reg;
  wire [4:0] _GEN_1083 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_912_clock;
  wire  line_912_reset;
  wire  line_912_valid;
  reg  line_912_valid_reg;
  wire [4:0] _GEN_1084 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_913_clock;
  wire  line_913_reset;
  wire  line_913_valid;
  reg  line_913_valid_reg;
  wire  _GEN_1085 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_914_clock;
  wire  line_914_reset;
  wire  line_914_valid;
  reg  line_914_valid_reg;
  wire  _GEN_1086 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_915_clock;
  wire  line_915_reset;
  wire  line_915_valid;
  reg  line_915_valid_reg;
  wire  _GEN_1087 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_916_clock;
  wire  line_916_reset;
  wire  line_916_valid;
  reg  line_916_valid_reg;
  wire  _GEN_1088 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_917_clock;
  wire  line_917_reset;
  wire  line_917_valid;
  reg  line_917_valid_reg;
  wire [4:0] _GEN_1089 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_918_clock;
  wire  line_918_reset;
  wire  line_918_valid;
  reg  line_918_valid_reg;
  wire [4:0] _GEN_1090 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_919_clock;
  wire  line_919_reset;
  wire  line_919_valid;
  reg  line_919_valid_reg;
  wire [4:0] _GEN_1091 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_920_clock;
  wire  line_920_reset;
  wire  line_920_valid;
  reg  line_920_valid_reg;
  wire [4:0] _GEN_1092 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_921_clock;
  wire  line_921_reset;
  wire  line_921_valid;
  reg  line_921_valid_reg;
  wire  _GEN_1093 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_922_clock;
  wire  line_922_reset;
  wire  line_922_valid;
  reg  line_922_valid_reg;
  wire  _GEN_1094 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_923_clock;
  wire  line_923_reset;
  wire  line_923_valid;
  reg  line_923_valid_reg;
  wire  _GEN_1095 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_924_clock;
  wire  line_924_reset;
  wire  line_924_valid;
  reg  line_924_valid_reg;
  wire  _GEN_1096 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_925_clock;
  wire  line_925_reset;
  wire  line_925_valid;
  reg  line_925_valid_reg;
  wire  line_926_clock;
  wire  line_926_reset;
  wire  line_926_valid;
  reg  line_926_valid_reg;
  wire  line_927_clock;
  wire  line_927_reset;
  wire  line_927_valid;
  reg  line_927_valid_reg;
  wire  line_928_clock;
  wire  line_928_reset;
  wire  line_928_valid;
  reg  line_928_valid_reg;
  wire  line_929_clock;
  wire  line_929_reset;
  wire  line_929_valid;
  reg  line_929_valid_reg;
  wire  line_930_clock;
  wire  line_930_reset;
  wire  line_930_valid;
  reg  line_930_valid_reg;
  wire  line_931_clock;
  wire  line_931_reset;
  wire  line_931_valid;
  reg  line_931_valid_reg;
  wire  line_932_clock;
  wire  line_932_reset;
  wire  line_932_valid;
  reg  line_932_valid_reg;
  wire  line_933_clock;
  wire  line_933_reset;
  wire  line_933_valid;
  reg  line_933_valid_reg;
  wire  line_934_clock;
  wire  line_934_reset;
  wire  line_934_valid;
  reg  line_934_valid_reg;
  wire  line_935_clock;
  wire  line_935_reset;
  wire  line_935_valid;
  reg  line_935_valid_reg;
  wire  line_936_clock;
  wire  line_936_reset;
  wire  line_936_valid;
  reg  line_936_valid_reg;
  wire  line_937_clock;
  wire  line_937_reset;
  wire  line_937_valid;
  reg  line_937_valid_reg;
  wire  line_938_clock;
  wire  line_938_reset;
  wire  line_938_valid;
  reg  line_938_valid_reg;
  wire  line_939_clock;
  wire  line_939_reset;
  wire  line_939_valid;
  reg  line_939_valid_reg;
  wire  line_940_clock;
  wire  line_940_reset;
  wire  line_940_valid;
  reg  line_940_valid_reg;
  wire  line_941_clock;
  wire  line_941_reset;
  wire  line_941_valid;
  reg  line_941_valid_reg;
  wire  line_942_clock;
  wire  line_942_reset;
  wire  line_942_valid;
  reg  line_942_valid_reg;
  wire  line_943_clock;
  wire  line_943_reset;
  wire  line_943_valid;
  reg  line_943_valid_reg;
  wire  line_944_clock;
  wire  line_944_reset;
  wire  line_944_valid;
  reg  line_944_valid_reg;
  wire  line_945_clock;
  wire  line_945_reset;
  wire  line_945_valid;
  reg  line_945_valid_reg;
  wire  line_946_clock;
  wire  line_946_reset;
  wire  line_946_valid;
  reg  line_946_valid_reg;
  wire  line_947_clock;
  wire  line_947_reset;
  wire  line_947_valid;
  reg  line_947_valid_reg;
  wire  line_948_clock;
  wire  line_948_reset;
  wire  line_948_valid;
  reg  line_948_valid_reg;
  wire  line_949_clock;
  wire  line_949_reset;
  wire  line_949_valid;
  reg  line_949_valid_reg;
  wire [63:0] _GEN_1121 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_950_clock;
  wire  line_950_reset;
  wire  line_950_valid;
  reg  line_950_valid_reg;
  wire [63:0] _GEN_1122 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_951_clock;
  wire  line_951_reset;
  wire  line_951_valid;
  reg  line_951_valid_reg;
  wire [63:0] _GEN_1123 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  line_952_clock;
  wire  line_952_reset;
  wire  line_952_valid;
  reg  line_952_valid_reg;
  wire [63:0] _GEN_1124 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1125 = enqueueFire_0 ? _GEN_901 : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1126 = enqueueFire_0 ? _GEN_902 : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1127 = enqueueFire_0 ? _GEN_903 : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1128 = enqueueFire_0 ? _GEN_904 : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1129 = enqueueFire_0 ? _GEN_905 : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1130 = enqueueFire_0 ? _GEN_906 : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1131 = enqueueFire_0 ? _GEN_907 : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1132 = enqueueFire_0 ? _GEN_908 : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1133 = enqueueFire_0 ? _GEN_909 : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1134 = enqueueFire_0 ? _GEN_910 : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1135 = enqueueFire_0 ? _GEN_911 : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_1136 = enqueueFire_0 ? _GEN_912 : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1153 = enqueueFire_0 ? _GEN_929 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1154 = enqueueFire_0 ? _GEN_930 : dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1155 = enqueueFire_0 ? _GEN_931 : dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1156 = enqueueFire_0 ? _GEN_932 : dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1157 = enqueueFire_0 ? _GEN_933 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1158 = enqueueFire_0 ? _GEN_934 : dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1159 = enqueueFire_0 ? _GEN_935 : dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1160 = enqueueFire_0 ? _GEN_936 : dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1197 = enqueueFire_0 ? _GEN_973 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1198 = enqueueFire_0 ? _GEN_974 : dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1199 = enqueueFire_0 ? _GEN_975 : dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1200 = enqueueFire_0 ? _GEN_976 : dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1217 = enqueueFire_0 ? _GEN_993 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1218 = enqueueFire_0 ? _GEN_994 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1219 = enqueueFire_0 ? _GEN_995 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1220 = enqueueFire_0 ? _GEN_996 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1225 = enqueueFire_0 ? _GEN_1001 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1226 = enqueueFire_0 ? _GEN_1002 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1227 = enqueueFire_0 ? _GEN_1003 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1228 = enqueueFire_0 ? _GEN_1004 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1233 = enqueueFire_0 ? _GEN_1009 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1234 = enqueueFire_0 ? _GEN_1010 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1235 = enqueueFire_0 ? _GEN_1011 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1236 = enqueueFire_0 ? _GEN_1012 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1241 = enqueueFire_0 ? _GEN_1017 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1242 = enqueueFire_0 ? _GEN_1018 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1243 = enqueueFire_0 ? _GEN_1019 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1244 = enqueueFire_0 ? _GEN_1020 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1249 = enqueueFire_0 ? _GEN_1025 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1250 = enqueueFire_0 ? _GEN_1026 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1251 = enqueueFire_0 ? _GEN_1027 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1252 = enqueueFire_0 ? _GEN_1028 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1257 = enqueueFire_0 ? _GEN_1033 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1258 = enqueueFire_0 ? _GEN_1034 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1259 = enqueueFire_0 ? _GEN_1035 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1260 = enqueueFire_0 ? _GEN_1036 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_1261 = enqueueFire_0 ? _GEN_1037 : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_1262 = enqueueFire_0 ? _GEN_1038 : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_1263 = enqueueFire_0 ? _GEN_1039 : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_1264 = enqueueFire_0 ? _GEN_1040 : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1269 = enqueueFire_0 ? _GEN_1045 : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1270 = enqueueFire_0 ? _GEN_1046 : dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1271 = enqueueFire_0 ? _GEN_1047 : dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1272 = enqueueFire_0 ? _GEN_1048 : dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1285 = enqueueFire_0 ? _GEN_1061 : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1286 = enqueueFire_0 ? _GEN_1062 : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1287 = enqueueFire_0 ? _GEN_1063 : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1288 = enqueueFire_0 ? _GEN_1064 : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1289 = enqueueFire_0 ? _GEN_1065 : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1290 = enqueueFire_0 ? _GEN_1066 : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1291 = enqueueFire_0 ? _GEN_1067 : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1292 = enqueueFire_0 ? _GEN_1068 : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_1293 = enqueueFire_0 ? _GEN_1069 : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_1294 = enqueueFire_0 ? _GEN_1070 : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_1295 = enqueueFire_0 ? _GEN_1071 : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_1296 = enqueueFire_0 ? _GEN_1072 : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_1297 = enqueueFire_0 ? _GEN_1073 : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_1298 = enqueueFire_0 ? _GEN_1074 : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_1299 = enqueueFire_0 ? _GEN_1075 : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_1300 = enqueueFire_0 ? _GEN_1076 : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1301 = enqueueFire_0 ? _GEN_1077 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1302 = enqueueFire_0 ? _GEN_1078 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1303 = enqueueFire_0 ? _GEN_1079 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1304 = enqueueFire_0 ? _GEN_1080 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1305 = enqueueFire_0 ? _GEN_1081 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1306 = enqueueFire_0 ? _GEN_1082 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1307 = enqueueFire_0 ? _GEN_1083 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1308 = enqueueFire_0 ? _GEN_1084 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1309 = enqueueFire_0 ? _GEN_1085 : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1310 = enqueueFire_0 ? _GEN_1086 : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1311 = enqueueFire_0 ? _GEN_1087 : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1312 = enqueueFire_0 ? _GEN_1088 : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1313 = enqueueFire_0 ? _GEN_1089 : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1314 = enqueueFire_0 ? _GEN_1090 : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1315 = enqueueFire_0 ? _GEN_1091 : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_1316 = enqueueFire_0 ? _GEN_1092 : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1317 = enqueueFire_0 ? _GEN_1093 : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1318 = enqueueFire_0 ? _GEN_1094 : dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1319 = enqueueFire_0 ? _GEN_1095 : dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_1320 = enqueueFire_0 ? _GEN_1096 : dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1345 = enqueueFire_0 ? _GEN_1121 : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1346 = enqueueFire_0 ? _GEN_1122 : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1347 = enqueueFire_0 ? _GEN_1123 : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_1348 = enqueueFire_0 ? _GEN_1124 : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  line_953_clock;
  wire  line_953_reset;
  wire  line_953_valid;
  reg  line_953_valid_reg;
  wire [1:0] _T_4 = 2'h1 + ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 46:45]
  wire  _GEN_225 = 2'h0 == _T_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
  wire  line_954_clock;
  wire  line_954_reset;
  wire  line_954_valid;
  reg  line_954_valid_reg;
  wire  _GEN_226 = 2'h1 == _T_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
  wire  line_955_clock;
  wire  line_955_reset;
  wire  line_955_valid;
  reg  line_955_valid_reg;
  wire  _GEN_227 = 2'h2 == _T_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
  wire  line_956_clock;
  wire  line_956_reset;
  wire  line_956_valid;
  reg  line_956_valid_reg;
  wire  _GEN_228 = 2'h3 == _T_4; // @[src/main/scala/utils/PipelineVector.scala 46:63]
  wire  line_957_clock;
  wire  line_957_reset;
  wire  line_957_valid;
  reg  line_957_valid_reg;
  wire  line_958_clock;
  wire  line_958_reset;
  wire  line_958_valid;
  reg  line_958_valid_reg;
  wire  line_959_clock;
  wire  line_959_reset;
  wire  line_959_valid;
  reg  line_959_valid_reg;
  wire  line_960_clock;
  wire  line_960_reset;
  wire  line_960_valid;
  reg  line_960_valid_reg;
  wire  line_961_clock;
  wire  line_961_reset;
  wire  line_961_valid;
  reg  line_961_valid_reg;
  wire  line_962_clock;
  wire  line_962_reset;
  wire  line_962_valid;
  reg  line_962_valid_reg;
  wire  line_963_clock;
  wire  line_963_reset;
  wire  line_963_valid;
  reg  line_963_valid_reg;
  wire  line_964_clock;
  wire  line_964_reset;
  wire  line_964_valid;
  reg  line_964_valid_reg;
  wire  line_965_clock;
  wire  line_965_reset;
  wire  line_965_valid;
  reg  line_965_valid_reg;
  wire  line_966_clock;
  wire  line_966_reset;
  wire  line_966_valid;
  reg  line_966_valid_reg;
  wire  line_967_clock;
  wire  line_967_reset;
  wire  line_967_valid;
  reg  line_967_valid_reg;
  wire  line_968_clock;
  wire  line_968_reset;
  wire  line_968_valid;
  reg  line_968_valid_reg;
  wire  line_969_clock;
  wire  line_969_reset;
  wire  line_969_valid;
  reg  line_969_valid_reg;
  wire  line_970_clock;
  wire  line_970_reset;
  wire  line_970_valid;
  reg  line_970_valid_reg;
  wire  line_971_clock;
  wire  line_971_reset;
  wire  line_971_valid;
  reg  line_971_valid_reg;
  wire  line_972_clock;
  wire  line_972_reset;
  wire  line_972_valid;
  reg  line_972_valid_reg;
  wire  line_973_clock;
  wire  line_973_reset;
  wire  line_973_valid;
  reg  line_973_valid_reg;
  wire  line_974_clock;
  wire  line_974_reset;
  wire  line_974_valid;
  reg  line_974_valid_reg;
  wire  line_975_clock;
  wire  line_975_reset;
  wire  line_975_valid;
  reg  line_975_valid_reg;
  wire  line_976_clock;
  wire  line_976_reset;
  wire  line_976_valid;
  reg  line_976_valid_reg;
  wire  line_977_clock;
  wire  line_977_reset;
  wire  line_977_valid;
  reg  line_977_valid_reg;
  wire  line_978_clock;
  wire  line_978_reset;
  wire  line_978_valid;
  reg  line_978_valid_reg;
  wire  line_979_clock;
  wire  line_979_reset;
  wire  line_979_valid;
  reg  line_979_valid_reg;
  wire  line_980_clock;
  wire  line_980_reset;
  wire  line_980_valid;
  reg  line_980_valid_reg;
  wire  line_981_clock;
  wire  line_981_reset;
  wire  line_981_valid;
  reg  line_981_valid_reg;
  wire  line_982_clock;
  wire  line_982_reset;
  wire  line_982_valid;
  reg  line_982_valid_reg;
  wire  line_983_clock;
  wire  line_983_reset;
  wire  line_983_valid;
  reg  line_983_valid_reg;
  wire  line_984_clock;
  wire  line_984_reset;
  wire  line_984_valid;
  reg  line_984_valid_reg;
  wire  line_985_clock;
  wire  line_985_reset;
  wire  line_985_valid;
  reg  line_985_valid_reg;
  wire  line_986_clock;
  wire  line_986_reset;
  wire  line_986_valid;
  reg  line_986_valid_reg;
  wire  line_987_clock;
  wire  line_987_reset;
  wire  line_987_valid;
  reg  line_987_valid_reg;
  wire  line_988_clock;
  wire  line_988_reset;
  wire  line_988_valid;
  reg  line_988_valid_reg;
  wire  line_989_clock;
  wire  line_989_reset;
  wire  line_989_valid;
  reg  line_989_valid_reg;
  wire  line_990_clock;
  wire  line_990_reset;
  wire  line_990_valid;
  reg  line_990_valid_reg;
  wire  line_991_clock;
  wire  line_991_reset;
  wire  line_991_valid;
  reg  line_991_valid_reg;
  wire  line_992_clock;
  wire  line_992_reset;
  wire  line_992_valid;
  reg  line_992_valid_reg;
  wire  line_993_clock;
  wire  line_993_reset;
  wire  line_993_valid;
  reg  line_993_valid_reg;
  wire  line_994_clock;
  wire  line_994_reset;
  wire  line_994_valid;
  reg  line_994_valid_reg;
  wire  line_995_clock;
  wire  line_995_reset;
  wire  line_995_valid;
  reg  line_995_valid_reg;
  wire  line_996_clock;
  wire  line_996_reset;
  wire  line_996_valid;
  reg  line_996_valid_reg;
  wire  line_997_clock;
  wire  line_997_reset;
  wire  line_997_valid;
  reg  line_997_valid_reg;
  wire  line_998_clock;
  wire  line_998_reset;
  wire  line_998_valid;
  reg  line_998_valid_reg;
  wire  line_999_clock;
  wire  line_999_reset;
  wire  line_999_valid;
  reg  line_999_valid_reg;
  wire  line_1000_clock;
  wire  line_1000_reset;
  wire  line_1000_valid;
  reg  line_1000_valid_reg;
  wire  line_1001_clock;
  wire  line_1001_reset;
  wire  line_1001_valid;
  reg  line_1001_valid_reg;
  wire  line_1002_clock;
  wire  line_1002_reset;
  wire  line_1002_valid;
  reg  line_1002_valid_reg;
  wire  line_1003_clock;
  wire  line_1003_reset;
  wire  line_1003_valid;
  reg  line_1003_valid_reg;
  wire  line_1004_clock;
  wire  line_1004_reset;
  wire  line_1004_valid;
  reg  line_1004_valid_reg;
  wire  line_1005_clock;
  wire  line_1005_reset;
  wire  line_1005_valid;
  reg  line_1005_valid_reg;
  wire  line_1006_clock;
  wire  line_1006_reset;
  wire  line_1006_valid;
  reg  line_1006_valid_reg;
  wire  line_1007_clock;
  wire  line_1007_reset;
  wire  line_1007_valid;
  reg  line_1007_valid_reg;
  wire  line_1008_clock;
  wire  line_1008_reset;
  wire  line_1008_valid;
  reg  line_1008_valid_reg;
  wire  line_1009_clock;
  wire  line_1009_reset;
  wire  line_1009_valid;
  reg  line_1009_valid_reg;
  wire  line_1010_clock;
  wire  line_1010_reset;
  wire  line_1010_valid;
  reg  line_1010_valid_reg;
  wire  line_1011_clock;
  wire  line_1011_reset;
  wire  line_1011_valid;
  reg  line_1011_valid_reg;
  wire  line_1012_clock;
  wire  line_1012_reset;
  wire  line_1012_valid;
  reg  line_1012_valid_reg;
  wire  line_1013_clock;
  wire  line_1013_reset;
  wire  line_1013_valid;
  reg  line_1013_valid_reg;
  wire  line_1014_clock;
  wire  line_1014_reset;
  wire  line_1014_valid;
  reg  line_1014_valid_reg;
  wire  line_1015_clock;
  wire  line_1015_reset;
  wire  line_1015_valid;
  reg  line_1015_valid_reg;
  wire  line_1016_clock;
  wire  line_1016_reset;
  wire  line_1016_valid;
  reg  line_1016_valid_reg;
  wire  line_1017_clock;
  wire  line_1017_reset;
  wire  line_1017_valid;
  reg  line_1017_valid_reg;
  wire  line_1018_clock;
  wire  line_1018_reset;
  wire  line_1018_valid;
  reg  line_1018_valid_reg;
  wire  line_1019_clock;
  wire  line_1019_reset;
  wire  line_1019_valid;
  reg  line_1019_valid_reg;
  wire  line_1020_clock;
  wire  line_1020_reset;
  wire  line_1020_valid;
  reg  line_1020_valid_reg;
  wire  line_1021_clock;
  wire  line_1021_reset;
  wire  line_1021_valid;
  reg  line_1021_valid_reg;
  wire  line_1022_clock;
  wire  line_1022_reset;
  wire  line_1022_valid;
  reg  line_1022_valid_reg;
  wire  line_1023_clock;
  wire  line_1023_reset;
  wire  line_1023_valid;
  reg  line_1023_valid_reg;
  wire  line_1024_clock;
  wire  line_1024_reset;
  wire  line_1024_valid;
  reg  line_1024_valid_reg;
  wire  line_1025_clock;
  wire  line_1025_reset;
  wire  line_1025_valid;
  reg  line_1025_valid_reg;
  wire  line_1026_clock;
  wire  line_1026_reset;
  wire  line_1026_valid;
  reg  line_1026_valid_reg;
  wire  line_1027_clock;
  wire  line_1027_reset;
  wire  line_1027_valid;
  reg  line_1027_valid_reg;
  wire  line_1028_clock;
  wire  line_1028_reset;
  wire  line_1028_valid;
  reg  line_1028_valid_reg;
  wire  line_1029_clock;
  wire  line_1029_reset;
  wire  line_1029_valid;
  reg  line_1029_valid_reg;
  wire  line_1030_clock;
  wire  line_1030_reset;
  wire  line_1030_valid;
  reg  line_1030_valid_reg;
  wire  line_1031_clock;
  wire  line_1031_reset;
  wire  line_1031_valid;
  reg  line_1031_valid_reg;
  wire  line_1032_clock;
  wire  line_1032_reset;
  wire  line_1032_valid;
  reg  line_1032_valid_reg;
  wire  line_1033_clock;
  wire  line_1033_reset;
  wire  line_1033_valid;
  reg  line_1033_valid_reg;
  wire  line_1034_clock;
  wire  line_1034_reset;
  wire  line_1034_valid;
  reg  line_1034_valid_reg;
  wire  line_1035_clock;
  wire  line_1035_reset;
  wire  line_1035_valid;
  reg  line_1035_valid_reg;
  wire  line_1036_clock;
  wire  line_1036_reset;
  wire  line_1036_valid;
  reg  line_1036_valid_reg;
  wire  line_1037_clock;
  wire  line_1037_reset;
  wire  line_1037_valid;
  reg  line_1037_valid_reg;
  wire  line_1038_clock;
  wire  line_1038_reset;
  wire  line_1038_valid;
  reg  line_1038_valid_reg;
  wire  line_1039_clock;
  wire  line_1039_reset;
  wire  line_1039_valid;
  reg  line_1039_valid_reg;
  wire  line_1040_clock;
  wire  line_1040_reset;
  wire  line_1040_valid;
  reg  line_1040_valid_reg;
  wire  line_1041_clock;
  wire  line_1041_reset;
  wire  line_1041_valid;
  reg  line_1041_valid_reg;
  wire  line_1042_clock;
  wire  line_1042_reset;
  wire  line_1042_valid;
  reg  line_1042_valid_reg;
  wire  line_1043_clock;
  wire  line_1043_reset;
  wire  line_1043_valid;
  reg  line_1043_valid_reg;
  wire  line_1044_clock;
  wire  line_1044_reset;
  wire  line_1044_valid;
  reg  line_1044_valid_reg;
  wire  line_1045_clock;
  wire  line_1045_reset;
  wire  line_1045_valid;
  reg  line_1045_valid_reg;
  wire  line_1046_clock;
  wire  line_1046_reset;
  wire  line_1046_valid;
  reg  line_1046_valid_reg;
  wire  line_1047_clock;
  wire  line_1047_reset;
  wire  line_1047_valid;
  reg  line_1047_valid_reg;
  wire  line_1048_clock;
  wire  line_1048_reset;
  wire  line_1048_valid;
  reg  line_1048_valid_reg;
  wire  line_1049_clock;
  wire  line_1049_reset;
  wire  line_1049_valid;
  reg  line_1049_valid_reg;
  wire  line_1050_clock;
  wire  line_1050_reset;
  wire  line_1050_valid;
  reg  line_1050_valid_reg;
  wire  line_1051_clock;
  wire  line_1051_reset;
  wire  line_1051_valid;
  reg  line_1051_valid_reg;
  wire  line_1052_clock;
  wire  line_1052_reset;
  wire  line_1052_valid;
  reg  line_1052_valid_reg;
  wire  line_1053_clock;
  wire  line_1053_reset;
  wire  line_1053_valid;
  reg  line_1053_valid_reg;
  wire  line_1054_clock;
  wire  line_1054_reset;
  wire  line_1054_valid;
  reg  line_1054_valid_reg;
  wire  line_1055_clock;
  wire  line_1055_reset;
  wire  line_1055_valid;
  reg  line_1055_valid_reg;
  wire  line_1056_clock;
  wire  line_1056_reset;
  wire  line_1056_valid;
  reg  line_1056_valid_reg;
  wire  line_1057_clock;
  wire  line_1057_reset;
  wire  line_1057_valid;
  reg  line_1057_valid_reg;
  wire  line_1058_clock;
  wire  line_1058_reset;
  wire  line_1058_valid;
  reg  line_1058_valid_reg;
  wire  line_1059_clock;
  wire  line_1059_reset;
  wire  line_1059_valid;
  reg  line_1059_valid_reg;
  wire  line_1060_clock;
  wire  line_1060_reset;
  wire  line_1060_valid;
  reg  line_1060_valid_reg;
  wire  line_1061_clock;
  wire  line_1061_reset;
  wire  line_1061_valid;
  reg  line_1061_valid_reg;
  wire  line_1062_clock;
  wire  line_1062_reset;
  wire  line_1062_valid;
  reg  line_1062_valid_reg;
  wire  line_1063_clock;
  wire  line_1063_reset;
  wire  line_1063_valid;
  reg  line_1063_valid_reg;
  wire  line_1064_clock;
  wire  line_1064_reset;
  wire  line_1064_valid;
  reg  line_1064_valid_reg;
  wire  line_1065_clock;
  wire  line_1065_reset;
  wire  line_1065_valid;
  reg  line_1065_valid_reg;
  wire  line_1066_clock;
  wire  line_1066_reset;
  wire  line_1066_valid;
  reg  line_1066_valid_reg;
  wire  line_1067_clock;
  wire  line_1067_reset;
  wire  line_1067_valid;
  reg  line_1067_valid_reg;
  wire  line_1068_clock;
  wire  line_1068_reset;
  wire  line_1068_valid;
  reg  line_1068_valid_reg;
  wire  line_1069_clock;
  wire  line_1069_reset;
  wire  line_1069_valid;
  reg  line_1069_valid_reg;
  wire  line_1070_clock;
  wire  line_1070_reset;
  wire  line_1070_valid;
  reg  line_1070_valid_reg;
  wire  line_1071_clock;
  wire  line_1071_reset;
  wire  line_1071_valid;
  reg  line_1071_valid_reg;
  wire  line_1072_clock;
  wire  line_1072_reset;
  wire  line_1072_valid;
  reg  line_1072_valid_reg;
  wire  line_1073_clock;
  wire  line_1073_reset;
  wire  line_1073_valid;
  reg  line_1073_valid_reg;
  wire  line_1074_clock;
  wire  line_1074_reset;
  wire  line_1074_valid;
  reg  line_1074_valid_reg;
  wire  line_1075_clock;
  wire  line_1075_reset;
  wire  line_1075_valid;
  reg  line_1075_valid_reg;
  wire  line_1076_clock;
  wire  line_1076_reset;
  wire  line_1076_valid;
  reg  line_1076_valid_reg;
  wire  line_1077_clock;
  wire  line_1077_reset;
  wire  line_1077_valid;
  reg  line_1077_valid_reg;
  wire  line_1078_clock;
  wire  line_1078_reset;
  wire  line_1078_valid;
  reg  line_1078_valid_reg;
  wire  line_1079_clock;
  wire  line_1079_reset;
  wire  line_1079_valid;
  reg  line_1079_valid_reg;
  wire  line_1080_clock;
  wire  line_1080_reset;
  wire  line_1080_valid;
  reg  line_1080_valid_reg;
  wire  line_1081_clock;
  wire  line_1081_reset;
  wire  line_1081_valid;
  reg  line_1081_valid_reg;
  wire  line_1082_clock;
  wire  line_1082_reset;
  wire  line_1082_valid;
  reg  line_1082_valid_reg;
  wire  line_1083_clock;
  wire  line_1083_reset;
  wire  line_1083_valid;
  reg  line_1083_valid_reg;
  wire  line_1084_clock;
  wire  line_1084_reset;
  wire  line_1084_valid;
  reg  line_1084_valid_reg;
  wire  line_1085_clock;
  wire  line_1085_reset;
  wire  line_1085_valid;
  reg  line_1085_valid_reg;
  wire  line_1086_clock;
  wire  line_1086_reset;
  wire  line_1086_valid;
  reg  line_1086_valid_reg;
  wire  line_1087_clock;
  wire  line_1087_reset;
  wire  line_1087_valid;
  reg  line_1087_valid_reg;
  wire  line_1088_clock;
  wire  line_1088_reset;
  wire  line_1088_valid;
  reg  line_1088_valid_reg;
  wire  line_1089_clock;
  wire  line_1089_reset;
  wire  line_1089_valid;
  reg  line_1089_valid_reg;
  wire  line_1090_clock;
  wire  line_1090_reset;
  wire  line_1090_valid;
  reg  line_1090_valid_reg;
  wire  line_1091_clock;
  wire  line_1091_reset;
  wire  line_1091_valid;
  reg  line_1091_valid_reg;
  wire  line_1092_clock;
  wire  line_1092_reset;
  wire  line_1092_valid;
  reg  line_1092_valid_reg;
  wire  line_1093_clock;
  wire  line_1093_reset;
  wire  line_1093_valid;
  reg  line_1093_valid_reg;
  wire  line_1094_clock;
  wire  line_1094_reset;
  wire  line_1094_valid;
  reg  line_1094_valid_reg;
  wire  line_1095_clock;
  wire  line_1095_reset;
  wire  line_1095_valid;
  reg  line_1095_valid_reg;
  wire  line_1096_clock;
  wire  line_1096_reset;
  wire  line_1096_valid;
  reg  line_1096_valid_reg;
  wire  line_1097_clock;
  wire  line_1097_reset;
  wire  line_1097_valid;
  reg  line_1097_valid_reg;
  wire  line_1098_clock;
  wire  line_1098_reset;
  wire  line_1098_valid;
  reg  line_1098_valid_reg;
  wire  line_1099_clock;
  wire  line_1099_reset;
  wire  line_1099_valid;
  reg  line_1099_valid_reg;
  wire  line_1100_clock;
  wire  line_1100_reset;
  wire  line_1100_valid;
  reg  line_1100_valid_reg;
  wire  line_1101_clock;
  wire  line_1101_reset;
  wire  line_1101_valid;
  reg  line_1101_valid_reg;
  wire  line_1102_clock;
  wire  line_1102_reset;
  wire  line_1102_valid;
  reg  line_1102_valid_reg;
  wire  line_1103_clock;
  wire  line_1103_reset;
  wire  line_1103_valid;
  reg  line_1103_valid_reg;
  wire  line_1104_clock;
  wire  line_1104_reset;
  wire  line_1104_valid;
  reg  line_1104_valid_reg;
  wire  line_1105_clock;
  wire  line_1105_reset;
  wire  line_1105_valid;
  reg  line_1105_valid_reg;
  wire  line_1106_clock;
  wire  line_1106_reset;
  wire  line_1106_valid;
  reg  line_1106_valid_reg;
  wire  line_1107_clock;
  wire  line_1107_reset;
  wire  line_1107_valid;
  reg  line_1107_valid_reg;
  wire  line_1108_clock;
  wire  line_1108_reset;
  wire  line_1108_valid;
  reg  line_1108_valid_reg;
  wire  line_1109_clock;
  wire  line_1109_reset;
  wire  line_1109_valid;
  reg  line_1109_valid_reg;
  wire  line_1110_clock;
  wire  line_1110_reset;
  wire  line_1110_valid;
  reg  line_1110_valid_reg;
  wire  line_1111_clock;
  wire  line_1111_reset;
  wire  line_1111_valid;
  reg  line_1111_valid_reg;
  wire  line_1112_clock;
  wire  line_1112_reset;
  wire  line_1112_valid;
  reg  line_1112_valid_reg;
  wire  line_1113_clock;
  wire  line_1113_reset;
  wire  line_1113_valid;
  reg  line_1113_valid_reg;
  wire  line_1114_clock;
  wire  line_1114_reset;
  wire  line_1114_valid;
  reg  line_1114_valid_reg;
  wire  line_1115_clock;
  wire  line_1115_reset;
  wire  line_1115_valid;
  reg  line_1115_valid_reg;
  wire  line_1116_clock;
  wire  line_1116_reset;
  wire  line_1116_valid;
  reg  line_1116_valid_reg;
  wire  line_1117_clock;
  wire  line_1117_reset;
  wire  line_1117_valid;
  reg  line_1117_valid_reg;
  wire  line_1118_clock;
  wire  line_1118_reset;
  wire  line_1118_valid;
  reg  line_1118_valid_reg;
  wire  line_1119_clock;
  wire  line_1119_reset;
  wire  line_1119_valid;
  reg  line_1119_valid_reg;
  wire  line_1120_clock;
  wire  line_1120_reset;
  wire  line_1120_valid;
  reg  line_1120_valid_reg;
  wire  line_1121_clock;
  wire  line_1121_reset;
  wire  line_1121_valid;
  reg  line_1121_valid_reg;
  wire  line_1122_clock;
  wire  line_1122_reset;
  wire  line_1122_valid;
  reg  line_1122_valid_reg;
  wire  line_1123_clock;
  wire  line_1123_reset;
  wire  line_1123_valid;
  reg  line_1123_valid_reg;
  wire  line_1124_clock;
  wire  line_1124_reset;
  wire  line_1124_valid;
  reg  line_1124_valid_reg;
  wire  line_1125_clock;
  wire  line_1125_reset;
  wire  line_1125_valid;
  reg  line_1125_valid_reg;
  wire  line_1126_clock;
  wire  line_1126_reset;
  wire  line_1126_valid;
  reg  line_1126_valid_reg;
  wire  line_1127_clock;
  wire  line_1127_reset;
  wire  line_1127_valid;
  reg  line_1127_valid_reg;
  wire  line_1128_clock;
  wire  line_1128_reset;
  wire  line_1128_valid;
  reg  line_1128_valid_reg;
  wire  line_1129_clock;
  wire  line_1129_reset;
  wire  line_1129_valid;
  reg  line_1129_valid_reg;
  wire  line_1130_clock;
  wire  line_1130_reset;
  wire  line_1130_valid;
  reg  line_1130_valid_reg;
  wire  line_1131_clock;
  wire  line_1131_reset;
  wire  line_1131_valid;
  reg  line_1131_valid_reg;
  wire  line_1132_clock;
  wire  line_1132_reset;
  wire  line_1132_valid;
  reg  line_1132_valid_reg;
  wire  line_1133_clock;
  wire  line_1133_reset;
  wire  line_1133_valid;
  reg  line_1133_valid_reg;
  wire  line_1134_clock;
  wire  line_1134_reset;
  wire  line_1134_valid;
  reg  line_1134_valid_reg;
  wire  line_1135_clock;
  wire  line_1135_reset;
  wire  line_1135_valid;
  reg  line_1135_valid_reg;
  wire  line_1136_clock;
  wire  line_1136_reset;
  wire  line_1136_valid;
  reg  line_1136_valid_reg;
  wire  line_1137_clock;
  wire  line_1137_reset;
  wire  line_1137_valid;
  reg  line_1137_valid_reg;
  wire  line_1138_clock;
  wire  line_1138_reset;
  wire  line_1138_valid;
  reg  line_1138_valid_reg;
  wire  line_1139_clock;
  wire  line_1139_reset;
  wire  line_1139_valid;
  reg  line_1139_valid_reg;
  wire  line_1140_clock;
  wire  line_1140_reset;
  wire  line_1140_valid;
  reg  line_1140_valid_reg;
  wire  line_1141_clock;
  wire  line_1141_reset;
  wire  line_1141_valid;
  reg  line_1141_valid_reg;
  wire  line_1142_clock;
  wire  line_1142_reset;
  wire  line_1142_valid;
  reg  line_1142_valid_reg;
  wire  line_1143_clock;
  wire  line_1143_reset;
  wire  line_1143_valid;
  reg  line_1143_valid_reg;
  wire  line_1144_clock;
  wire  line_1144_reset;
  wire  line_1144_valid;
  reg  line_1144_valid_reg;
  wire  line_1145_clock;
  wire  line_1145_reset;
  wire  line_1145_valid;
  reg  line_1145_valid_reg;
  wire  line_1146_clock;
  wire  line_1146_reset;
  wire  line_1146_valid;
  reg  line_1146_valid_reg;
  wire  line_1147_clock;
  wire  line_1147_reset;
  wire  line_1147_valid;
  reg  line_1147_valid_reg;
  wire  line_1148_clock;
  wire  line_1148_reset;
  wire  line_1148_valid;
  reg  line_1148_valid_reg;
  wire  line_1149_clock;
  wire  line_1149_reset;
  wire  line_1149_valid;
  reg  line_1149_valid_reg;
  wire  line_1150_clock;
  wire  line_1150_reset;
  wire  line_1150_valid;
  reg  line_1150_valid_reg;
  wire  line_1151_clock;
  wire  line_1151_reset;
  wire  line_1151_valid;
  reg  line_1151_valid_reg;
  wire  line_1152_clock;
  wire  line_1152_reset;
  wire  line_1152_valid;
  reg  line_1152_valid_reg;
  wire  line_1153_clock;
  wire  line_1153_reset;
  wire  line_1153_valid;
  reg  line_1153_valid_reg;
  wire  line_1154_clock;
  wire  line_1154_reset;
  wire  line_1154_valid;
  reg  line_1154_valid_reg;
  wire  line_1155_clock;
  wire  line_1155_reset;
  wire  line_1155_valid;
  reg  line_1155_valid_reg;
  wire  line_1156_clock;
  wire  line_1156_reset;
  wire  line_1156_valid;
  reg  line_1156_valid_reg;
  wire  line_1157_clock;
  wire  line_1157_reset;
  wire  line_1157_valid;
  reg  line_1157_valid_reg;
  wire  line_1158_clock;
  wire  line_1158_reset;
  wire  line_1158_valid;
  reg  line_1158_valid_reg;
  wire  line_1159_clock;
  wire  line_1159_reset;
  wire  line_1159_valid;
  reg  line_1159_valid_reg;
  wire  line_1160_clock;
  wire  line_1160_reset;
  wire  line_1160_valid;
  reg  line_1160_valid_reg;
  wire  line_1161_clock;
  wire  line_1161_reset;
  wire  line_1161_valid;
  reg  line_1161_valid_reg;
  wire  line_1162_clock;
  wire  line_1162_reset;
  wire  line_1162_valid;
  reg  line_1162_valid_reg;
  wire  line_1163_clock;
  wire  line_1163_reset;
  wire  line_1163_valid;
  reg  line_1163_valid_reg;
  wire  line_1164_clock;
  wire  line_1164_reset;
  wire  line_1164_valid;
  reg  line_1164_valid_reg;
  wire  line_1165_clock;
  wire  line_1165_reset;
  wire  line_1165_valid;
  reg  line_1165_valid_reg;
  wire  line_1166_clock;
  wire  line_1166_reset;
  wire  line_1166_valid;
  reg  line_1166_valid_reg;
  wire  line_1167_clock;
  wire  line_1167_reset;
  wire  line_1167_valid;
  reg  line_1167_valid_reg;
  wire  line_1168_clock;
  wire  line_1168_reset;
  wire  line_1168_valid;
  reg  line_1168_valid_reg;
  wire  line_1169_clock;
  wire  line_1169_reset;
  wire  line_1169_valid;
  reg  line_1169_valid_reg;
  wire  line_1170_clock;
  wire  line_1170_reset;
  wire  line_1170_valid;
  reg  line_1170_valid_reg;
  wire  line_1171_clock;
  wire  line_1171_reset;
  wire  line_1171_valid;
  reg  line_1171_valid_reg;
  wire  line_1172_clock;
  wire  line_1172_reset;
  wire  line_1172_valid;
  reg  line_1172_valid_reg;
  wire  line_1173_clock;
  wire  line_1173_reset;
  wire  line_1173_valid;
  reg  line_1173_valid_reg;
  wire  line_1174_clock;
  wire  line_1174_reset;
  wire  line_1174_valid;
  reg  line_1174_valid_reg;
  wire  line_1175_clock;
  wire  line_1175_reset;
  wire  line_1175_valid;
  reg  line_1175_valid_reg;
  wire  line_1176_clock;
  wire  line_1176_reset;
  wire  line_1176_valid;
  reg  line_1176_valid_reg;
  wire  line_1177_clock;
  wire  line_1177_reset;
  wire  line_1177_valid;
  reg  line_1177_valid_reg;
  wire [1:0] _ringBufferHead_T_1 = ringBufferHead + enqueueSize; // @[src/main/scala/utils/PipelineVector.scala 47:42]
  wire  line_1178_clock;
  wire  line_1178_reset;
  wire  line_1178_valid;
  reg  line_1178_valid_reg;
  wire  line_1179_clock;
  wire  line_1179_reset;
  wire  line_1179_valid;
  reg  line_1179_valid_reg;
  wire [63:0] _GEN_2023 = 2'h1 == ringBufferTail ? dataBuffer_1_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1180_clock;
  wire  line_1180_reset;
  wire  line_1180_valid;
  reg  line_1180_valid_reg;
  wire [63:0] _GEN_2024 = 2'h2 == ringBufferTail ? dataBuffer_2_data_imm : _GEN_2023; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1181_clock;
  wire  line_1181_reset;
  wire  line_1181_valid;
  reg  line_1181_valid_reg;
  wire  line_1182_clock;
  wire  line_1182_reset;
  wire  line_1182_valid;
  reg  line_1182_valid_reg;
  wire  line_1183_clock;
  wire  line_1183_reset;
  wire  line_1183_valid;
  reg  line_1183_valid_reg;
  wire  line_1184_clock;
  wire  line_1184_reset;
  wire  line_1184_valid;
  reg  line_1184_valid_reg;
  wire  line_1185_clock;
  wire  line_1185_reset;
  wire  line_1185_valid;
  reg  line_1185_valid_reg;
  wire  line_1186_clock;
  wire  line_1186_reset;
  wire  line_1186_valid;
  reg  line_1186_valid_reg;
  wire  line_1187_clock;
  wire  line_1187_reset;
  wire  line_1187_valid;
  reg  line_1187_valid_reg;
  wire  line_1188_clock;
  wire  line_1188_reset;
  wire  line_1188_valid;
  reg  line_1188_valid_reg;
  wire  line_1189_clock;
  wire  line_1189_reset;
  wire  line_1189_valid;
  reg  line_1189_valid_reg;
  wire  line_1190_clock;
  wire  line_1190_reset;
  wire  line_1190_valid;
  reg  line_1190_valid_reg;
  wire  line_1191_clock;
  wire  line_1191_reset;
  wire  line_1191_valid;
  reg  line_1191_valid_reg;
  wire  line_1192_clock;
  wire  line_1192_reset;
  wire  line_1192_valid;
  reg  line_1192_valid_reg;
  wire  line_1193_clock;
  wire  line_1193_reset;
  wire  line_1193_valid;
  reg  line_1193_valid_reg;
  wire  line_1194_clock;
  wire  line_1194_reset;
  wire  line_1194_valid;
  reg  line_1194_valid_reg;
  wire  line_1195_clock;
  wire  line_1195_reset;
  wire  line_1195_valid;
  reg  line_1195_valid_reg;
  wire  line_1196_clock;
  wire  line_1196_reset;
  wire  line_1196_valid;
  reg  line_1196_valid_reg;
  wire  line_1197_clock;
  wire  line_1197_reset;
  wire  line_1197_valid;
  reg  line_1197_valid_reg;
  wire  line_1198_clock;
  wire  line_1198_reset;
  wire  line_1198_valid;
  reg  line_1198_valid_reg;
  wire  line_1199_clock;
  wire  line_1199_reset;
  wire  line_1199_valid;
  reg  line_1199_valid_reg;
  wire  line_1200_clock;
  wire  line_1200_reset;
  wire  line_1200_valid;
  reg  line_1200_valid_reg;
  wire  line_1201_clock;
  wire  line_1201_reset;
  wire  line_1201_valid;
  reg  line_1201_valid_reg;
  wire  line_1202_clock;
  wire  line_1202_reset;
  wire  line_1202_valid;
  reg  line_1202_valid_reg;
  wire  line_1203_clock;
  wire  line_1203_reset;
  wire  line_1203_valid;
  reg  line_1203_valid_reg;
  wire  line_1204_clock;
  wire  line_1204_reset;
  wire  line_1204_valid;
  reg  line_1204_valid_reg;
  wire  line_1205_clock;
  wire  line_1205_reset;
  wire  line_1205_valid;
  reg  line_1205_valid_reg;
  wire  line_1206_clock;
  wire  line_1206_reset;
  wire  line_1206_valid;
  reg  line_1206_valid_reg;
  wire  line_1207_clock;
  wire  line_1207_reset;
  wire  line_1207_valid;
  reg  line_1207_valid_reg;
  wire  _GEN_2051 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_isNutCoreTrap : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1208_clock;
  wire  line_1208_reset;
  wire  line_1208_valid;
  reg  line_1208_valid_reg;
  wire  _GEN_2052 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_isNutCoreTrap : _GEN_2051; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1209_clock;
  wire  line_1209_reset;
  wire  line_1209_valid;
  reg  line_1209_valid_reg;
  wire  line_1210_clock;
  wire  line_1210_reset;
  wire  line_1210_valid;
  reg  line_1210_valid_reg;
  wire  line_1211_clock;
  wire  line_1211_reset;
  wire  line_1211_valid;
  reg  line_1211_valid_reg;
  wire [4:0] _GEN_2055 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1212_clock;
  wire  line_1212_reset;
  wire  line_1212_valid;
  reg  line_1212_valid_reg;
  wire [4:0] _GEN_2056 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfDest : _GEN_2055; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1213_clock;
  wire  line_1213_reset;
  wire  line_1213_valid;
  reg  line_1213_valid_reg;
  wire  line_1214_clock;
  wire  line_1214_reset;
  wire  line_1214_valid;
  reg  line_1214_valid_reg;
  wire  line_1215_clock;
  wire  line_1215_reset;
  wire  line_1215_valid;
  reg  line_1215_valid_reg;
  wire  _GEN_2059 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1216_clock;
  wire  line_1216_reset;
  wire  line_1216_valid;
  reg  line_1216_valid_reg;
  wire  _GEN_2060 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfWen : _GEN_2059; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1217_clock;
  wire  line_1217_reset;
  wire  line_1217_valid;
  reg  line_1217_valid_reg;
  wire  line_1218_clock;
  wire  line_1218_reset;
  wire  line_1218_valid;
  reg  line_1218_valid_reg;
  wire  line_1219_clock;
  wire  line_1219_reset;
  wire  line_1219_valid;
  reg  line_1219_valid_reg;
  wire [4:0] _GEN_2063 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1220_clock;
  wire  line_1220_reset;
  wire  line_1220_valid;
  reg  line_1220_valid_reg;
  wire [4:0] _GEN_2064 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc2 : _GEN_2063; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1221_clock;
  wire  line_1221_reset;
  wire  line_1221_valid;
  reg  line_1221_valid_reg;
  wire  line_1222_clock;
  wire  line_1222_reset;
  wire  line_1222_valid;
  reg  line_1222_valid_reg;
  wire  line_1223_clock;
  wire  line_1223_reset;
  wire  line_1223_valid;
  reg  line_1223_valid_reg;
  wire [4:0] _GEN_2067 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1224_clock;
  wire  line_1224_reset;
  wire  line_1224_valid;
  reg  line_1224_valid_reg;
  wire [4:0] _GEN_2068 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc1 : _GEN_2067; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1225_clock;
  wire  line_1225_reset;
  wire  line_1225_valid;
  reg  line_1225_valid_reg;
  wire  line_1226_clock;
  wire  line_1226_reset;
  wire  line_1226_valid;
  reg  line_1226_valid_reg;
  wire  line_1227_clock;
  wire  line_1227_reset;
  wire  line_1227_valid;
  reg  line_1227_valid_reg;
  wire [6:0] _GEN_2071 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1228_clock;
  wire  line_1228_reset;
  wire  line_1228_valid;
  reg  line_1228_valid_reg;
  wire [6:0] _GEN_2072 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuOpType : _GEN_2071; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1229_clock;
  wire  line_1229_reset;
  wire  line_1229_valid;
  reg  line_1229_valid_reg;
  wire  line_1230_clock;
  wire  line_1230_reset;
  wire  line_1230_valid;
  reg  line_1230_valid_reg;
  wire  line_1231_clock;
  wire  line_1231_reset;
  wire  line_1231_valid;
  reg  line_1231_valid_reg;
  wire [2:0] _GEN_2075 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1232_clock;
  wire  line_1232_reset;
  wire  line_1232_valid;
  reg  line_1232_valid_reg;
  wire [2:0] _GEN_2076 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuType : _GEN_2075; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1233_clock;
  wire  line_1233_reset;
  wire  line_1233_valid;
  reg  line_1233_valid_reg;
  wire  line_1234_clock;
  wire  line_1234_reset;
  wire  line_1234_valid;
  reg  line_1234_valid_reg;
  wire  line_1235_clock;
  wire  line_1235_reset;
  wire  line_1235_valid;
  reg  line_1235_valid_reg;
  wire  _GEN_2079 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1236_clock;
  wire  line_1236_reset;
  wire  line_1236_valid;
  reg  line_1236_valid_reg;
  wire  _GEN_2080 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src2Type : _GEN_2079; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1237_clock;
  wire  line_1237_reset;
  wire  line_1237_valid;
  reg  line_1237_valid_reg;
  wire  line_1238_clock;
  wire  line_1238_reset;
  wire  line_1238_valid;
  reg  line_1238_valid_reg;
  wire  line_1239_clock;
  wire  line_1239_reset;
  wire  line_1239_valid;
  reg  line_1239_valid_reg;
  wire  _GEN_2083 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1240_clock;
  wire  line_1240_reset;
  wire  line_1240_valid;
  reg  line_1240_valid_reg;
  wire  _GEN_2084 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src1Type : _GEN_2083; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1241_clock;
  wire  line_1241_reset;
  wire  line_1241_valid;
  reg  line_1241_valid_reg;
  wire  line_1242_clock;
  wire  line_1242_reset;
  wire  line_1242_valid;
  reg  line_1242_valid_reg;
  wire  line_1243_clock;
  wire  line_1243_reset;
  wire  line_1243_valid;
  reg  line_1243_valid_reg;
  wire  line_1244_clock;
  wire  line_1244_reset;
  wire  line_1244_valid;
  reg  line_1244_valid_reg;
  wire  line_1245_clock;
  wire  line_1245_reset;
  wire  line_1245_valid;
  reg  line_1245_valid_reg;
  wire  line_1246_clock;
  wire  line_1246_reset;
  wire  line_1246_valid;
  reg  line_1246_valid_reg;
  wire  line_1247_clock;
  wire  line_1247_reset;
  wire  line_1247_valid;
  reg  line_1247_valid_reg;
  wire  line_1248_clock;
  wire  line_1248_reset;
  wire  line_1248_valid;
  reg  line_1248_valid_reg;
  wire  line_1249_clock;
  wire  line_1249_reset;
  wire  line_1249_valid;
  reg  line_1249_valid_reg;
  wire  line_1250_clock;
  wire  line_1250_reset;
  wire  line_1250_valid;
  reg  line_1250_valid_reg;
  wire  line_1251_clock;
  wire  line_1251_reset;
  wire  line_1251_valid;
  reg  line_1251_valid_reg;
  wire  line_1252_clock;
  wire  line_1252_reset;
  wire  line_1252_valid;
  reg  line_1252_valid_reg;
  wire  line_1253_clock;
  wire  line_1253_reset;
  wire  line_1253_valid;
  reg  line_1253_valid_reg;
  wire  line_1254_clock;
  wire  line_1254_reset;
  wire  line_1254_valid;
  reg  line_1254_valid_reg;
  wire  line_1255_clock;
  wire  line_1255_reset;
  wire  line_1255_valid;
  reg  line_1255_valid_reg;
  wire  _GEN_2099 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_crossBoundaryFault : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1256_clock;
  wire  line_1256_reset;
  wire  line_1256_valid;
  reg  line_1256_valid_reg;
  wire  _GEN_2100 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_crossBoundaryFault : _GEN_2099; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1257_clock;
  wire  line_1257_reset;
  wire  line_1257_valid;
  reg  line_1257_valid_reg;
  wire  line_1258_clock;
  wire  line_1258_reset;
  wire  line_1258_valid;
  reg  line_1258_valid_reg;
  wire  line_1259_clock;
  wire  line_1259_reset;
  wire  line_1259_valid;
  reg  line_1259_valid_reg;
  wire  line_1260_clock;
  wire  line_1260_reset;
  wire  line_1260_valid;
  reg  line_1260_valid_reg;
  wire  line_1261_clock;
  wire  line_1261_reset;
  wire  line_1261_valid;
  reg  line_1261_valid_reg;
  wire  line_1262_clock;
  wire  line_1262_reset;
  wire  line_1262_valid;
  reg  line_1262_valid_reg;
  wire  line_1263_clock;
  wire  line_1263_reset;
  wire  line_1263_valid;
  reg  line_1263_valid_reg;
  wire [3:0] _GEN_2107 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1264_clock;
  wire  line_1264_reset;
  wire  line_1264_valid;
  reg  line_1264_valid_reg;
  wire [3:0] _GEN_2108 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_brIdx : _GEN_2107; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1265_clock;
  wire  line_1265_reset;
  wire  line_1265_valid;
  reg  line_1265_valid_reg;
  wire  line_1266_clock;
  wire  line_1266_reset;
  wire  line_1266_valid;
  reg  line_1266_valid_reg;
  wire  line_1267_clock;
  wire  line_1267_reset;
  wire  line_1267_valid;
  reg  line_1267_valid_reg;
  wire  line_1268_clock;
  wire  line_1268_reset;
  wire  line_1268_valid;
  reg  line_1268_valid_reg;
  wire  line_1269_clock;
  wire  line_1269_reset;
  wire  line_1269_valid;
  reg  line_1269_valid_reg;
  wire  line_1270_clock;
  wire  line_1270_reset;
  wire  line_1270_valid;
  reg  line_1270_valid_reg;
  wire  line_1271_clock;
  wire  line_1271_reset;
  wire  line_1271_valid;
  reg  line_1271_valid_reg;
  wire  _GEN_2115 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1272_clock;
  wire  line_1272_reset;
  wire  line_1272_valid;
  reg  line_1272_valid_reg;
  wire  _GEN_2116 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_1 : _GEN_2115; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1273_clock;
  wire  line_1273_reset;
  wire  line_1273_valid;
  reg  line_1273_valid_reg;
  wire  line_1274_clock;
  wire  line_1274_reset;
  wire  line_1274_valid;
  reg  line_1274_valid_reg;
  wire  line_1275_clock;
  wire  line_1275_reset;
  wire  line_1275_valid;
  reg  line_1275_valid_reg;
  wire  line_1276_clock;
  wire  line_1276_reset;
  wire  line_1276_valid;
  reg  line_1276_valid_reg;
  wire  line_1277_clock;
  wire  line_1277_reset;
  wire  line_1277_valid;
  reg  line_1277_valid_reg;
  wire  line_1278_clock;
  wire  line_1278_reset;
  wire  line_1278_valid;
  reg  line_1278_valid_reg;
  wire  line_1279_clock;
  wire  line_1279_reset;
  wire  line_1279_valid;
  reg  line_1279_valid_reg;
  wire  _GEN_2123 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1280_clock;
  wire  line_1280_reset;
  wire  line_1280_valid;
  reg  line_1280_valid_reg;
  wire  _GEN_2124 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_3 : _GEN_2123; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1281_clock;
  wire  line_1281_reset;
  wire  line_1281_valid;
  reg  line_1281_valid_reg;
  wire  line_1282_clock;
  wire  line_1282_reset;
  wire  line_1282_valid;
  reg  line_1282_valid_reg;
  wire  line_1283_clock;
  wire  line_1283_reset;
  wire  line_1283_valid;
  reg  line_1283_valid_reg;
  wire  line_1284_clock;
  wire  line_1284_reset;
  wire  line_1284_valid;
  reg  line_1284_valid_reg;
  wire  line_1285_clock;
  wire  line_1285_reset;
  wire  line_1285_valid;
  reg  line_1285_valid_reg;
  wire  line_1286_clock;
  wire  line_1286_reset;
  wire  line_1286_valid;
  reg  line_1286_valid_reg;
  wire  line_1287_clock;
  wire  line_1287_reset;
  wire  line_1287_valid;
  reg  line_1287_valid_reg;
  wire  _GEN_2131 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1288_clock;
  wire  line_1288_reset;
  wire  line_1288_valid;
  reg  line_1288_valid_reg;
  wire  _GEN_2132 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_5 : _GEN_2131; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1289_clock;
  wire  line_1289_reset;
  wire  line_1289_valid;
  reg  line_1289_valid_reg;
  wire  line_1290_clock;
  wire  line_1290_reset;
  wire  line_1290_valid;
  reg  line_1290_valid_reg;
  wire  line_1291_clock;
  wire  line_1291_reset;
  wire  line_1291_valid;
  reg  line_1291_valid_reg;
  wire  line_1292_clock;
  wire  line_1292_reset;
  wire  line_1292_valid;
  reg  line_1292_valid_reg;
  wire  line_1293_clock;
  wire  line_1293_reset;
  wire  line_1293_valid;
  reg  line_1293_valid_reg;
  wire  line_1294_clock;
  wire  line_1294_reset;
  wire  line_1294_valid;
  reg  line_1294_valid_reg;
  wire  line_1295_clock;
  wire  line_1295_reset;
  wire  line_1295_valid;
  reg  line_1295_valid_reg;
  wire  _GEN_2139 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1296_clock;
  wire  line_1296_reset;
  wire  line_1296_valid;
  reg  line_1296_valid_reg;
  wire  _GEN_2140 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_7 : _GEN_2139; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1297_clock;
  wire  line_1297_reset;
  wire  line_1297_valid;
  reg  line_1297_valid_reg;
  wire  line_1298_clock;
  wire  line_1298_reset;
  wire  line_1298_valid;
  reg  line_1298_valid_reg;
  wire  line_1299_clock;
  wire  line_1299_reset;
  wire  line_1299_valid;
  reg  line_1299_valid_reg;
  wire  line_1300_clock;
  wire  line_1300_reset;
  wire  line_1300_valid;
  reg  line_1300_valid_reg;
  wire  line_1301_clock;
  wire  line_1301_reset;
  wire  line_1301_valid;
  reg  line_1301_valid_reg;
  wire  line_1302_clock;
  wire  line_1302_reset;
  wire  line_1302_valid;
  reg  line_1302_valid_reg;
  wire  line_1303_clock;
  wire  line_1303_reset;
  wire  line_1303_valid;
  reg  line_1303_valid_reg;
  wire  _GEN_2147 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1304_clock;
  wire  line_1304_reset;
  wire  line_1304_valid;
  reg  line_1304_valid_reg;
  wire  _GEN_2148 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_9 : _GEN_2147; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1305_clock;
  wire  line_1305_reset;
  wire  line_1305_valid;
  reg  line_1305_valid_reg;
  wire  line_1306_clock;
  wire  line_1306_reset;
  wire  line_1306_valid;
  reg  line_1306_valid_reg;
  wire  line_1307_clock;
  wire  line_1307_reset;
  wire  line_1307_valid;
  reg  line_1307_valid_reg;
  wire  line_1308_clock;
  wire  line_1308_reset;
  wire  line_1308_valid;
  reg  line_1308_valid_reg;
  wire  line_1309_clock;
  wire  line_1309_reset;
  wire  line_1309_valid;
  reg  line_1309_valid_reg;
  wire  line_1310_clock;
  wire  line_1310_reset;
  wire  line_1310_valid;
  reg  line_1310_valid_reg;
  wire  line_1311_clock;
  wire  line_1311_reset;
  wire  line_1311_valid;
  reg  line_1311_valid_reg;
  wire  _GEN_2155 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1312_clock;
  wire  line_1312_reset;
  wire  line_1312_valid;
  reg  line_1312_valid_reg;
  wire  _GEN_2156 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_11 : _GEN_2155; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1313_clock;
  wire  line_1313_reset;
  wire  line_1313_valid;
  reg  line_1313_valid_reg;
  wire  line_1314_clock;
  wire  line_1314_reset;
  wire  line_1314_valid;
  reg  line_1314_valid_reg;
  wire  line_1315_clock;
  wire  line_1315_reset;
  wire  line_1315_valid;
  reg  line_1315_valid_reg;
  wire  line_1316_clock;
  wire  line_1316_reset;
  wire  line_1316_valid;
  reg  line_1316_valid_reg;
  wire  line_1317_clock;
  wire  line_1317_reset;
  wire  line_1317_valid;
  reg  line_1317_valid_reg;
  wire  line_1318_clock;
  wire  line_1318_reset;
  wire  line_1318_valid;
  reg  line_1318_valid_reg;
  wire  line_1319_clock;
  wire  line_1319_reset;
  wire  line_1319_valid;
  reg  line_1319_valid_reg;
  wire  _GEN_2163 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_1 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1320_clock;
  wire  line_1320_reset;
  wire  line_1320_valid;
  reg  line_1320_valid_reg;
  wire  _GEN_2164 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_1 : _GEN_2163; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1321_clock;
  wire  line_1321_reset;
  wire  line_1321_valid;
  reg  line_1321_valid_reg;
  wire  line_1322_clock;
  wire  line_1322_reset;
  wire  line_1322_valid;
  reg  line_1322_valid_reg;
  wire  line_1323_clock;
  wire  line_1323_reset;
  wire  line_1323_valid;
  reg  line_1323_valid_reg;
  wire  _GEN_2167 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_2 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1324_clock;
  wire  line_1324_reset;
  wire  line_1324_valid;
  reg  line_1324_valid_reg;
  wire  _GEN_2168 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_2 : _GEN_2167; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1325_clock;
  wire  line_1325_reset;
  wire  line_1325_valid;
  reg  line_1325_valid_reg;
  wire  line_1326_clock;
  wire  line_1326_reset;
  wire  line_1326_valid;
  reg  line_1326_valid_reg;
  wire  line_1327_clock;
  wire  line_1327_reset;
  wire  line_1327_valid;
  reg  line_1327_valid_reg;
  wire  line_1328_clock;
  wire  line_1328_reset;
  wire  line_1328_valid;
  reg  line_1328_valid_reg;
  wire  line_1329_clock;
  wire  line_1329_reset;
  wire  line_1329_valid;
  reg  line_1329_valid_reg;
  wire  line_1330_clock;
  wire  line_1330_reset;
  wire  line_1330_valid;
  reg  line_1330_valid_reg;
  wire  line_1331_clock;
  wire  line_1331_reset;
  wire  line_1331_valid;
  reg  line_1331_valid_reg;
  wire  line_1332_clock;
  wire  line_1332_reset;
  wire  line_1332_valid;
  reg  line_1332_valid_reg;
  wire  line_1333_clock;
  wire  line_1333_reset;
  wire  line_1333_valid;
  reg  line_1333_valid_reg;
  wire  line_1334_clock;
  wire  line_1334_reset;
  wire  line_1334_valid;
  reg  line_1334_valid_reg;
  wire  line_1335_clock;
  wire  line_1335_reset;
  wire  line_1335_valid;
  reg  line_1335_valid_reg;
  wire  line_1336_clock;
  wire  line_1336_reset;
  wire  line_1336_valid;
  reg  line_1336_valid_reg;
  wire  line_1337_clock;
  wire  line_1337_reset;
  wire  line_1337_valid;
  reg  line_1337_valid_reg;
  wire  line_1338_clock;
  wire  line_1338_reset;
  wire  line_1338_valid;
  reg  line_1338_valid_reg;
  wire  line_1339_clock;
  wire  line_1339_reset;
  wire  line_1339_valid;
  reg  line_1339_valid_reg;
  wire  line_1340_clock;
  wire  line_1340_reset;
  wire  line_1340_valid;
  reg  line_1340_valid_reg;
  wire  line_1341_clock;
  wire  line_1341_reset;
  wire  line_1341_valid;
  reg  line_1341_valid_reg;
  wire  line_1342_clock;
  wire  line_1342_reset;
  wire  line_1342_valid;
  reg  line_1342_valid_reg;
  wire  line_1343_clock;
  wire  line_1343_reset;
  wire  line_1343_valid;
  reg  line_1343_valid_reg;
  wire  line_1344_clock;
  wire  line_1344_reset;
  wire  line_1344_valid;
  reg  line_1344_valid_reg;
  wire  line_1345_clock;
  wire  line_1345_reset;
  wire  line_1345_valid;
  reg  line_1345_valid_reg;
  wire  line_1346_clock;
  wire  line_1346_reset;
  wire  line_1346_valid;
  reg  line_1346_valid_reg;
  wire  line_1347_clock;
  wire  line_1347_reset;
  wire  line_1347_valid;
  reg  line_1347_valid_reg;
  wire  line_1348_clock;
  wire  line_1348_reset;
  wire  line_1348_valid;
  reg  line_1348_valid_reg;
  wire  line_1349_clock;
  wire  line_1349_reset;
  wire  line_1349_valid;
  reg  line_1349_valid_reg;
  wire  line_1350_clock;
  wire  line_1350_reset;
  wire  line_1350_valid;
  reg  line_1350_valid_reg;
  wire  line_1351_clock;
  wire  line_1351_reset;
  wire  line_1351_valid;
  reg  line_1351_valid_reg;
  wire  line_1352_clock;
  wire  line_1352_reset;
  wire  line_1352_valid;
  reg  line_1352_valid_reg;
  wire  line_1353_clock;
  wire  line_1353_reset;
  wire  line_1353_valid;
  reg  line_1353_valid_reg;
  wire  line_1354_clock;
  wire  line_1354_reset;
  wire  line_1354_valid;
  reg  line_1354_valid_reg;
  wire  line_1355_clock;
  wire  line_1355_reset;
  wire  line_1355_valid;
  reg  line_1355_valid_reg;
  wire  line_1356_clock;
  wire  line_1356_reset;
  wire  line_1356_valid;
  reg  line_1356_valid_reg;
  wire  line_1357_clock;
  wire  line_1357_reset;
  wire  line_1357_valid;
  reg  line_1357_valid_reg;
  wire  line_1358_clock;
  wire  line_1358_reset;
  wire  line_1358_valid;
  reg  line_1358_valid_reg;
  wire  line_1359_clock;
  wire  line_1359_reset;
  wire  line_1359_valid;
  reg  line_1359_valid_reg;
  wire  line_1360_clock;
  wire  line_1360_reset;
  wire  line_1360_valid;
  reg  line_1360_valid_reg;
  wire  line_1361_clock;
  wire  line_1361_reset;
  wire  line_1361_valid;
  reg  line_1361_valid_reg;
  wire  line_1362_clock;
  wire  line_1362_reset;
  wire  line_1362_valid;
  reg  line_1362_valid_reg;
  wire  line_1363_clock;
  wire  line_1363_reset;
  wire  line_1363_valid;
  reg  line_1363_valid_reg;
  wire  _GEN_2207 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_12 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1364_clock;
  wire  line_1364_reset;
  wire  line_1364_valid;
  reg  line_1364_valid_reg;
  wire  _GEN_2208 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_12 : _GEN_2207; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1365_clock;
  wire  line_1365_reset;
  wire  line_1365_valid;
  reg  line_1365_valid_reg;
  wire  line_1366_clock;
  wire  line_1366_reset;
  wire  line_1366_valid;
  reg  line_1366_valid_reg;
  wire  line_1367_clock;
  wire  line_1367_reset;
  wire  line_1367_valid;
  reg  line_1367_valid_reg;
  wire  line_1368_clock;
  wire  line_1368_reset;
  wire  line_1368_valid;
  reg  line_1368_valid_reg;
  wire  line_1369_clock;
  wire  line_1369_reset;
  wire  line_1369_valid;
  reg  line_1369_valid_reg;
  wire  line_1370_clock;
  wire  line_1370_reset;
  wire  line_1370_valid;
  reg  line_1370_valid_reg;
  wire  line_1371_clock;
  wire  line_1371_reset;
  wire  line_1371_valid;
  reg  line_1371_valid_reg;
  wire  line_1372_clock;
  wire  line_1372_reset;
  wire  line_1372_valid;
  reg  line_1372_valid_reg;
  wire  line_1373_clock;
  wire  line_1373_reset;
  wire  line_1373_valid;
  reg  line_1373_valid_reg;
  wire  line_1374_clock;
  wire  line_1374_reset;
  wire  line_1374_valid;
  reg  line_1374_valid_reg;
  wire  line_1375_clock;
  wire  line_1375_reset;
  wire  line_1375_valid;
  reg  line_1375_valid_reg;
  wire  line_1376_clock;
  wire  line_1376_reset;
  wire  line_1376_valid;
  reg  line_1376_valid_reg;
  wire  line_1377_clock;
  wire  line_1377_reset;
  wire  line_1377_valid;
  reg  line_1377_valid_reg;
  wire  line_1378_clock;
  wire  line_1378_reset;
  wire  line_1378_valid;
  reg  line_1378_valid_reg;
  wire  line_1379_clock;
  wire  line_1379_reset;
  wire  line_1379_valid;
  reg  line_1379_valid_reg;
  wire  line_1380_clock;
  wire  line_1380_reset;
  wire  line_1380_valid;
  reg  line_1380_valid_reg;
  wire  line_1381_clock;
  wire  line_1381_reset;
  wire  line_1381_valid;
  reg  line_1381_valid_reg;
  wire  line_1382_clock;
  wire  line_1382_reset;
  wire  line_1382_valid;
  reg  line_1382_valid_reg;
  wire  line_1383_clock;
  wire  line_1383_reset;
  wire  line_1383_valid;
  reg  line_1383_valid_reg;
  wire  line_1384_clock;
  wire  line_1384_reset;
  wire  line_1384_valid;
  reg  line_1384_valid_reg;
  wire  line_1385_clock;
  wire  line_1385_reset;
  wire  line_1385_valid;
  reg  line_1385_valid_reg;
  wire  line_1386_clock;
  wire  line_1386_reset;
  wire  line_1386_valid;
  reg  line_1386_valid_reg;
  wire  line_1387_clock;
  wire  line_1387_reset;
  wire  line_1387_valid;
  reg  line_1387_valid_reg;
  wire  line_1388_clock;
  wire  line_1388_reset;
  wire  line_1388_valid;
  reg  line_1388_valid_reg;
  wire  line_1389_clock;
  wire  line_1389_reset;
  wire  line_1389_valid;
  reg  line_1389_valid_reg;
  wire  line_1390_clock;
  wire  line_1390_reset;
  wire  line_1390_valid;
  reg  line_1390_valid_reg;
  wire  line_1391_clock;
  wire  line_1391_reset;
  wire  line_1391_valid;
  reg  line_1391_valid_reg;
  wire [38:0] _GEN_2235 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1392_clock;
  wire  line_1392_reset;
  wire  line_1392_valid;
  reg  line_1392_valid_reg;
  wire [38:0] _GEN_2236 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pnpc : _GEN_2235; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1393_clock;
  wire  line_1393_reset;
  wire  line_1393_valid;
  reg  line_1393_valid_reg;
  wire  line_1394_clock;
  wire  line_1394_reset;
  wire  line_1394_valid;
  reg  line_1394_valid_reg;
  wire  line_1395_clock;
  wire  line_1395_reset;
  wire  line_1395_valid;
  reg  line_1395_valid_reg;
  wire [38:0] _GEN_2239 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1396_clock;
  wire  line_1396_reset;
  wire  line_1396_valid;
  reg  line_1396_valid_reg;
  wire [38:0] _GEN_2240 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pc : _GEN_2239; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1397_clock;
  wire  line_1397_reset;
  wire  line_1397_valid;
  reg  line_1397_valid_reg;
  wire  line_1398_clock;
  wire  line_1398_reset;
  wire  line_1398_valid;
  reg  line_1398_valid_reg;
  wire  line_1399_clock;
  wire  line_1399_reset;
  wire  line_1399_valid;
  reg  line_1399_valid_reg;
  wire [63:0] _GEN_2243 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1400_clock;
  wire  line_1400_reset;
  wire  line_1400_valid;
  reg  line_1400_valid_reg;
  wire [63:0] _GEN_2244 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_instr : _GEN_2243; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  line_1401_clock;
  wire  line_1401_reset;
  wire  line_1401_valid;
  reg  line_1401_valid_reg;
  wire [1:0] deq2_StartIndex = ringBufferTail + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 59:42]
  wire  line_1402_clock;
  wire  line_1402_reset;
  wire  line_1402_valid;
  reg  line_1402_valid_reg;
  wire  line_1403_clock;
  wire  line_1403_reset;
  wire  line_1403_valid;
  reg  line_1403_valid_reg;
  wire  line_1404_clock;
  wire  line_1404_reset;
  wire  line_1404_valid;
  reg  line_1404_valid_reg;
  wire  line_1405_clock;
  wire  line_1405_reset;
  wire  line_1405_valid;
  reg  line_1405_valid_reg;
  wire  line_1406_clock;
  wire  line_1406_reset;
  wire  line_1406_valid;
  reg  line_1406_valid_reg;
  wire  line_1407_clock;
  wire  line_1407_reset;
  wire  line_1407_valid;
  reg  line_1407_valid_reg;
  wire  line_1408_clock;
  wire  line_1408_reset;
  wire  line_1408_valid;
  reg  line_1408_valid_reg;
  wire  line_1409_clock;
  wire  line_1409_reset;
  wire  line_1409_valid;
  reg  line_1409_valid_reg;
  wire  line_1410_clock;
  wire  line_1410_reset;
  wire  line_1410_valid;
  reg  line_1410_valid_reg;
  wire  line_1411_clock;
  wire  line_1411_reset;
  wire  line_1411_valid;
  reg  line_1411_valid_reg;
  wire  line_1412_clock;
  wire  line_1412_reset;
  wire  line_1412_valid;
  reg  line_1412_valid_reg;
  wire  line_1413_clock;
  wire  line_1413_reset;
  wire  line_1413_valid;
  reg  line_1413_valid_reg;
  wire  line_1414_clock;
  wire  line_1414_reset;
  wire  line_1414_valid;
  reg  line_1414_valid_reg;
  wire  line_1415_clock;
  wire  line_1415_reset;
  wire  line_1415_valid;
  reg  line_1415_valid_reg;
  wire  line_1416_clock;
  wire  line_1416_reset;
  wire  line_1416_valid;
  reg  line_1416_valid_reg;
  wire  line_1417_clock;
  wire  line_1417_reset;
  wire  line_1417_valid;
  reg  line_1417_valid_reg;
  wire  line_1418_clock;
  wire  line_1418_reset;
  wire  line_1418_valid;
  reg  line_1418_valid_reg;
  wire  line_1419_clock;
  wire  line_1419_reset;
  wire  line_1419_valid;
  reg  line_1419_valid_reg;
  wire  line_1420_clock;
  wire  line_1420_reset;
  wire  line_1420_valid;
  reg  line_1420_valid_reg;
  wire  line_1421_clock;
  wire  line_1421_reset;
  wire  line_1421_valid;
  reg  line_1421_valid_reg;
  wire  line_1422_clock;
  wire  line_1422_reset;
  wire  line_1422_valid;
  reg  line_1422_valid_reg;
  wire  line_1423_clock;
  wire  line_1423_reset;
  wire  line_1423_valid;
  reg  line_1423_valid_reg;
  wire  line_1424_clock;
  wire  line_1424_reset;
  wire  line_1424_valid;
  reg  line_1424_valid_reg;
  wire  line_1425_clock;
  wire  line_1425_reset;
  wire  line_1425_valid;
  reg  line_1425_valid_reg;
  wire  line_1426_clock;
  wire  line_1426_reset;
  wire  line_1426_valid;
  reg  line_1426_valid_reg;
  wire  line_1427_clock;
  wire  line_1427_reset;
  wire  line_1427_valid;
  reg  line_1427_valid_reg;
  wire  line_1428_clock;
  wire  line_1428_reset;
  wire  line_1428_valid;
  reg  line_1428_valid_reg;
  wire  line_1429_clock;
  wire  line_1429_reset;
  wire  line_1429_valid;
  reg  line_1429_valid_reg;
  wire  line_1430_clock;
  wire  line_1430_reset;
  wire  line_1430_valid;
  reg  line_1430_valid_reg;
  wire  line_1431_clock;
  wire  line_1431_reset;
  wire  line_1431_valid;
  reg  line_1431_valid_reg;
  wire  line_1432_clock;
  wire  line_1432_reset;
  wire  line_1432_valid;
  reg  line_1432_valid_reg;
  wire  line_1433_clock;
  wire  line_1433_reset;
  wire  line_1433_valid;
  reg  line_1433_valid_reg;
  wire  line_1434_clock;
  wire  line_1434_reset;
  wire  line_1434_valid;
  reg  line_1434_valid_reg;
  wire  line_1435_clock;
  wire  line_1435_reset;
  wire  line_1435_valid;
  reg  line_1435_valid_reg;
  wire  line_1436_clock;
  wire  line_1436_reset;
  wire  line_1436_valid;
  reg  line_1436_valid_reg;
  wire  line_1437_clock;
  wire  line_1437_reset;
  wire  line_1437_valid;
  reg  line_1437_valid_reg;
  wire  line_1438_clock;
  wire  line_1438_reset;
  wire  line_1438_valid;
  reg  line_1438_valid_reg;
  wire  line_1439_clock;
  wire  line_1439_reset;
  wire  line_1439_valid;
  reg  line_1439_valid_reg;
  wire  line_1440_clock;
  wire  line_1440_reset;
  wire  line_1440_valid;
  reg  line_1440_valid_reg;
  wire  line_1441_clock;
  wire  line_1441_reset;
  wire  line_1441_valid;
  reg  line_1441_valid_reg;
  wire  line_1442_clock;
  wire  line_1442_reset;
  wire  line_1442_valid;
  reg  line_1442_valid_reg;
  wire  line_1443_clock;
  wire  line_1443_reset;
  wire  line_1443_valid;
  reg  line_1443_valid_reg;
  wire  line_1444_clock;
  wire  line_1444_reset;
  wire  line_1444_valid;
  reg  line_1444_valid_reg;
  wire  line_1445_clock;
  wire  line_1445_reset;
  wire  line_1445_valid;
  reg  line_1445_valid_reg;
  wire  line_1446_clock;
  wire  line_1446_reset;
  wire  line_1446_valid;
  reg  line_1446_valid_reg;
  wire  line_1447_clock;
  wire  line_1447_reset;
  wire  line_1447_valid;
  reg  line_1447_valid_reg;
  wire  line_1448_clock;
  wire  line_1448_reset;
  wire  line_1448_valid;
  reg  line_1448_valid_reg;
  wire  line_1449_clock;
  wire  line_1449_reset;
  wire  line_1449_valid;
  reg  line_1449_valid_reg;
  wire  line_1450_clock;
  wire  line_1450_reset;
  wire  line_1450_valid;
  reg  line_1450_valid_reg;
  wire  line_1451_clock;
  wire  line_1451_reset;
  wire  line_1451_valid;
  reg  line_1451_valid_reg;
  wire  line_1452_clock;
  wire  line_1452_reset;
  wire  line_1452_valid;
  reg  line_1452_valid_reg;
  wire  line_1453_clock;
  wire  line_1453_reset;
  wire  line_1453_valid;
  reg  line_1453_valid_reg;
  wire  line_1454_clock;
  wire  line_1454_reset;
  wire  line_1454_valid;
  reg  line_1454_valid_reg;
  wire  line_1455_clock;
  wire  line_1455_reset;
  wire  line_1455_valid;
  reg  line_1455_valid_reg;
  wire  line_1456_clock;
  wire  line_1456_reset;
  wire  line_1456_valid;
  reg  line_1456_valid_reg;
  wire  line_1457_clock;
  wire  line_1457_reset;
  wire  line_1457_valid;
  reg  line_1457_valid_reg;
  wire  line_1458_clock;
  wire  line_1458_reset;
  wire  line_1458_valid;
  reg  line_1458_valid_reg;
  wire  line_1459_clock;
  wire  line_1459_reset;
  wire  line_1459_valid;
  reg  line_1459_valid_reg;
  wire  line_1460_clock;
  wire  line_1460_reset;
  wire  line_1460_valid;
  reg  line_1460_valid_reg;
  wire  line_1461_clock;
  wire  line_1461_reset;
  wire  line_1461_valid;
  reg  line_1461_valid_reg;
  wire  line_1462_clock;
  wire  line_1462_reset;
  wire  line_1462_valid;
  reg  line_1462_valid_reg;
  wire  line_1463_clock;
  wire  line_1463_reset;
  wire  line_1463_valid;
  reg  line_1463_valid_reg;
  wire  line_1464_clock;
  wire  line_1464_reset;
  wire  line_1464_valid;
  reg  line_1464_valid_reg;
  wire  line_1465_clock;
  wire  line_1465_reset;
  wire  line_1465_valid;
  reg  line_1465_valid_reg;
  wire  line_1466_clock;
  wire  line_1466_reset;
  wire  line_1466_valid;
  reg  line_1466_valid_reg;
  wire  line_1467_clock;
  wire  line_1467_reset;
  wire  line_1467_valid;
  reg  line_1467_valid_reg;
  wire  line_1468_clock;
  wire  line_1468_reset;
  wire  line_1468_valid;
  reg  line_1468_valid_reg;
  wire  line_1469_clock;
  wire  line_1469_reset;
  wire  line_1469_valid;
  reg  line_1469_valid_reg;
  wire  line_1470_clock;
  wire  line_1470_reset;
  wire  line_1470_valid;
  reg  line_1470_valid_reg;
  wire  line_1471_clock;
  wire  line_1471_reset;
  wire  line_1471_valid;
  reg  line_1471_valid_reg;
  wire  line_1472_clock;
  wire  line_1472_reset;
  wire  line_1472_valid;
  reg  line_1472_valid_reg;
  wire  line_1473_clock;
  wire  line_1473_reset;
  wire  line_1473_valid;
  reg  line_1473_valid_reg;
  wire  line_1474_clock;
  wire  line_1474_reset;
  wire  line_1474_valid;
  reg  line_1474_valid_reg;
  wire  line_1475_clock;
  wire  line_1475_reset;
  wire  line_1475_valid;
  reg  line_1475_valid_reg;
  wire  line_1476_clock;
  wire  line_1476_reset;
  wire  line_1476_valid;
  reg  line_1476_valid_reg;
  wire  line_1477_clock;
  wire  line_1477_reset;
  wire  line_1477_valid;
  reg  line_1477_valid_reg;
  wire  line_1478_clock;
  wire  line_1478_reset;
  wire  line_1478_valid;
  reg  line_1478_valid_reg;
  wire  line_1479_clock;
  wire  line_1479_reset;
  wire  line_1479_valid;
  reg  line_1479_valid_reg;
  wire  line_1480_clock;
  wire  line_1480_reset;
  wire  line_1480_valid;
  reg  line_1480_valid_reg;
  wire  line_1481_clock;
  wire  line_1481_reset;
  wire  line_1481_valid;
  reg  line_1481_valid_reg;
  wire  line_1482_clock;
  wire  line_1482_reset;
  wire  line_1482_valid;
  reg  line_1482_valid_reg;
  wire  line_1483_clock;
  wire  line_1483_reset;
  wire  line_1483_valid;
  reg  line_1483_valid_reg;
  wire  line_1484_clock;
  wire  line_1484_reset;
  wire  line_1484_valid;
  reg  line_1484_valid_reg;
  wire  line_1485_clock;
  wire  line_1485_reset;
  wire  line_1485_valid;
  reg  line_1485_valid_reg;
  wire  line_1486_clock;
  wire  line_1486_reset;
  wire  line_1486_valid;
  reg  line_1486_valid_reg;
  wire  line_1487_clock;
  wire  line_1487_reset;
  wire  line_1487_valid;
  reg  line_1487_valid_reg;
  wire  line_1488_clock;
  wire  line_1488_reset;
  wire  line_1488_valid;
  reg  line_1488_valid_reg;
  wire  line_1489_clock;
  wire  line_1489_reset;
  wire  line_1489_valid;
  reg  line_1489_valid_reg;
  wire  line_1490_clock;
  wire  line_1490_reset;
  wire  line_1490_valid;
  reg  line_1490_valid_reg;
  wire  line_1491_clock;
  wire  line_1491_reset;
  wire  line_1491_valid;
  reg  line_1491_valid_reg;
  wire  line_1492_clock;
  wire  line_1492_reset;
  wire  line_1492_valid;
  reg  line_1492_valid_reg;
  wire  line_1493_clock;
  wire  line_1493_reset;
  wire  line_1493_valid;
  reg  line_1493_valid_reg;
  wire  line_1494_clock;
  wire  line_1494_reset;
  wire  line_1494_valid;
  reg  line_1494_valid_reg;
  wire  line_1495_clock;
  wire  line_1495_reset;
  wire  line_1495_valid;
  reg  line_1495_valid_reg;
  wire  line_1496_clock;
  wire  line_1496_reset;
  wire  line_1496_valid;
  reg  line_1496_valid_reg;
  wire  line_1497_clock;
  wire  line_1497_reset;
  wire  line_1497_valid;
  reg  line_1497_valid_reg;
  wire  line_1498_clock;
  wire  line_1498_reset;
  wire  line_1498_valid;
  reg  line_1498_valid_reg;
  wire  line_1499_clock;
  wire  line_1499_reset;
  wire  line_1499_valid;
  reg  line_1499_valid_reg;
  wire  line_1500_clock;
  wire  line_1500_reset;
  wire  line_1500_valid;
  reg  line_1500_valid_reg;
  wire  line_1501_clock;
  wire  line_1501_reset;
  wire  line_1501_valid;
  reg  line_1501_valid_reg;
  wire  line_1502_clock;
  wire  line_1502_reset;
  wire  line_1502_valid;
  reg  line_1502_valid_reg;
  wire  line_1503_clock;
  wire  line_1503_reset;
  wire  line_1503_valid;
  reg  line_1503_valid_reg;
  wire  line_1504_clock;
  wire  line_1504_reset;
  wire  line_1504_valid;
  reg  line_1504_valid_reg;
  wire  line_1505_clock;
  wire  line_1505_reset;
  wire  line_1505_valid;
  reg  line_1505_valid_reg;
  wire  line_1506_clock;
  wire  line_1506_reset;
  wire  line_1506_valid;
  reg  line_1506_valid_reg;
  wire  line_1507_clock;
  wire  line_1507_reset;
  wire  line_1507_valid;
  reg  line_1507_valid_reg;
  wire  line_1508_clock;
  wire  line_1508_reset;
  wire  line_1508_valid;
  reg  line_1508_valid_reg;
  wire  line_1509_clock;
  wire  line_1509_reset;
  wire  line_1509_valid;
  reg  line_1509_valid_reg;
  wire  line_1510_clock;
  wire  line_1510_reset;
  wire  line_1510_valid;
  reg  line_1510_valid_reg;
  wire  line_1511_clock;
  wire  line_1511_reset;
  wire  line_1511_valid;
  reg  line_1511_valid_reg;
  wire  line_1512_clock;
  wire  line_1512_reset;
  wire  line_1512_valid;
  reg  line_1512_valid_reg;
  wire  line_1513_clock;
  wire  line_1513_reset;
  wire  line_1513_valid;
  reg  line_1513_valid_reg;
  wire  line_1514_clock;
  wire  line_1514_reset;
  wire  line_1514_valid;
  reg  line_1514_valid_reg;
  wire  line_1515_clock;
  wire  line_1515_reset;
  wire  line_1515_valid;
  reg  line_1515_valid_reg;
  wire  line_1516_clock;
  wire  line_1516_reset;
  wire  line_1516_valid;
  reg  line_1516_valid_reg;
  wire  line_1517_clock;
  wire  line_1517_reset;
  wire  line_1517_valid;
  reg  line_1517_valid_reg;
  wire  line_1518_clock;
  wire  line_1518_reset;
  wire  line_1518_valid;
  reg  line_1518_valid_reg;
  wire  line_1519_clock;
  wire  line_1519_reset;
  wire  line_1519_valid;
  reg  line_1519_valid_reg;
  wire  line_1520_clock;
  wire  line_1520_reset;
  wire  line_1520_valid;
  reg  line_1520_valid_reg;
  wire  line_1521_clock;
  wire  line_1521_reset;
  wire  line_1521_valid;
  reg  line_1521_valid_reg;
  wire  line_1522_clock;
  wire  line_1522_reset;
  wire  line_1522_valid;
  reg  line_1522_valid_reg;
  wire  line_1523_clock;
  wire  line_1523_reset;
  wire  line_1523_valid;
  reg  line_1523_valid_reg;
  wire  line_1524_clock;
  wire  line_1524_reset;
  wire  line_1524_valid;
  reg  line_1524_valid_reg;
  wire  line_1525_clock;
  wire  line_1525_reset;
  wire  line_1525_valid;
  reg  line_1525_valid_reg;
  wire  line_1526_clock;
  wire  line_1526_reset;
  wire  line_1526_valid;
  reg  line_1526_valid_reg;
  wire  line_1527_clock;
  wire  line_1527_reset;
  wire  line_1527_valid;
  reg  line_1527_valid_reg;
  wire  line_1528_clock;
  wire  line_1528_reset;
  wire  line_1528_valid;
  reg  line_1528_valid_reg;
  wire  line_1529_clock;
  wire  line_1529_reset;
  wire  line_1529_valid;
  reg  line_1529_valid_reg;
  wire  line_1530_clock;
  wire  line_1530_reset;
  wire  line_1530_valid;
  reg  line_1530_valid_reg;
  wire  line_1531_clock;
  wire  line_1531_reset;
  wire  line_1531_valid;
  reg  line_1531_valid_reg;
  wire  line_1532_clock;
  wire  line_1532_reset;
  wire  line_1532_valid;
  reg  line_1532_valid_reg;
  wire  line_1533_clock;
  wire  line_1533_reset;
  wire  line_1533_valid;
  reg  line_1533_valid_reg;
  wire  line_1534_clock;
  wire  line_1534_reset;
  wire  line_1534_valid;
  reg  line_1534_valid_reg;
  wire  line_1535_clock;
  wire  line_1535_reset;
  wire  line_1535_valid;
  reg  line_1535_valid_reg;
  wire  line_1536_clock;
  wire  line_1536_reset;
  wire  line_1536_valid;
  reg  line_1536_valid_reg;
  wire  line_1537_clock;
  wire  line_1537_reset;
  wire  line_1537_valid;
  reg  line_1537_valid_reg;
  wire  line_1538_clock;
  wire  line_1538_reset;
  wire  line_1538_valid;
  reg  line_1538_valid_reg;
  wire  line_1539_clock;
  wire  line_1539_reset;
  wire  line_1539_valid;
  reg  line_1539_valid_reg;
  wire  line_1540_clock;
  wire  line_1540_reset;
  wire  line_1540_valid;
  reg  line_1540_valid_reg;
  wire  line_1541_clock;
  wire  line_1541_reset;
  wire  line_1541_valid;
  reg  line_1541_valid_reg;
  wire  line_1542_clock;
  wire  line_1542_reset;
  wire  line_1542_valid;
  reg  line_1542_valid_reg;
  wire  line_1543_clock;
  wire  line_1543_reset;
  wire  line_1543_valid;
  reg  line_1543_valid_reg;
  wire  line_1544_clock;
  wire  line_1544_reset;
  wire  line_1544_valid;
  reg  line_1544_valid_reg;
  wire  line_1545_clock;
  wire  line_1545_reset;
  wire  line_1545_valid;
  reg  line_1545_valid_reg;
  wire  line_1546_clock;
  wire  line_1546_reset;
  wire  line_1546_valid;
  reg  line_1546_valid_reg;
  wire  line_1547_clock;
  wire  line_1547_reset;
  wire  line_1547_valid;
  reg  line_1547_valid_reg;
  wire  line_1548_clock;
  wire  line_1548_reset;
  wire  line_1548_valid;
  reg  line_1548_valid_reg;
  wire  line_1549_clock;
  wire  line_1549_reset;
  wire  line_1549_valid;
  reg  line_1549_valid_reg;
  wire  line_1550_clock;
  wire  line_1550_reset;
  wire  line_1550_valid;
  reg  line_1550_valid_reg;
  wire  line_1551_clock;
  wire  line_1551_reset;
  wire  line_1551_valid;
  reg  line_1551_valid_reg;
  wire  line_1552_clock;
  wire  line_1552_reset;
  wire  line_1552_valid;
  reg  line_1552_valid_reg;
  wire  line_1553_clock;
  wire  line_1553_reset;
  wire  line_1553_valid;
  reg  line_1553_valid_reg;
  wire  line_1554_clock;
  wire  line_1554_reset;
  wire  line_1554_valid;
  reg  line_1554_valid_reg;
  wire  line_1555_clock;
  wire  line_1555_reset;
  wire  line_1555_valid;
  reg  line_1555_valid_reg;
  wire  line_1556_clock;
  wire  line_1556_reset;
  wire  line_1556_valid;
  reg  line_1556_valid_reg;
  wire  line_1557_clock;
  wire  line_1557_reset;
  wire  line_1557_valid;
  reg  line_1557_valid_reg;
  wire  line_1558_clock;
  wire  line_1558_reset;
  wire  line_1558_valid;
  reg  line_1558_valid_reg;
  wire  line_1559_clock;
  wire  line_1559_reset;
  wire  line_1559_valid;
  reg  line_1559_valid_reg;
  wire  line_1560_clock;
  wire  line_1560_reset;
  wire  line_1560_valid;
  reg  line_1560_valid_reg;
  wire  line_1561_clock;
  wire  line_1561_reset;
  wire  line_1561_valid;
  reg  line_1561_valid_reg;
  wire  line_1562_clock;
  wire  line_1562_reset;
  wire  line_1562_valid;
  reg  line_1562_valid_reg;
  wire  line_1563_clock;
  wire  line_1563_reset;
  wire  line_1563_valid;
  reg  line_1563_valid_reg;
  wire  line_1564_clock;
  wire  line_1564_reset;
  wire  line_1564_valid;
  reg  line_1564_valid_reg;
  wire  line_1565_clock;
  wire  line_1565_reset;
  wire  line_1565_valid;
  reg  line_1565_valid_reg;
  wire  line_1566_clock;
  wire  line_1566_reset;
  wire  line_1566_valid;
  reg  line_1566_valid_reg;
  wire  line_1567_clock;
  wire  line_1567_reset;
  wire  line_1567_valid;
  reg  line_1567_valid_reg;
  wire  line_1568_clock;
  wire  line_1568_reset;
  wire  line_1568_valid;
  reg  line_1568_valid_reg;
  wire  line_1569_clock;
  wire  line_1569_reset;
  wire  line_1569_valid;
  reg  line_1569_valid_reg;
  wire  line_1570_clock;
  wire  line_1570_reset;
  wire  line_1570_valid;
  reg  line_1570_valid_reg;
  wire  line_1571_clock;
  wire  line_1571_reset;
  wire  line_1571_valid;
  reg  line_1571_valid_reg;
  wire  line_1572_clock;
  wire  line_1572_reset;
  wire  line_1572_valid;
  reg  line_1572_valid_reg;
  wire  line_1573_clock;
  wire  line_1573_reset;
  wire  line_1573_valid;
  reg  line_1573_valid_reg;
  wire  line_1574_clock;
  wire  line_1574_reset;
  wire  line_1574_valid;
  reg  line_1574_valid_reg;
  wire  line_1575_clock;
  wire  line_1575_reset;
  wire  line_1575_valid;
  reg  line_1575_valid_reg;
  wire  line_1576_clock;
  wire  line_1576_reset;
  wire  line_1576_valid;
  reg  line_1576_valid_reg;
  wire  line_1577_clock;
  wire  line_1577_reset;
  wire  line_1577_valid;
  reg  line_1577_valid_reg;
  wire  line_1578_clock;
  wire  line_1578_reset;
  wire  line_1578_valid;
  reg  line_1578_valid_reg;
  wire  line_1579_clock;
  wire  line_1579_reset;
  wire  line_1579_valid;
  reg  line_1579_valid_reg;
  wire  line_1580_clock;
  wire  line_1580_reset;
  wire  line_1580_valid;
  reg  line_1580_valid_reg;
  wire  line_1581_clock;
  wire  line_1581_reset;
  wire  line_1581_valid;
  reg  line_1581_valid_reg;
  wire  line_1582_clock;
  wire  line_1582_reset;
  wire  line_1582_valid;
  reg  line_1582_valid_reg;
  wire  line_1583_clock;
  wire  line_1583_reset;
  wire  line_1583_valid;
  reg  line_1583_valid_reg;
  wire  line_1584_clock;
  wire  line_1584_reset;
  wire  line_1584_valid;
  reg  line_1584_valid_reg;
  wire  line_1585_clock;
  wire  line_1585_reset;
  wire  line_1585_valid;
  reg  line_1585_valid_reg;
  wire  line_1586_clock;
  wire  line_1586_reset;
  wire  line_1586_valid;
  reg  line_1586_valid_reg;
  wire  line_1587_clock;
  wire  line_1587_reset;
  wire  line_1587_valid;
  reg  line_1587_valid_reg;
  wire  line_1588_clock;
  wire  line_1588_reset;
  wire  line_1588_valid;
  reg  line_1588_valid_reg;
  wire  line_1589_clock;
  wire  line_1589_reset;
  wire  line_1589_valid;
  reg  line_1589_valid_reg;
  wire  line_1590_clock;
  wire  line_1590_reset;
  wire  line_1590_valid;
  reg  line_1590_valid_reg;
  wire  line_1591_clock;
  wire  line_1591_reset;
  wire  line_1591_valid;
  reg  line_1591_valid_reg;
  wire  line_1592_clock;
  wire  line_1592_reset;
  wire  line_1592_valid;
  reg  line_1592_valid_reg;
  wire  line_1593_clock;
  wire  line_1593_reset;
  wire  line_1593_valid;
  reg  line_1593_valid_reg;
  wire  line_1594_clock;
  wire  line_1594_reset;
  wire  line_1594_valid;
  reg  line_1594_valid_reg;
  wire  line_1595_clock;
  wire  line_1595_reset;
  wire  line_1595_valid;
  reg  line_1595_valid_reg;
  wire  line_1596_clock;
  wire  line_1596_reset;
  wire  line_1596_valid;
  reg  line_1596_valid_reg;
  wire  line_1597_clock;
  wire  line_1597_reset;
  wire  line_1597_valid;
  reg  line_1597_valid_reg;
  wire  line_1598_clock;
  wire  line_1598_reset;
  wire  line_1598_valid;
  reg  line_1598_valid_reg;
  wire  line_1599_clock;
  wire  line_1599_reset;
  wire  line_1599_valid;
  reg  line_1599_valid_reg;
  wire  line_1600_clock;
  wire  line_1600_reset;
  wire  line_1600_valid;
  reg  line_1600_valid_reg;
  wire  line_1601_clock;
  wire  line_1601_reset;
  wire  line_1601_valid;
  reg  line_1601_valid_reg;
  wire  line_1602_clock;
  wire  line_1602_reset;
  wire  line_1602_valid;
  reg  line_1602_valid_reg;
  wire  line_1603_clock;
  wire  line_1603_reset;
  wire  line_1603_valid;
  reg  line_1603_valid_reg;
  wire  line_1604_clock;
  wire  line_1604_reset;
  wire  line_1604_valid;
  reg  line_1604_valid_reg;
  wire  line_1605_clock;
  wire  line_1605_reset;
  wire  line_1605_valid;
  reg  line_1605_valid_reg;
  wire  line_1606_clock;
  wire  line_1606_reset;
  wire  line_1606_valid;
  reg  line_1606_valid_reg;
  wire  line_1607_clock;
  wire  line_1607_reset;
  wire  line_1607_valid;
  reg  line_1607_valid_reg;
  wire  line_1608_clock;
  wire  line_1608_reset;
  wire  line_1608_valid;
  reg  line_1608_valid_reg;
  wire  line_1609_clock;
  wire  line_1609_reset;
  wire  line_1609_valid;
  reg  line_1609_valid_reg;
  wire  line_1610_clock;
  wire  line_1610_reset;
  wire  line_1610_valid;
  reg  line_1610_valid_reg;
  wire  line_1611_clock;
  wire  line_1611_reset;
  wire  line_1611_valid;
  reg  line_1611_valid_reg;
  wire  line_1612_clock;
  wire  line_1612_reset;
  wire  line_1612_valid;
  reg  line_1612_valid_reg;
  wire  line_1613_clock;
  wire  line_1613_reset;
  wire  line_1613_valid;
  reg  line_1613_valid_reg;
  wire  line_1614_clock;
  wire  line_1614_reset;
  wire  line_1614_valid;
  reg  line_1614_valid_reg;
  wire  line_1615_clock;
  wire  line_1615_reset;
  wire  line_1615_valid;
  reg  line_1615_valid_reg;
  wire  line_1616_clock;
  wire  line_1616_reset;
  wire  line_1616_valid;
  reg  line_1616_valid_reg;
  wire  line_1617_clock;
  wire  line_1617_reset;
  wire  line_1617_valid;
  reg  line_1617_valid_reg;
  wire  line_1618_clock;
  wire  line_1618_reset;
  wire  line_1618_valid;
  reg  line_1618_valid_reg;
  wire  line_1619_clock;
  wire  line_1619_reset;
  wire  line_1619_valid;
  reg  line_1619_valid_reg;
  wire  line_1620_clock;
  wire  line_1620_reset;
  wire  line_1620_valid;
  reg  line_1620_valid_reg;
  wire  line_1621_clock;
  wire  line_1621_reset;
  wire  line_1621_valid;
  reg  line_1621_valid_reg;
  wire  line_1622_clock;
  wire  line_1622_reset;
  wire  line_1622_valid;
  reg  line_1622_valid_reg;
  wire  line_1623_clock;
  wire  line_1623_reset;
  wire  line_1623_valid;
  reg  line_1623_valid_reg;
  wire  line_1624_clock;
  wire  line_1624_reset;
  wire  line_1624_valid;
  reg  line_1624_valid_reg;
  wire  line_1625_clock;
  wire  line_1625_reset;
  wire  line_1625_valid;
  reg  line_1625_valid_reg;
  wire  _dequeueSize_T = backend_io_in_0_ready & backend_io_in_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] dequeueSize = {{1'd0}, _dequeueSize_T}; // @[src/main/scala/utils/PipelineVector.scala 64:42]
  wire  dequeueFire = dequeueSize > 2'h0; // @[src/main/scala/utils/PipelineVector.scala 65:35]
  wire  line_1626_clock;
  wire  line_1626_reset;
  wire  line_1626_valid;
  reg  line_1626_valid_reg;
  wire [1:0] _ringBufferTail_T_1 = ringBufferTail + dequeueSize; // @[src/main/scala/utils/PipelineVector.scala 67:42]
  wire  line_1627_clock;
  wire  line_1627_reset;
  wire  line_1627_valid;
  reg  line_1627_valid_reg;
  Frontend_inorder frontend ( // @[src/main/scala/nutcore/NutCore.scala 131:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(frontend_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(frontend_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_iaf(frontend_io_iaf),
    .io_sfence_vma_invalid(frontend_io_sfence_vma_invalid),
    .io_wfi_invalid(frontend_io_wfi_invalid),
    .REG_valid(frontend_REG_valid),
    .REG_pc(frontend_REG_pc),
    .REG_isMissPredict(frontend_REG_isMissPredict),
    .REG_actualTarget(frontend_REG_actualTarget),
    .REG_actualTaken(frontend_REG_actualTaken),
    .REG_fuOpType(frontend_REG_fuOpType),
    .REG_btbType(frontend_REG_btbType),
    .REG_isRVC(frontend_REG_isRVC),
    .isWFI(frontend_isWFI),
    .flushICache(frontend_flushICache),
    .flushTLB(frontend_flushTLB),
    .intrVecIDU(frontend_intrVecIDU)
  );
  Backend_inorder backend ( // @[src/main/scala/nutcore/NutCore.scala 174:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(backend_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(backend_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(backend_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(backend_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(backend_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(backend_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(backend_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(backend_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(backend_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_laf(backend_io_memMMU_dmem_laf),
    .io_memMMU_dmem_saf(backend_io_memMMU_dmem_saf),
    .io_sfence_vma_invalid(backend_io_sfence_vma_invalid),
    .io_wfi_invalid(backend_io_wfi_invalid),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    .lr(backend_lr),
    .io_extra_meip_0(backend_io_extra_meip_0),
    .scInflight(backend_scInflight),
    .REG_valid(backend_REG_valid),
    .REG_pc(backend_REG_pc),
    .REG_isMissPredict(backend_REG_isMissPredict),
    .REG_actualTarget(backend_REG_actualTarget),
    .REG_actualTaken(backend_REG_actualTaken),
    .REG_fuOpType(backend_REG_fuOpType),
    .REG_btbType(backend_REG_btbType),
    .REG_isRVC(backend_REG_isRVC),
    .amoReq(backend_amoReq),
    .lrAddr(backend_lrAddr),
    .paddr(backend_paddr),
    .satp(backend_satp),
    ._T_12(backend__T_12),
    .scIsSuccess(backend_scIsSuccess),
    .io_extra_mtip(backend_io_extra_mtip),
    .flushICache(backend_flushICache),
    .vmEnable(backend_vmEnable),
    .flushTLB(backend_flushTLB),
    .intrVecIDU(backend_intrVecIDU),
    .tlbFinish(backend_tlbFinish),
    .ismmio(backend_ismmio),
    ._T_13_0(backend__T_13_0),
    .io_extra_msip(backend_io_extra_msip)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[src/main/scala/nutcore/NutCore.scala 178:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[src/main/scala/nutcore/NutCore.scala 179:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(dmemXbar_io_in_1_req_ready),
    .io_in_1_req_valid(dmemXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(dmemXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(dmemXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(dmemXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(dmemXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(dmemXbar_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(dmemXbar_io_in_2_req_ready),
    .io_in_2_req_valid(dmemXbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(dmemXbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(dmemXbar_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(dmemXbar_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(dmemXbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(dmemXbar_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(dmemXbar_io_in_3_req_ready),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  EmbeddedTLB itlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user),
    .io_mem_req_ready(itlb_io_mem_req_ready),
    .io_mem_req_valid(itlb_io_mem_req_valid),
    .io_mem_req_bits_addr(itlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(itlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(itlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(itlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(itlb_io_mem_resp_bits_rdata),
    .io_flush(itlb_io_flush),
    .io_csrMMU_priviledgeMode(itlb_io_csrMMU_priviledgeMode),
    .io_iaf(itlb_io_iaf),
    .CSRSATP(itlb_CSRSATP),
    .MOUFlushTLB(itlb_MOUFlushTLB)
  );
  PTERequestFilter filter ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_in_req_ready(filter_io_in_req_ready),
    .io_in_req_valid(filter_io_in_req_valid),
    .io_in_req_bits_addr(filter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_io_out_req_ready),
    .io_out_req_valid(filter_io_out_req_valid),
    .io_out_req_bits_addr(filter_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_io_out_resp_bits_rdata),
    .io_u(filter_io_u)
  );
  Cache_fake io_imem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_imem_cache_clock),
    .reset(io_imem_cache_reset),
    .io_in_req_ready(io_imem_cache_io_in_req_ready),
    .io_in_req_valid(io_imem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_imem_cache_io_in_req_bits_addr),
    .io_in_req_bits_user(io_imem_cache_io_in_req_bits_user),
    .io_in_resp_ready(io_imem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_imem_cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(io_imem_cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(io_imem_cache_io_in_resp_bits_user),
    .io_flush(io_imem_cache_io_flush),
    .io_out_mem_req_ready(io_imem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_imem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_imem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(io_imem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_imem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_rdata(io_imem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_imem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_imem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_imem_cache_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(io_imem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_imem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_imem_cache_io_mmio_resp_bits_rdata)
  );
  EmbeddedTLB_1 dtlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(dtlb_clock),
    .reset(dtlb_reset),
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata),
    .io_mem_req_ready(dtlb_io_mem_req_ready),
    .io_mem_req_valid(dtlb_io_mem_req_valid),
    .io_mem_req_bits_addr(dtlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(dtlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(dtlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(dtlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(dtlb_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(dtlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(dtlb_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(dtlb_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(dtlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(dtlb_io_csrMMU_storePF),
    .io_csrMMU_laf(dtlb_io_csrMMU_laf),
    .io_csrMMU_saf(dtlb_io_csrMMU_saf),
    .lr(dtlb_lr),
    .scInflight(dtlb_scInflight),
    .amoReq(dtlb_amoReq),
    .lrAddr(dtlb_lrAddr),
    .paddr(dtlb_paddr),
    .CSRSATP(dtlb_CSRSATP),
    ._T_12_0(dtlb__T_12_0),
    .scIsSuccess_0(dtlb_scIsSuccess_0),
    .vmEnable_0(dtlb_vmEnable_0),
    .MOUFlushTLB(dtlb_MOUFlushTLB),
    .tlbFinish_0(dtlb_tlbFinish_0),
    ._T_13_1(dtlb__T_13_1)
  );
  PTERequestFilter_1 filter_1 ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_1_clock),
    .reset(filter_1_reset),
    .io_in_req_ready(filter_1_io_in_req_ready),
    .io_in_req_valid(filter_1_io_in_req_valid),
    .io_in_req_bits_addr(filter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_1_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_1_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_1_io_out_req_ready),
    .io_out_req_valid(filter_1_io_out_req_valid),
    .io_out_req_bits_addr(filter_1_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_1_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_1_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_1_io_out_resp_bits_rdata),
    .io_u(filter_1_io_u)
  );
  Cache_fake_1 io_dmem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_dmem_cache_clock),
    .reset(io_dmem_cache_reset),
    .io_in_req_ready(io_dmem_cache_io_in_req_ready),
    .io_in_req_valid(io_dmem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_dmem_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(io_dmem_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_dmem_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_dmem_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_dmem_cache_io_in_req_bits_wdata),
    .io_in_resp_valid(io_dmem_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_dmem_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_dmem_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(io_dmem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_dmem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_dmem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_size(io_dmem_cache_io_out_mem_req_bits_size),
    .io_out_mem_req_bits_cmd(io_dmem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wmask(io_dmem_cache_io_out_mem_req_bits_wmask),
    .io_out_mem_req_bits_wdata(io_dmem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(io_dmem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_dmem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_dmem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_dmem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_dmem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_dmem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_dmem_cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(io_dmem_cache_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(io_dmem_cache_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(io_dmem_cache_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(io_dmem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_dmem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(io_dmem_cache_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(io_dmem_cache_io_mmio_resp_bits_rdata),
    .ismmio_0(io_dmem_cache_ismmio_0)
  );
  GEN_w1_line #(.COVER_INDEX(727)) line_727 (
    .clock(line_727_clock),
    .reset(line_727_reset),
    .valid(line_727_valid)
  );
  GEN_w1_line #(.COVER_INDEX(728)) line_728 (
    .clock(line_728_clock),
    .reset(line_728_reset),
    .valid(line_728_valid)
  );
  GEN_w1_line #(.COVER_INDEX(729)) line_729 (
    .clock(line_729_clock),
    .reset(line_729_reset),
    .valid(line_729_valid)
  );
  GEN_w1_line #(.COVER_INDEX(730)) line_730 (
    .clock(line_730_clock),
    .reset(line_730_reset),
    .valid(line_730_valid)
  );
  GEN_w1_line #(.COVER_INDEX(731)) line_731 (
    .clock(line_731_clock),
    .reset(line_731_reset),
    .valid(line_731_valid)
  );
  GEN_w1_line #(.COVER_INDEX(732)) line_732 (
    .clock(line_732_clock),
    .reset(line_732_reset),
    .valid(line_732_valid)
  );
  GEN_w1_line #(.COVER_INDEX(733)) line_733 (
    .clock(line_733_clock),
    .reset(line_733_reset),
    .valid(line_733_valid)
  );
  GEN_w1_line #(.COVER_INDEX(734)) line_734 (
    .clock(line_734_clock),
    .reset(line_734_reset),
    .valid(line_734_valid)
  );
  GEN_w1_line #(.COVER_INDEX(735)) line_735 (
    .clock(line_735_clock),
    .reset(line_735_reset),
    .valid(line_735_valid)
  );
  GEN_w1_line #(.COVER_INDEX(736)) line_736 (
    .clock(line_736_clock),
    .reset(line_736_reset),
    .valid(line_736_valid)
  );
  GEN_w1_line #(.COVER_INDEX(737)) line_737 (
    .clock(line_737_clock),
    .reset(line_737_reset),
    .valid(line_737_valid)
  );
  GEN_w1_line #(.COVER_INDEX(738)) line_738 (
    .clock(line_738_clock),
    .reset(line_738_reset),
    .valid(line_738_valid)
  );
  GEN_w1_line #(.COVER_INDEX(739)) line_739 (
    .clock(line_739_clock),
    .reset(line_739_reset),
    .valid(line_739_valid)
  );
  GEN_w1_line #(.COVER_INDEX(740)) line_740 (
    .clock(line_740_clock),
    .reset(line_740_reset),
    .valid(line_740_valid)
  );
  GEN_w1_line #(.COVER_INDEX(741)) line_741 (
    .clock(line_741_clock),
    .reset(line_741_reset),
    .valid(line_741_valid)
  );
  GEN_w1_line #(.COVER_INDEX(742)) line_742 (
    .clock(line_742_clock),
    .reset(line_742_reset),
    .valid(line_742_valid)
  );
  GEN_w1_line #(.COVER_INDEX(743)) line_743 (
    .clock(line_743_clock),
    .reset(line_743_reset),
    .valid(line_743_valid)
  );
  GEN_w1_line #(.COVER_INDEX(744)) line_744 (
    .clock(line_744_clock),
    .reset(line_744_reset),
    .valid(line_744_valid)
  );
  GEN_w1_line #(.COVER_INDEX(745)) line_745 (
    .clock(line_745_clock),
    .reset(line_745_reset),
    .valid(line_745_valid)
  );
  GEN_w1_line #(.COVER_INDEX(746)) line_746 (
    .clock(line_746_clock),
    .reset(line_746_reset),
    .valid(line_746_valid)
  );
  GEN_w1_line #(.COVER_INDEX(747)) line_747 (
    .clock(line_747_clock),
    .reset(line_747_reset),
    .valid(line_747_valid)
  );
  GEN_w1_line #(.COVER_INDEX(748)) line_748 (
    .clock(line_748_clock),
    .reset(line_748_reset),
    .valid(line_748_valid)
  );
  GEN_w1_line #(.COVER_INDEX(749)) line_749 (
    .clock(line_749_clock),
    .reset(line_749_reset),
    .valid(line_749_valid)
  );
  GEN_w1_line #(.COVER_INDEX(750)) line_750 (
    .clock(line_750_clock),
    .reset(line_750_reset),
    .valid(line_750_valid)
  );
  GEN_w1_line #(.COVER_INDEX(751)) line_751 (
    .clock(line_751_clock),
    .reset(line_751_reset),
    .valid(line_751_valid)
  );
  GEN_w1_line #(.COVER_INDEX(752)) line_752 (
    .clock(line_752_clock),
    .reset(line_752_reset),
    .valid(line_752_valid)
  );
  GEN_w1_line #(.COVER_INDEX(753)) line_753 (
    .clock(line_753_clock),
    .reset(line_753_reset),
    .valid(line_753_valid)
  );
  GEN_w1_line #(.COVER_INDEX(754)) line_754 (
    .clock(line_754_clock),
    .reset(line_754_reset),
    .valid(line_754_valid)
  );
  GEN_w1_line #(.COVER_INDEX(755)) line_755 (
    .clock(line_755_clock),
    .reset(line_755_reset),
    .valid(line_755_valid)
  );
  GEN_w1_line #(.COVER_INDEX(756)) line_756 (
    .clock(line_756_clock),
    .reset(line_756_reset),
    .valid(line_756_valid)
  );
  GEN_w1_line #(.COVER_INDEX(757)) line_757 (
    .clock(line_757_clock),
    .reset(line_757_reset),
    .valid(line_757_valid)
  );
  GEN_w1_line #(.COVER_INDEX(758)) line_758 (
    .clock(line_758_clock),
    .reset(line_758_reset),
    .valid(line_758_valid)
  );
  GEN_w1_line #(.COVER_INDEX(759)) line_759 (
    .clock(line_759_clock),
    .reset(line_759_reset),
    .valid(line_759_valid)
  );
  GEN_w1_line #(.COVER_INDEX(760)) line_760 (
    .clock(line_760_clock),
    .reset(line_760_reset),
    .valid(line_760_valid)
  );
  GEN_w1_line #(.COVER_INDEX(761)) line_761 (
    .clock(line_761_clock),
    .reset(line_761_reset),
    .valid(line_761_valid)
  );
  GEN_w1_line #(.COVER_INDEX(762)) line_762 (
    .clock(line_762_clock),
    .reset(line_762_reset),
    .valid(line_762_valid)
  );
  GEN_w1_line #(.COVER_INDEX(763)) line_763 (
    .clock(line_763_clock),
    .reset(line_763_reset),
    .valid(line_763_valid)
  );
  GEN_w1_line #(.COVER_INDEX(764)) line_764 (
    .clock(line_764_clock),
    .reset(line_764_reset),
    .valid(line_764_valid)
  );
  GEN_w1_line #(.COVER_INDEX(765)) line_765 (
    .clock(line_765_clock),
    .reset(line_765_reset),
    .valid(line_765_valid)
  );
  GEN_w1_line #(.COVER_INDEX(766)) line_766 (
    .clock(line_766_clock),
    .reset(line_766_reset),
    .valid(line_766_valid)
  );
  GEN_w1_line #(.COVER_INDEX(767)) line_767 (
    .clock(line_767_clock),
    .reset(line_767_reset),
    .valid(line_767_valid)
  );
  GEN_w1_line #(.COVER_INDEX(768)) line_768 (
    .clock(line_768_clock),
    .reset(line_768_reset),
    .valid(line_768_valid)
  );
  GEN_w1_line #(.COVER_INDEX(769)) line_769 (
    .clock(line_769_clock),
    .reset(line_769_reset),
    .valid(line_769_valid)
  );
  GEN_w1_line #(.COVER_INDEX(770)) line_770 (
    .clock(line_770_clock),
    .reset(line_770_reset),
    .valid(line_770_valid)
  );
  GEN_w1_line #(.COVER_INDEX(771)) line_771 (
    .clock(line_771_clock),
    .reset(line_771_reset),
    .valid(line_771_valid)
  );
  GEN_w1_line #(.COVER_INDEX(772)) line_772 (
    .clock(line_772_clock),
    .reset(line_772_reset),
    .valid(line_772_valid)
  );
  GEN_w1_line #(.COVER_INDEX(773)) line_773 (
    .clock(line_773_clock),
    .reset(line_773_reset),
    .valid(line_773_valid)
  );
  GEN_w1_line #(.COVER_INDEX(774)) line_774 (
    .clock(line_774_clock),
    .reset(line_774_reset),
    .valid(line_774_valid)
  );
  GEN_w1_line #(.COVER_INDEX(775)) line_775 (
    .clock(line_775_clock),
    .reset(line_775_reset),
    .valid(line_775_valid)
  );
  GEN_w1_line #(.COVER_INDEX(776)) line_776 (
    .clock(line_776_clock),
    .reset(line_776_reset),
    .valid(line_776_valid)
  );
  GEN_w1_line #(.COVER_INDEX(777)) line_777 (
    .clock(line_777_clock),
    .reset(line_777_reset),
    .valid(line_777_valid)
  );
  GEN_w1_line #(.COVER_INDEX(778)) line_778 (
    .clock(line_778_clock),
    .reset(line_778_reset),
    .valid(line_778_valid)
  );
  GEN_w1_line #(.COVER_INDEX(779)) line_779 (
    .clock(line_779_clock),
    .reset(line_779_reset),
    .valid(line_779_valid)
  );
  GEN_w1_line #(.COVER_INDEX(780)) line_780 (
    .clock(line_780_clock),
    .reset(line_780_reset),
    .valid(line_780_valid)
  );
  GEN_w1_line #(.COVER_INDEX(781)) line_781 (
    .clock(line_781_clock),
    .reset(line_781_reset),
    .valid(line_781_valid)
  );
  GEN_w1_line #(.COVER_INDEX(782)) line_782 (
    .clock(line_782_clock),
    .reset(line_782_reset),
    .valid(line_782_valid)
  );
  GEN_w1_line #(.COVER_INDEX(783)) line_783 (
    .clock(line_783_clock),
    .reset(line_783_reset),
    .valid(line_783_valid)
  );
  GEN_w1_line #(.COVER_INDEX(784)) line_784 (
    .clock(line_784_clock),
    .reset(line_784_reset),
    .valid(line_784_valid)
  );
  GEN_w1_line #(.COVER_INDEX(785)) line_785 (
    .clock(line_785_clock),
    .reset(line_785_reset),
    .valid(line_785_valid)
  );
  GEN_w1_line #(.COVER_INDEX(786)) line_786 (
    .clock(line_786_clock),
    .reset(line_786_reset),
    .valid(line_786_valid)
  );
  GEN_w1_line #(.COVER_INDEX(787)) line_787 (
    .clock(line_787_clock),
    .reset(line_787_reset),
    .valid(line_787_valid)
  );
  GEN_w1_line #(.COVER_INDEX(788)) line_788 (
    .clock(line_788_clock),
    .reset(line_788_reset),
    .valid(line_788_valid)
  );
  GEN_w1_line #(.COVER_INDEX(789)) line_789 (
    .clock(line_789_clock),
    .reset(line_789_reset),
    .valid(line_789_valid)
  );
  GEN_w1_line #(.COVER_INDEX(790)) line_790 (
    .clock(line_790_clock),
    .reset(line_790_reset),
    .valid(line_790_valid)
  );
  GEN_w1_line #(.COVER_INDEX(791)) line_791 (
    .clock(line_791_clock),
    .reset(line_791_reset),
    .valid(line_791_valid)
  );
  GEN_w1_line #(.COVER_INDEX(792)) line_792 (
    .clock(line_792_clock),
    .reset(line_792_reset),
    .valid(line_792_valid)
  );
  GEN_w1_line #(.COVER_INDEX(793)) line_793 (
    .clock(line_793_clock),
    .reset(line_793_reset),
    .valid(line_793_valid)
  );
  GEN_w1_line #(.COVER_INDEX(794)) line_794 (
    .clock(line_794_clock),
    .reset(line_794_reset),
    .valid(line_794_valid)
  );
  GEN_w1_line #(.COVER_INDEX(795)) line_795 (
    .clock(line_795_clock),
    .reset(line_795_reset),
    .valid(line_795_valid)
  );
  GEN_w1_line #(.COVER_INDEX(796)) line_796 (
    .clock(line_796_clock),
    .reset(line_796_reset),
    .valid(line_796_valid)
  );
  GEN_w1_line #(.COVER_INDEX(797)) line_797 (
    .clock(line_797_clock),
    .reset(line_797_reset),
    .valid(line_797_valid)
  );
  GEN_w1_line #(.COVER_INDEX(798)) line_798 (
    .clock(line_798_clock),
    .reset(line_798_reset),
    .valid(line_798_valid)
  );
  GEN_w1_line #(.COVER_INDEX(799)) line_799 (
    .clock(line_799_clock),
    .reset(line_799_reset),
    .valid(line_799_valid)
  );
  GEN_w1_line #(.COVER_INDEX(800)) line_800 (
    .clock(line_800_clock),
    .reset(line_800_reset),
    .valid(line_800_valid)
  );
  GEN_w1_line #(.COVER_INDEX(801)) line_801 (
    .clock(line_801_clock),
    .reset(line_801_reset),
    .valid(line_801_valid)
  );
  GEN_w1_line #(.COVER_INDEX(802)) line_802 (
    .clock(line_802_clock),
    .reset(line_802_reset),
    .valid(line_802_valid)
  );
  GEN_w1_line #(.COVER_INDEX(803)) line_803 (
    .clock(line_803_clock),
    .reset(line_803_reset),
    .valid(line_803_valid)
  );
  GEN_w1_line #(.COVER_INDEX(804)) line_804 (
    .clock(line_804_clock),
    .reset(line_804_reset),
    .valid(line_804_valid)
  );
  GEN_w1_line #(.COVER_INDEX(805)) line_805 (
    .clock(line_805_clock),
    .reset(line_805_reset),
    .valid(line_805_valid)
  );
  GEN_w1_line #(.COVER_INDEX(806)) line_806 (
    .clock(line_806_clock),
    .reset(line_806_reset),
    .valid(line_806_valid)
  );
  GEN_w1_line #(.COVER_INDEX(807)) line_807 (
    .clock(line_807_clock),
    .reset(line_807_reset),
    .valid(line_807_valid)
  );
  GEN_w1_line #(.COVER_INDEX(808)) line_808 (
    .clock(line_808_clock),
    .reset(line_808_reset),
    .valid(line_808_valid)
  );
  GEN_w1_line #(.COVER_INDEX(809)) line_809 (
    .clock(line_809_clock),
    .reset(line_809_reset),
    .valid(line_809_valid)
  );
  GEN_w1_line #(.COVER_INDEX(810)) line_810 (
    .clock(line_810_clock),
    .reset(line_810_reset),
    .valid(line_810_valid)
  );
  GEN_w1_line #(.COVER_INDEX(811)) line_811 (
    .clock(line_811_clock),
    .reset(line_811_reset),
    .valid(line_811_valid)
  );
  GEN_w1_line #(.COVER_INDEX(812)) line_812 (
    .clock(line_812_clock),
    .reset(line_812_reset),
    .valid(line_812_valid)
  );
  GEN_w1_line #(.COVER_INDEX(813)) line_813 (
    .clock(line_813_clock),
    .reset(line_813_reset),
    .valid(line_813_valid)
  );
  GEN_w1_line #(.COVER_INDEX(814)) line_814 (
    .clock(line_814_clock),
    .reset(line_814_reset),
    .valid(line_814_valid)
  );
  GEN_w1_line #(.COVER_INDEX(815)) line_815 (
    .clock(line_815_clock),
    .reset(line_815_reset),
    .valid(line_815_valid)
  );
  GEN_w1_line #(.COVER_INDEX(816)) line_816 (
    .clock(line_816_clock),
    .reset(line_816_reset),
    .valid(line_816_valid)
  );
  GEN_w1_line #(.COVER_INDEX(817)) line_817 (
    .clock(line_817_clock),
    .reset(line_817_reset),
    .valid(line_817_valid)
  );
  GEN_w1_line #(.COVER_INDEX(818)) line_818 (
    .clock(line_818_clock),
    .reset(line_818_reset),
    .valid(line_818_valid)
  );
  GEN_w1_line #(.COVER_INDEX(819)) line_819 (
    .clock(line_819_clock),
    .reset(line_819_reset),
    .valid(line_819_valid)
  );
  GEN_w1_line #(.COVER_INDEX(820)) line_820 (
    .clock(line_820_clock),
    .reset(line_820_reset),
    .valid(line_820_valid)
  );
  GEN_w1_line #(.COVER_INDEX(821)) line_821 (
    .clock(line_821_clock),
    .reset(line_821_reset),
    .valid(line_821_valid)
  );
  GEN_w1_line #(.COVER_INDEX(822)) line_822 (
    .clock(line_822_clock),
    .reset(line_822_reset),
    .valid(line_822_valid)
  );
  GEN_w1_line #(.COVER_INDEX(823)) line_823 (
    .clock(line_823_clock),
    .reset(line_823_reset),
    .valid(line_823_valid)
  );
  GEN_w1_line #(.COVER_INDEX(824)) line_824 (
    .clock(line_824_clock),
    .reset(line_824_reset),
    .valid(line_824_valid)
  );
  GEN_w1_line #(.COVER_INDEX(825)) line_825 (
    .clock(line_825_clock),
    .reset(line_825_reset),
    .valid(line_825_valid)
  );
  GEN_w1_line #(.COVER_INDEX(826)) line_826 (
    .clock(line_826_clock),
    .reset(line_826_reset),
    .valid(line_826_valid)
  );
  GEN_w1_line #(.COVER_INDEX(827)) line_827 (
    .clock(line_827_clock),
    .reset(line_827_reset),
    .valid(line_827_valid)
  );
  GEN_w1_line #(.COVER_INDEX(828)) line_828 (
    .clock(line_828_clock),
    .reset(line_828_reset),
    .valid(line_828_valid)
  );
  GEN_w1_line #(.COVER_INDEX(829)) line_829 (
    .clock(line_829_clock),
    .reset(line_829_reset),
    .valid(line_829_valid)
  );
  GEN_w1_line #(.COVER_INDEX(830)) line_830 (
    .clock(line_830_clock),
    .reset(line_830_reset),
    .valid(line_830_valid)
  );
  GEN_w1_line #(.COVER_INDEX(831)) line_831 (
    .clock(line_831_clock),
    .reset(line_831_reset),
    .valid(line_831_valid)
  );
  GEN_w1_line #(.COVER_INDEX(832)) line_832 (
    .clock(line_832_clock),
    .reset(line_832_reset),
    .valid(line_832_valid)
  );
  GEN_w1_line #(.COVER_INDEX(833)) line_833 (
    .clock(line_833_clock),
    .reset(line_833_reset),
    .valid(line_833_valid)
  );
  GEN_w1_line #(.COVER_INDEX(834)) line_834 (
    .clock(line_834_clock),
    .reset(line_834_reset),
    .valid(line_834_valid)
  );
  GEN_w1_line #(.COVER_INDEX(835)) line_835 (
    .clock(line_835_clock),
    .reset(line_835_reset),
    .valid(line_835_valid)
  );
  GEN_w1_line #(.COVER_INDEX(836)) line_836 (
    .clock(line_836_clock),
    .reset(line_836_reset),
    .valid(line_836_valid)
  );
  GEN_w1_line #(.COVER_INDEX(837)) line_837 (
    .clock(line_837_clock),
    .reset(line_837_reset),
    .valid(line_837_valid)
  );
  GEN_w1_line #(.COVER_INDEX(838)) line_838 (
    .clock(line_838_clock),
    .reset(line_838_reset),
    .valid(line_838_valid)
  );
  GEN_w1_line #(.COVER_INDEX(839)) line_839 (
    .clock(line_839_clock),
    .reset(line_839_reset),
    .valid(line_839_valid)
  );
  GEN_w1_line #(.COVER_INDEX(840)) line_840 (
    .clock(line_840_clock),
    .reset(line_840_reset),
    .valid(line_840_valid)
  );
  GEN_w1_line #(.COVER_INDEX(841)) line_841 (
    .clock(line_841_clock),
    .reset(line_841_reset),
    .valid(line_841_valid)
  );
  GEN_w1_line #(.COVER_INDEX(842)) line_842 (
    .clock(line_842_clock),
    .reset(line_842_reset),
    .valid(line_842_valid)
  );
  GEN_w1_line #(.COVER_INDEX(843)) line_843 (
    .clock(line_843_clock),
    .reset(line_843_reset),
    .valid(line_843_valid)
  );
  GEN_w1_line #(.COVER_INDEX(844)) line_844 (
    .clock(line_844_clock),
    .reset(line_844_reset),
    .valid(line_844_valid)
  );
  GEN_w1_line #(.COVER_INDEX(845)) line_845 (
    .clock(line_845_clock),
    .reset(line_845_reset),
    .valid(line_845_valid)
  );
  GEN_w1_line #(.COVER_INDEX(846)) line_846 (
    .clock(line_846_clock),
    .reset(line_846_reset),
    .valid(line_846_valid)
  );
  GEN_w1_line #(.COVER_INDEX(847)) line_847 (
    .clock(line_847_clock),
    .reset(line_847_reset),
    .valid(line_847_valid)
  );
  GEN_w1_line #(.COVER_INDEX(848)) line_848 (
    .clock(line_848_clock),
    .reset(line_848_reset),
    .valid(line_848_valid)
  );
  GEN_w1_line #(.COVER_INDEX(849)) line_849 (
    .clock(line_849_clock),
    .reset(line_849_reset),
    .valid(line_849_valid)
  );
  GEN_w1_line #(.COVER_INDEX(850)) line_850 (
    .clock(line_850_clock),
    .reset(line_850_reset),
    .valid(line_850_valid)
  );
  GEN_w1_line #(.COVER_INDEX(851)) line_851 (
    .clock(line_851_clock),
    .reset(line_851_reset),
    .valid(line_851_valid)
  );
  GEN_w1_line #(.COVER_INDEX(852)) line_852 (
    .clock(line_852_clock),
    .reset(line_852_reset),
    .valid(line_852_valid)
  );
  GEN_w1_line #(.COVER_INDEX(853)) line_853 (
    .clock(line_853_clock),
    .reset(line_853_reset),
    .valid(line_853_valid)
  );
  GEN_w1_line #(.COVER_INDEX(854)) line_854 (
    .clock(line_854_clock),
    .reset(line_854_reset),
    .valid(line_854_valid)
  );
  GEN_w1_line #(.COVER_INDEX(855)) line_855 (
    .clock(line_855_clock),
    .reset(line_855_reset),
    .valid(line_855_valid)
  );
  GEN_w1_line #(.COVER_INDEX(856)) line_856 (
    .clock(line_856_clock),
    .reset(line_856_reset),
    .valid(line_856_valid)
  );
  GEN_w1_line #(.COVER_INDEX(857)) line_857 (
    .clock(line_857_clock),
    .reset(line_857_reset),
    .valid(line_857_valid)
  );
  GEN_w1_line #(.COVER_INDEX(858)) line_858 (
    .clock(line_858_clock),
    .reset(line_858_reset),
    .valid(line_858_valid)
  );
  GEN_w1_line #(.COVER_INDEX(859)) line_859 (
    .clock(line_859_clock),
    .reset(line_859_reset),
    .valid(line_859_valid)
  );
  GEN_w1_line #(.COVER_INDEX(860)) line_860 (
    .clock(line_860_clock),
    .reset(line_860_reset),
    .valid(line_860_valid)
  );
  GEN_w1_line #(.COVER_INDEX(861)) line_861 (
    .clock(line_861_clock),
    .reset(line_861_reset),
    .valid(line_861_valid)
  );
  GEN_w1_line #(.COVER_INDEX(862)) line_862 (
    .clock(line_862_clock),
    .reset(line_862_reset),
    .valid(line_862_valid)
  );
  GEN_w1_line #(.COVER_INDEX(863)) line_863 (
    .clock(line_863_clock),
    .reset(line_863_reset),
    .valid(line_863_valid)
  );
  GEN_w1_line #(.COVER_INDEX(864)) line_864 (
    .clock(line_864_clock),
    .reset(line_864_reset),
    .valid(line_864_valid)
  );
  GEN_w1_line #(.COVER_INDEX(865)) line_865 (
    .clock(line_865_clock),
    .reset(line_865_reset),
    .valid(line_865_valid)
  );
  GEN_w1_line #(.COVER_INDEX(866)) line_866 (
    .clock(line_866_clock),
    .reset(line_866_reset),
    .valid(line_866_valid)
  );
  GEN_w1_line #(.COVER_INDEX(867)) line_867 (
    .clock(line_867_clock),
    .reset(line_867_reset),
    .valid(line_867_valid)
  );
  GEN_w1_line #(.COVER_INDEX(868)) line_868 (
    .clock(line_868_clock),
    .reset(line_868_reset),
    .valid(line_868_valid)
  );
  GEN_w1_line #(.COVER_INDEX(869)) line_869 (
    .clock(line_869_clock),
    .reset(line_869_reset),
    .valid(line_869_valid)
  );
  GEN_w1_line #(.COVER_INDEX(870)) line_870 (
    .clock(line_870_clock),
    .reset(line_870_reset),
    .valid(line_870_valid)
  );
  GEN_w1_line #(.COVER_INDEX(871)) line_871 (
    .clock(line_871_clock),
    .reset(line_871_reset),
    .valid(line_871_valid)
  );
  GEN_w1_line #(.COVER_INDEX(872)) line_872 (
    .clock(line_872_clock),
    .reset(line_872_reset),
    .valid(line_872_valid)
  );
  GEN_w1_line #(.COVER_INDEX(873)) line_873 (
    .clock(line_873_clock),
    .reset(line_873_reset),
    .valid(line_873_valid)
  );
  GEN_w1_line #(.COVER_INDEX(874)) line_874 (
    .clock(line_874_clock),
    .reset(line_874_reset),
    .valid(line_874_valid)
  );
  GEN_w1_line #(.COVER_INDEX(875)) line_875 (
    .clock(line_875_clock),
    .reset(line_875_reset),
    .valid(line_875_valid)
  );
  GEN_w1_line #(.COVER_INDEX(876)) line_876 (
    .clock(line_876_clock),
    .reset(line_876_reset),
    .valid(line_876_valid)
  );
  GEN_w1_line #(.COVER_INDEX(877)) line_877 (
    .clock(line_877_clock),
    .reset(line_877_reset),
    .valid(line_877_valid)
  );
  GEN_w1_line #(.COVER_INDEX(878)) line_878 (
    .clock(line_878_clock),
    .reset(line_878_reset),
    .valid(line_878_valid)
  );
  GEN_w1_line #(.COVER_INDEX(879)) line_879 (
    .clock(line_879_clock),
    .reset(line_879_reset),
    .valid(line_879_valid)
  );
  GEN_w1_line #(.COVER_INDEX(880)) line_880 (
    .clock(line_880_clock),
    .reset(line_880_reset),
    .valid(line_880_valid)
  );
  GEN_w1_line #(.COVER_INDEX(881)) line_881 (
    .clock(line_881_clock),
    .reset(line_881_reset),
    .valid(line_881_valid)
  );
  GEN_w1_line #(.COVER_INDEX(882)) line_882 (
    .clock(line_882_clock),
    .reset(line_882_reset),
    .valid(line_882_valid)
  );
  GEN_w1_line #(.COVER_INDEX(883)) line_883 (
    .clock(line_883_clock),
    .reset(line_883_reset),
    .valid(line_883_valid)
  );
  GEN_w1_line #(.COVER_INDEX(884)) line_884 (
    .clock(line_884_clock),
    .reset(line_884_reset),
    .valid(line_884_valid)
  );
  GEN_w1_line #(.COVER_INDEX(885)) line_885 (
    .clock(line_885_clock),
    .reset(line_885_reset),
    .valid(line_885_valid)
  );
  GEN_w1_line #(.COVER_INDEX(886)) line_886 (
    .clock(line_886_clock),
    .reset(line_886_reset),
    .valid(line_886_valid)
  );
  GEN_w1_line #(.COVER_INDEX(887)) line_887 (
    .clock(line_887_clock),
    .reset(line_887_reset),
    .valid(line_887_valid)
  );
  GEN_w1_line #(.COVER_INDEX(888)) line_888 (
    .clock(line_888_clock),
    .reset(line_888_reset),
    .valid(line_888_valid)
  );
  GEN_w1_line #(.COVER_INDEX(889)) line_889 (
    .clock(line_889_clock),
    .reset(line_889_reset),
    .valid(line_889_valid)
  );
  GEN_w1_line #(.COVER_INDEX(890)) line_890 (
    .clock(line_890_clock),
    .reset(line_890_reset),
    .valid(line_890_valid)
  );
  GEN_w1_line #(.COVER_INDEX(891)) line_891 (
    .clock(line_891_clock),
    .reset(line_891_reset),
    .valid(line_891_valid)
  );
  GEN_w1_line #(.COVER_INDEX(892)) line_892 (
    .clock(line_892_clock),
    .reset(line_892_reset),
    .valid(line_892_valid)
  );
  GEN_w1_line #(.COVER_INDEX(893)) line_893 (
    .clock(line_893_clock),
    .reset(line_893_reset),
    .valid(line_893_valid)
  );
  GEN_w1_line #(.COVER_INDEX(894)) line_894 (
    .clock(line_894_clock),
    .reset(line_894_reset),
    .valid(line_894_valid)
  );
  GEN_w1_line #(.COVER_INDEX(895)) line_895 (
    .clock(line_895_clock),
    .reset(line_895_reset),
    .valid(line_895_valid)
  );
  GEN_w1_line #(.COVER_INDEX(896)) line_896 (
    .clock(line_896_clock),
    .reset(line_896_reset),
    .valid(line_896_valid)
  );
  GEN_w1_line #(.COVER_INDEX(897)) line_897 (
    .clock(line_897_clock),
    .reset(line_897_reset),
    .valid(line_897_valid)
  );
  GEN_w1_line #(.COVER_INDEX(898)) line_898 (
    .clock(line_898_clock),
    .reset(line_898_reset),
    .valid(line_898_valid)
  );
  GEN_w1_line #(.COVER_INDEX(899)) line_899 (
    .clock(line_899_clock),
    .reset(line_899_reset),
    .valid(line_899_valid)
  );
  GEN_w1_line #(.COVER_INDEX(900)) line_900 (
    .clock(line_900_clock),
    .reset(line_900_reset),
    .valid(line_900_valid)
  );
  GEN_w1_line #(.COVER_INDEX(901)) line_901 (
    .clock(line_901_clock),
    .reset(line_901_reset),
    .valid(line_901_valid)
  );
  GEN_w1_line #(.COVER_INDEX(902)) line_902 (
    .clock(line_902_clock),
    .reset(line_902_reset),
    .valid(line_902_valid)
  );
  GEN_w1_line #(.COVER_INDEX(903)) line_903 (
    .clock(line_903_clock),
    .reset(line_903_reset),
    .valid(line_903_valid)
  );
  GEN_w1_line #(.COVER_INDEX(904)) line_904 (
    .clock(line_904_clock),
    .reset(line_904_reset),
    .valid(line_904_valid)
  );
  GEN_w1_line #(.COVER_INDEX(905)) line_905 (
    .clock(line_905_clock),
    .reset(line_905_reset),
    .valid(line_905_valid)
  );
  GEN_w1_line #(.COVER_INDEX(906)) line_906 (
    .clock(line_906_clock),
    .reset(line_906_reset),
    .valid(line_906_valid)
  );
  GEN_w1_line #(.COVER_INDEX(907)) line_907 (
    .clock(line_907_clock),
    .reset(line_907_reset),
    .valid(line_907_valid)
  );
  GEN_w1_line #(.COVER_INDEX(908)) line_908 (
    .clock(line_908_clock),
    .reset(line_908_reset),
    .valid(line_908_valid)
  );
  GEN_w1_line #(.COVER_INDEX(909)) line_909 (
    .clock(line_909_clock),
    .reset(line_909_reset),
    .valid(line_909_valid)
  );
  GEN_w1_line #(.COVER_INDEX(910)) line_910 (
    .clock(line_910_clock),
    .reset(line_910_reset),
    .valid(line_910_valid)
  );
  GEN_w1_line #(.COVER_INDEX(911)) line_911 (
    .clock(line_911_clock),
    .reset(line_911_reset),
    .valid(line_911_valid)
  );
  GEN_w1_line #(.COVER_INDEX(912)) line_912 (
    .clock(line_912_clock),
    .reset(line_912_reset),
    .valid(line_912_valid)
  );
  GEN_w1_line #(.COVER_INDEX(913)) line_913 (
    .clock(line_913_clock),
    .reset(line_913_reset),
    .valid(line_913_valid)
  );
  GEN_w1_line #(.COVER_INDEX(914)) line_914 (
    .clock(line_914_clock),
    .reset(line_914_reset),
    .valid(line_914_valid)
  );
  GEN_w1_line #(.COVER_INDEX(915)) line_915 (
    .clock(line_915_clock),
    .reset(line_915_reset),
    .valid(line_915_valid)
  );
  GEN_w1_line #(.COVER_INDEX(916)) line_916 (
    .clock(line_916_clock),
    .reset(line_916_reset),
    .valid(line_916_valid)
  );
  GEN_w1_line #(.COVER_INDEX(917)) line_917 (
    .clock(line_917_clock),
    .reset(line_917_reset),
    .valid(line_917_valid)
  );
  GEN_w1_line #(.COVER_INDEX(918)) line_918 (
    .clock(line_918_clock),
    .reset(line_918_reset),
    .valid(line_918_valid)
  );
  GEN_w1_line #(.COVER_INDEX(919)) line_919 (
    .clock(line_919_clock),
    .reset(line_919_reset),
    .valid(line_919_valid)
  );
  GEN_w1_line #(.COVER_INDEX(920)) line_920 (
    .clock(line_920_clock),
    .reset(line_920_reset),
    .valid(line_920_valid)
  );
  GEN_w1_line #(.COVER_INDEX(921)) line_921 (
    .clock(line_921_clock),
    .reset(line_921_reset),
    .valid(line_921_valid)
  );
  GEN_w1_line #(.COVER_INDEX(922)) line_922 (
    .clock(line_922_clock),
    .reset(line_922_reset),
    .valid(line_922_valid)
  );
  GEN_w1_line #(.COVER_INDEX(923)) line_923 (
    .clock(line_923_clock),
    .reset(line_923_reset),
    .valid(line_923_valid)
  );
  GEN_w1_line #(.COVER_INDEX(924)) line_924 (
    .clock(line_924_clock),
    .reset(line_924_reset),
    .valid(line_924_valid)
  );
  GEN_w1_line #(.COVER_INDEX(925)) line_925 (
    .clock(line_925_clock),
    .reset(line_925_reset),
    .valid(line_925_valid)
  );
  GEN_w1_line #(.COVER_INDEX(926)) line_926 (
    .clock(line_926_clock),
    .reset(line_926_reset),
    .valid(line_926_valid)
  );
  GEN_w1_line #(.COVER_INDEX(927)) line_927 (
    .clock(line_927_clock),
    .reset(line_927_reset),
    .valid(line_927_valid)
  );
  GEN_w1_line #(.COVER_INDEX(928)) line_928 (
    .clock(line_928_clock),
    .reset(line_928_reset),
    .valid(line_928_valid)
  );
  GEN_w1_line #(.COVER_INDEX(929)) line_929 (
    .clock(line_929_clock),
    .reset(line_929_reset),
    .valid(line_929_valid)
  );
  GEN_w1_line #(.COVER_INDEX(930)) line_930 (
    .clock(line_930_clock),
    .reset(line_930_reset),
    .valid(line_930_valid)
  );
  GEN_w1_line #(.COVER_INDEX(931)) line_931 (
    .clock(line_931_clock),
    .reset(line_931_reset),
    .valid(line_931_valid)
  );
  GEN_w1_line #(.COVER_INDEX(932)) line_932 (
    .clock(line_932_clock),
    .reset(line_932_reset),
    .valid(line_932_valid)
  );
  GEN_w1_line #(.COVER_INDEX(933)) line_933 (
    .clock(line_933_clock),
    .reset(line_933_reset),
    .valid(line_933_valid)
  );
  GEN_w1_line #(.COVER_INDEX(934)) line_934 (
    .clock(line_934_clock),
    .reset(line_934_reset),
    .valid(line_934_valid)
  );
  GEN_w1_line #(.COVER_INDEX(935)) line_935 (
    .clock(line_935_clock),
    .reset(line_935_reset),
    .valid(line_935_valid)
  );
  GEN_w1_line #(.COVER_INDEX(936)) line_936 (
    .clock(line_936_clock),
    .reset(line_936_reset),
    .valid(line_936_valid)
  );
  GEN_w1_line #(.COVER_INDEX(937)) line_937 (
    .clock(line_937_clock),
    .reset(line_937_reset),
    .valid(line_937_valid)
  );
  GEN_w1_line #(.COVER_INDEX(938)) line_938 (
    .clock(line_938_clock),
    .reset(line_938_reset),
    .valid(line_938_valid)
  );
  GEN_w1_line #(.COVER_INDEX(939)) line_939 (
    .clock(line_939_clock),
    .reset(line_939_reset),
    .valid(line_939_valid)
  );
  GEN_w1_line #(.COVER_INDEX(940)) line_940 (
    .clock(line_940_clock),
    .reset(line_940_reset),
    .valid(line_940_valid)
  );
  GEN_w1_line #(.COVER_INDEX(941)) line_941 (
    .clock(line_941_clock),
    .reset(line_941_reset),
    .valid(line_941_valid)
  );
  GEN_w1_line #(.COVER_INDEX(942)) line_942 (
    .clock(line_942_clock),
    .reset(line_942_reset),
    .valid(line_942_valid)
  );
  GEN_w1_line #(.COVER_INDEX(943)) line_943 (
    .clock(line_943_clock),
    .reset(line_943_reset),
    .valid(line_943_valid)
  );
  GEN_w1_line #(.COVER_INDEX(944)) line_944 (
    .clock(line_944_clock),
    .reset(line_944_reset),
    .valid(line_944_valid)
  );
  GEN_w1_line #(.COVER_INDEX(945)) line_945 (
    .clock(line_945_clock),
    .reset(line_945_reset),
    .valid(line_945_valid)
  );
  GEN_w1_line #(.COVER_INDEX(946)) line_946 (
    .clock(line_946_clock),
    .reset(line_946_reset),
    .valid(line_946_valid)
  );
  GEN_w1_line #(.COVER_INDEX(947)) line_947 (
    .clock(line_947_clock),
    .reset(line_947_reset),
    .valid(line_947_valid)
  );
  GEN_w1_line #(.COVER_INDEX(948)) line_948 (
    .clock(line_948_clock),
    .reset(line_948_reset),
    .valid(line_948_valid)
  );
  GEN_w1_line #(.COVER_INDEX(949)) line_949 (
    .clock(line_949_clock),
    .reset(line_949_reset),
    .valid(line_949_valid)
  );
  GEN_w1_line #(.COVER_INDEX(950)) line_950 (
    .clock(line_950_clock),
    .reset(line_950_reset),
    .valid(line_950_valid)
  );
  GEN_w1_line #(.COVER_INDEX(951)) line_951 (
    .clock(line_951_clock),
    .reset(line_951_reset),
    .valid(line_951_valid)
  );
  GEN_w1_line #(.COVER_INDEX(952)) line_952 (
    .clock(line_952_clock),
    .reset(line_952_reset),
    .valid(line_952_valid)
  );
  GEN_w1_line #(.COVER_INDEX(953)) line_953 (
    .clock(line_953_clock),
    .reset(line_953_reset),
    .valid(line_953_valid)
  );
  GEN_w1_line #(.COVER_INDEX(954)) line_954 (
    .clock(line_954_clock),
    .reset(line_954_reset),
    .valid(line_954_valid)
  );
  GEN_w1_line #(.COVER_INDEX(955)) line_955 (
    .clock(line_955_clock),
    .reset(line_955_reset),
    .valid(line_955_valid)
  );
  GEN_w1_line #(.COVER_INDEX(956)) line_956 (
    .clock(line_956_clock),
    .reset(line_956_reset),
    .valid(line_956_valid)
  );
  GEN_w1_line #(.COVER_INDEX(957)) line_957 (
    .clock(line_957_clock),
    .reset(line_957_reset),
    .valid(line_957_valid)
  );
  GEN_w1_line #(.COVER_INDEX(958)) line_958 (
    .clock(line_958_clock),
    .reset(line_958_reset),
    .valid(line_958_valid)
  );
  GEN_w1_line #(.COVER_INDEX(959)) line_959 (
    .clock(line_959_clock),
    .reset(line_959_reset),
    .valid(line_959_valid)
  );
  GEN_w1_line #(.COVER_INDEX(960)) line_960 (
    .clock(line_960_clock),
    .reset(line_960_reset),
    .valid(line_960_valid)
  );
  GEN_w1_line #(.COVER_INDEX(961)) line_961 (
    .clock(line_961_clock),
    .reset(line_961_reset),
    .valid(line_961_valid)
  );
  GEN_w1_line #(.COVER_INDEX(962)) line_962 (
    .clock(line_962_clock),
    .reset(line_962_reset),
    .valid(line_962_valid)
  );
  GEN_w1_line #(.COVER_INDEX(963)) line_963 (
    .clock(line_963_clock),
    .reset(line_963_reset),
    .valid(line_963_valid)
  );
  GEN_w1_line #(.COVER_INDEX(964)) line_964 (
    .clock(line_964_clock),
    .reset(line_964_reset),
    .valid(line_964_valid)
  );
  GEN_w1_line #(.COVER_INDEX(965)) line_965 (
    .clock(line_965_clock),
    .reset(line_965_reset),
    .valid(line_965_valid)
  );
  GEN_w1_line #(.COVER_INDEX(966)) line_966 (
    .clock(line_966_clock),
    .reset(line_966_reset),
    .valid(line_966_valid)
  );
  GEN_w1_line #(.COVER_INDEX(967)) line_967 (
    .clock(line_967_clock),
    .reset(line_967_reset),
    .valid(line_967_valid)
  );
  GEN_w1_line #(.COVER_INDEX(968)) line_968 (
    .clock(line_968_clock),
    .reset(line_968_reset),
    .valid(line_968_valid)
  );
  GEN_w1_line #(.COVER_INDEX(969)) line_969 (
    .clock(line_969_clock),
    .reset(line_969_reset),
    .valid(line_969_valid)
  );
  GEN_w1_line #(.COVER_INDEX(970)) line_970 (
    .clock(line_970_clock),
    .reset(line_970_reset),
    .valid(line_970_valid)
  );
  GEN_w1_line #(.COVER_INDEX(971)) line_971 (
    .clock(line_971_clock),
    .reset(line_971_reset),
    .valid(line_971_valid)
  );
  GEN_w1_line #(.COVER_INDEX(972)) line_972 (
    .clock(line_972_clock),
    .reset(line_972_reset),
    .valid(line_972_valid)
  );
  GEN_w1_line #(.COVER_INDEX(973)) line_973 (
    .clock(line_973_clock),
    .reset(line_973_reset),
    .valid(line_973_valid)
  );
  GEN_w1_line #(.COVER_INDEX(974)) line_974 (
    .clock(line_974_clock),
    .reset(line_974_reset),
    .valid(line_974_valid)
  );
  GEN_w1_line #(.COVER_INDEX(975)) line_975 (
    .clock(line_975_clock),
    .reset(line_975_reset),
    .valid(line_975_valid)
  );
  GEN_w1_line #(.COVER_INDEX(976)) line_976 (
    .clock(line_976_clock),
    .reset(line_976_reset),
    .valid(line_976_valid)
  );
  GEN_w1_line #(.COVER_INDEX(977)) line_977 (
    .clock(line_977_clock),
    .reset(line_977_reset),
    .valid(line_977_valid)
  );
  GEN_w1_line #(.COVER_INDEX(978)) line_978 (
    .clock(line_978_clock),
    .reset(line_978_reset),
    .valid(line_978_valid)
  );
  GEN_w1_line #(.COVER_INDEX(979)) line_979 (
    .clock(line_979_clock),
    .reset(line_979_reset),
    .valid(line_979_valid)
  );
  GEN_w1_line #(.COVER_INDEX(980)) line_980 (
    .clock(line_980_clock),
    .reset(line_980_reset),
    .valid(line_980_valid)
  );
  GEN_w1_line #(.COVER_INDEX(981)) line_981 (
    .clock(line_981_clock),
    .reset(line_981_reset),
    .valid(line_981_valid)
  );
  GEN_w1_line #(.COVER_INDEX(982)) line_982 (
    .clock(line_982_clock),
    .reset(line_982_reset),
    .valid(line_982_valid)
  );
  GEN_w1_line #(.COVER_INDEX(983)) line_983 (
    .clock(line_983_clock),
    .reset(line_983_reset),
    .valid(line_983_valid)
  );
  GEN_w1_line #(.COVER_INDEX(984)) line_984 (
    .clock(line_984_clock),
    .reset(line_984_reset),
    .valid(line_984_valid)
  );
  GEN_w1_line #(.COVER_INDEX(985)) line_985 (
    .clock(line_985_clock),
    .reset(line_985_reset),
    .valid(line_985_valid)
  );
  GEN_w1_line #(.COVER_INDEX(986)) line_986 (
    .clock(line_986_clock),
    .reset(line_986_reset),
    .valid(line_986_valid)
  );
  GEN_w1_line #(.COVER_INDEX(987)) line_987 (
    .clock(line_987_clock),
    .reset(line_987_reset),
    .valid(line_987_valid)
  );
  GEN_w1_line #(.COVER_INDEX(988)) line_988 (
    .clock(line_988_clock),
    .reset(line_988_reset),
    .valid(line_988_valid)
  );
  GEN_w1_line #(.COVER_INDEX(989)) line_989 (
    .clock(line_989_clock),
    .reset(line_989_reset),
    .valid(line_989_valid)
  );
  GEN_w1_line #(.COVER_INDEX(990)) line_990 (
    .clock(line_990_clock),
    .reset(line_990_reset),
    .valid(line_990_valid)
  );
  GEN_w1_line #(.COVER_INDEX(991)) line_991 (
    .clock(line_991_clock),
    .reset(line_991_reset),
    .valid(line_991_valid)
  );
  GEN_w1_line #(.COVER_INDEX(992)) line_992 (
    .clock(line_992_clock),
    .reset(line_992_reset),
    .valid(line_992_valid)
  );
  GEN_w1_line #(.COVER_INDEX(993)) line_993 (
    .clock(line_993_clock),
    .reset(line_993_reset),
    .valid(line_993_valid)
  );
  GEN_w1_line #(.COVER_INDEX(994)) line_994 (
    .clock(line_994_clock),
    .reset(line_994_reset),
    .valid(line_994_valid)
  );
  GEN_w1_line #(.COVER_INDEX(995)) line_995 (
    .clock(line_995_clock),
    .reset(line_995_reset),
    .valid(line_995_valid)
  );
  GEN_w1_line #(.COVER_INDEX(996)) line_996 (
    .clock(line_996_clock),
    .reset(line_996_reset),
    .valid(line_996_valid)
  );
  GEN_w1_line #(.COVER_INDEX(997)) line_997 (
    .clock(line_997_clock),
    .reset(line_997_reset),
    .valid(line_997_valid)
  );
  GEN_w1_line #(.COVER_INDEX(998)) line_998 (
    .clock(line_998_clock),
    .reset(line_998_reset),
    .valid(line_998_valid)
  );
  GEN_w1_line #(.COVER_INDEX(999)) line_999 (
    .clock(line_999_clock),
    .reset(line_999_reset),
    .valid(line_999_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1000)) line_1000 (
    .clock(line_1000_clock),
    .reset(line_1000_reset),
    .valid(line_1000_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1001)) line_1001 (
    .clock(line_1001_clock),
    .reset(line_1001_reset),
    .valid(line_1001_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1002)) line_1002 (
    .clock(line_1002_clock),
    .reset(line_1002_reset),
    .valid(line_1002_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1003)) line_1003 (
    .clock(line_1003_clock),
    .reset(line_1003_reset),
    .valid(line_1003_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1004)) line_1004 (
    .clock(line_1004_clock),
    .reset(line_1004_reset),
    .valid(line_1004_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1005)) line_1005 (
    .clock(line_1005_clock),
    .reset(line_1005_reset),
    .valid(line_1005_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1006)) line_1006 (
    .clock(line_1006_clock),
    .reset(line_1006_reset),
    .valid(line_1006_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1007)) line_1007 (
    .clock(line_1007_clock),
    .reset(line_1007_reset),
    .valid(line_1007_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1008)) line_1008 (
    .clock(line_1008_clock),
    .reset(line_1008_reset),
    .valid(line_1008_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1009)) line_1009 (
    .clock(line_1009_clock),
    .reset(line_1009_reset),
    .valid(line_1009_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1010)) line_1010 (
    .clock(line_1010_clock),
    .reset(line_1010_reset),
    .valid(line_1010_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1011)) line_1011 (
    .clock(line_1011_clock),
    .reset(line_1011_reset),
    .valid(line_1011_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1012)) line_1012 (
    .clock(line_1012_clock),
    .reset(line_1012_reset),
    .valid(line_1012_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1013)) line_1013 (
    .clock(line_1013_clock),
    .reset(line_1013_reset),
    .valid(line_1013_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1014)) line_1014 (
    .clock(line_1014_clock),
    .reset(line_1014_reset),
    .valid(line_1014_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1015)) line_1015 (
    .clock(line_1015_clock),
    .reset(line_1015_reset),
    .valid(line_1015_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1016)) line_1016 (
    .clock(line_1016_clock),
    .reset(line_1016_reset),
    .valid(line_1016_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1017)) line_1017 (
    .clock(line_1017_clock),
    .reset(line_1017_reset),
    .valid(line_1017_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1018)) line_1018 (
    .clock(line_1018_clock),
    .reset(line_1018_reset),
    .valid(line_1018_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1019)) line_1019 (
    .clock(line_1019_clock),
    .reset(line_1019_reset),
    .valid(line_1019_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1020)) line_1020 (
    .clock(line_1020_clock),
    .reset(line_1020_reset),
    .valid(line_1020_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1021)) line_1021 (
    .clock(line_1021_clock),
    .reset(line_1021_reset),
    .valid(line_1021_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1022)) line_1022 (
    .clock(line_1022_clock),
    .reset(line_1022_reset),
    .valid(line_1022_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1023)) line_1023 (
    .clock(line_1023_clock),
    .reset(line_1023_reset),
    .valid(line_1023_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1024)) line_1024 (
    .clock(line_1024_clock),
    .reset(line_1024_reset),
    .valid(line_1024_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1025)) line_1025 (
    .clock(line_1025_clock),
    .reset(line_1025_reset),
    .valid(line_1025_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1026)) line_1026 (
    .clock(line_1026_clock),
    .reset(line_1026_reset),
    .valid(line_1026_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1027)) line_1027 (
    .clock(line_1027_clock),
    .reset(line_1027_reset),
    .valid(line_1027_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1028)) line_1028 (
    .clock(line_1028_clock),
    .reset(line_1028_reset),
    .valid(line_1028_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1029)) line_1029 (
    .clock(line_1029_clock),
    .reset(line_1029_reset),
    .valid(line_1029_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1030)) line_1030 (
    .clock(line_1030_clock),
    .reset(line_1030_reset),
    .valid(line_1030_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1031)) line_1031 (
    .clock(line_1031_clock),
    .reset(line_1031_reset),
    .valid(line_1031_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1032)) line_1032 (
    .clock(line_1032_clock),
    .reset(line_1032_reset),
    .valid(line_1032_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1033)) line_1033 (
    .clock(line_1033_clock),
    .reset(line_1033_reset),
    .valid(line_1033_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1034)) line_1034 (
    .clock(line_1034_clock),
    .reset(line_1034_reset),
    .valid(line_1034_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1035)) line_1035 (
    .clock(line_1035_clock),
    .reset(line_1035_reset),
    .valid(line_1035_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1036)) line_1036 (
    .clock(line_1036_clock),
    .reset(line_1036_reset),
    .valid(line_1036_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1037)) line_1037 (
    .clock(line_1037_clock),
    .reset(line_1037_reset),
    .valid(line_1037_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1038)) line_1038 (
    .clock(line_1038_clock),
    .reset(line_1038_reset),
    .valid(line_1038_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1039)) line_1039 (
    .clock(line_1039_clock),
    .reset(line_1039_reset),
    .valid(line_1039_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1040)) line_1040 (
    .clock(line_1040_clock),
    .reset(line_1040_reset),
    .valid(line_1040_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1041)) line_1041 (
    .clock(line_1041_clock),
    .reset(line_1041_reset),
    .valid(line_1041_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1042)) line_1042 (
    .clock(line_1042_clock),
    .reset(line_1042_reset),
    .valid(line_1042_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1043)) line_1043 (
    .clock(line_1043_clock),
    .reset(line_1043_reset),
    .valid(line_1043_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1044)) line_1044 (
    .clock(line_1044_clock),
    .reset(line_1044_reset),
    .valid(line_1044_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1045)) line_1045 (
    .clock(line_1045_clock),
    .reset(line_1045_reset),
    .valid(line_1045_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1046)) line_1046 (
    .clock(line_1046_clock),
    .reset(line_1046_reset),
    .valid(line_1046_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1047)) line_1047 (
    .clock(line_1047_clock),
    .reset(line_1047_reset),
    .valid(line_1047_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1048)) line_1048 (
    .clock(line_1048_clock),
    .reset(line_1048_reset),
    .valid(line_1048_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1049)) line_1049 (
    .clock(line_1049_clock),
    .reset(line_1049_reset),
    .valid(line_1049_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1050)) line_1050 (
    .clock(line_1050_clock),
    .reset(line_1050_reset),
    .valid(line_1050_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1051)) line_1051 (
    .clock(line_1051_clock),
    .reset(line_1051_reset),
    .valid(line_1051_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1052)) line_1052 (
    .clock(line_1052_clock),
    .reset(line_1052_reset),
    .valid(line_1052_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1053)) line_1053 (
    .clock(line_1053_clock),
    .reset(line_1053_reset),
    .valid(line_1053_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1054)) line_1054 (
    .clock(line_1054_clock),
    .reset(line_1054_reset),
    .valid(line_1054_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1055)) line_1055 (
    .clock(line_1055_clock),
    .reset(line_1055_reset),
    .valid(line_1055_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1056)) line_1056 (
    .clock(line_1056_clock),
    .reset(line_1056_reset),
    .valid(line_1056_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1057)) line_1057 (
    .clock(line_1057_clock),
    .reset(line_1057_reset),
    .valid(line_1057_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1058)) line_1058 (
    .clock(line_1058_clock),
    .reset(line_1058_reset),
    .valid(line_1058_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1059)) line_1059 (
    .clock(line_1059_clock),
    .reset(line_1059_reset),
    .valid(line_1059_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1060)) line_1060 (
    .clock(line_1060_clock),
    .reset(line_1060_reset),
    .valid(line_1060_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1061)) line_1061 (
    .clock(line_1061_clock),
    .reset(line_1061_reset),
    .valid(line_1061_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1062)) line_1062 (
    .clock(line_1062_clock),
    .reset(line_1062_reset),
    .valid(line_1062_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1063)) line_1063 (
    .clock(line_1063_clock),
    .reset(line_1063_reset),
    .valid(line_1063_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1064)) line_1064 (
    .clock(line_1064_clock),
    .reset(line_1064_reset),
    .valid(line_1064_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1065)) line_1065 (
    .clock(line_1065_clock),
    .reset(line_1065_reset),
    .valid(line_1065_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1066)) line_1066 (
    .clock(line_1066_clock),
    .reset(line_1066_reset),
    .valid(line_1066_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1067)) line_1067 (
    .clock(line_1067_clock),
    .reset(line_1067_reset),
    .valid(line_1067_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1068)) line_1068 (
    .clock(line_1068_clock),
    .reset(line_1068_reset),
    .valid(line_1068_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1069)) line_1069 (
    .clock(line_1069_clock),
    .reset(line_1069_reset),
    .valid(line_1069_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1070)) line_1070 (
    .clock(line_1070_clock),
    .reset(line_1070_reset),
    .valid(line_1070_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1071)) line_1071 (
    .clock(line_1071_clock),
    .reset(line_1071_reset),
    .valid(line_1071_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1072)) line_1072 (
    .clock(line_1072_clock),
    .reset(line_1072_reset),
    .valid(line_1072_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1073)) line_1073 (
    .clock(line_1073_clock),
    .reset(line_1073_reset),
    .valid(line_1073_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1074)) line_1074 (
    .clock(line_1074_clock),
    .reset(line_1074_reset),
    .valid(line_1074_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1075)) line_1075 (
    .clock(line_1075_clock),
    .reset(line_1075_reset),
    .valid(line_1075_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1076)) line_1076 (
    .clock(line_1076_clock),
    .reset(line_1076_reset),
    .valid(line_1076_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1077)) line_1077 (
    .clock(line_1077_clock),
    .reset(line_1077_reset),
    .valid(line_1077_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1078)) line_1078 (
    .clock(line_1078_clock),
    .reset(line_1078_reset),
    .valid(line_1078_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1079)) line_1079 (
    .clock(line_1079_clock),
    .reset(line_1079_reset),
    .valid(line_1079_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1080)) line_1080 (
    .clock(line_1080_clock),
    .reset(line_1080_reset),
    .valid(line_1080_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1081)) line_1081 (
    .clock(line_1081_clock),
    .reset(line_1081_reset),
    .valid(line_1081_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1082)) line_1082 (
    .clock(line_1082_clock),
    .reset(line_1082_reset),
    .valid(line_1082_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1083)) line_1083 (
    .clock(line_1083_clock),
    .reset(line_1083_reset),
    .valid(line_1083_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1084)) line_1084 (
    .clock(line_1084_clock),
    .reset(line_1084_reset),
    .valid(line_1084_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1085)) line_1085 (
    .clock(line_1085_clock),
    .reset(line_1085_reset),
    .valid(line_1085_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1086)) line_1086 (
    .clock(line_1086_clock),
    .reset(line_1086_reset),
    .valid(line_1086_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1087)) line_1087 (
    .clock(line_1087_clock),
    .reset(line_1087_reset),
    .valid(line_1087_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1088)) line_1088 (
    .clock(line_1088_clock),
    .reset(line_1088_reset),
    .valid(line_1088_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1089)) line_1089 (
    .clock(line_1089_clock),
    .reset(line_1089_reset),
    .valid(line_1089_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1090)) line_1090 (
    .clock(line_1090_clock),
    .reset(line_1090_reset),
    .valid(line_1090_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1091)) line_1091 (
    .clock(line_1091_clock),
    .reset(line_1091_reset),
    .valid(line_1091_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1092)) line_1092 (
    .clock(line_1092_clock),
    .reset(line_1092_reset),
    .valid(line_1092_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1093)) line_1093 (
    .clock(line_1093_clock),
    .reset(line_1093_reset),
    .valid(line_1093_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1094)) line_1094 (
    .clock(line_1094_clock),
    .reset(line_1094_reset),
    .valid(line_1094_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1095)) line_1095 (
    .clock(line_1095_clock),
    .reset(line_1095_reset),
    .valid(line_1095_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1096)) line_1096 (
    .clock(line_1096_clock),
    .reset(line_1096_reset),
    .valid(line_1096_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1097)) line_1097 (
    .clock(line_1097_clock),
    .reset(line_1097_reset),
    .valid(line_1097_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1098)) line_1098 (
    .clock(line_1098_clock),
    .reset(line_1098_reset),
    .valid(line_1098_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1099)) line_1099 (
    .clock(line_1099_clock),
    .reset(line_1099_reset),
    .valid(line_1099_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1100)) line_1100 (
    .clock(line_1100_clock),
    .reset(line_1100_reset),
    .valid(line_1100_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1101)) line_1101 (
    .clock(line_1101_clock),
    .reset(line_1101_reset),
    .valid(line_1101_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1102)) line_1102 (
    .clock(line_1102_clock),
    .reset(line_1102_reset),
    .valid(line_1102_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1103)) line_1103 (
    .clock(line_1103_clock),
    .reset(line_1103_reset),
    .valid(line_1103_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1104)) line_1104 (
    .clock(line_1104_clock),
    .reset(line_1104_reset),
    .valid(line_1104_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1105)) line_1105 (
    .clock(line_1105_clock),
    .reset(line_1105_reset),
    .valid(line_1105_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1106)) line_1106 (
    .clock(line_1106_clock),
    .reset(line_1106_reset),
    .valid(line_1106_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1107)) line_1107 (
    .clock(line_1107_clock),
    .reset(line_1107_reset),
    .valid(line_1107_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1108)) line_1108 (
    .clock(line_1108_clock),
    .reset(line_1108_reset),
    .valid(line_1108_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1109)) line_1109 (
    .clock(line_1109_clock),
    .reset(line_1109_reset),
    .valid(line_1109_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1110)) line_1110 (
    .clock(line_1110_clock),
    .reset(line_1110_reset),
    .valid(line_1110_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1111)) line_1111 (
    .clock(line_1111_clock),
    .reset(line_1111_reset),
    .valid(line_1111_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1112)) line_1112 (
    .clock(line_1112_clock),
    .reset(line_1112_reset),
    .valid(line_1112_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1113)) line_1113 (
    .clock(line_1113_clock),
    .reset(line_1113_reset),
    .valid(line_1113_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1114)) line_1114 (
    .clock(line_1114_clock),
    .reset(line_1114_reset),
    .valid(line_1114_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1115)) line_1115 (
    .clock(line_1115_clock),
    .reset(line_1115_reset),
    .valid(line_1115_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1116)) line_1116 (
    .clock(line_1116_clock),
    .reset(line_1116_reset),
    .valid(line_1116_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1117)) line_1117 (
    .clock(line_1117_clock),
    .reset(line_1117_reset),
    .valid(line_1117_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1118)) line_1118 (
    .clock(line_1118_clock),
    .reset(line_1118_reset),
    .valid(line_1118_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1119)) line_1119 (
    .clock(line_1119_clock),
    .reset(line_1119_reset),
    .valid(line_1119_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1120)) line_1120 (
    .clock(line_1120_clock),
    .reset(line_1120_reset),
    .valid(line_1120_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1121)) line_1121 (
    .clock(line_1121_clock),
    .reset(line_1121_reset),
    .valid(line_1121_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1122)) line_1122 (
    .clock(line_1122_clock),
    .reset(line_1122_reset),
    .valid(line_1122_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1123)) line_1123 (
    .clock(line_1123_clock),
    .reset(line_1123_reset),
    .valid(line_1123_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1124)) line_1124 (
    .clock(line_1124_clock),
    .reset(line_1124_reset),
    .valid(line_1124_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1125)) line_1125 (
    .clock(line_1125_clock),
    .reset(line_1125_reset),
    .valid(line_1125_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1126)) line_1126 (
    .clock(line_1126_clock),
    .reset(line_1126_reset),
    .valid(line_1126_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1127)) line_1127 (
    .clock(line_1127_clock),
    .reset(line_1127_reset),
    .valid(line_1127_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1128)) line_1128 (
    .clock(line_1128_clock),
    .reset(line_1128_reset),
    .valid(line_1128_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1129)) line_1129 (
    .clock(line_1129_clock),
    .reset(line_1129_reset),
    .valid(line_1129_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1130)) line_1130 (
    .clock(line_1130_clock),
    .reset(line_1130_reset),
    .valid(line_1130_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1131)) line_1131 (
    .clock(line_1131_clock),
    .reset(line_1131_reset),
    .valid(line_1131_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1132)) line_1132 (
    .clock(line_1132_clock),
    .reset(line_1132_reset),
    .valid(line_1132_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1133)) line_1133 (
    .clock(line_1133_clock),
    .reset(line_1133_reset),
    .valid(line_1133_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1134)) line_1134 (
    .clock(line_1134_clock),
    .reset(line_1134_reset),
    .valid(line_1134_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1135)) line_1135 (
    .clock(line_1135_clock),
    .reset(line_1135_reset),
    .valid(line_1135_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1136)) line_1136 (
    .clock(line_1136_clock),
    .reset(line_1136_reset),
    .valid(line_1136_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1137)) line_1137 (
    .clock(line_1137_clock),
    .reset(line_1137_reset),
    .valid(line_1137_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1138)) line_1138 (
    .clock(line_1138_clock),
    .reset(line_1138_reset),
    .valid(line_1138_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1139)) line_1139 (
    .clock(line_1139_clock),
    .reset(line_1139_reset),
    .valid(line_1139_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1140)) line_1140 (
    .clock(line_1140_clock),
    .reset(line_1140_reset),
    .valid(line_1140_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1141)) line_1141 (
    .clock(line_1141_clock),
    .reset(line_1141_reset),
    .valid(line_1141_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1142)) line_1142 (
    .clock(line_1142_clock),
    .reset(line_1142_reset),
    .valid(line_1142_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1143)) line_1143 (
    .clock(line_1143_clock),
    .reset(line_1143_reset),
    .valid(line_1143_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1144)) line_1144 (
    .clock(line_1144_clock),
    .reset(line_1144_reset),
    .valid(line_1144_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1145)) line_1145 (
    .clock(line_1145_clock),
    .reset(line_1145_reset),
    .valid(line_1145_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1146)) line_1146 (
    .clock(line_1146_clock),
    .reset(line_1146_reset),
    .valid(line_1146_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1147)) line_1147 (
    .clock(line_1147_clock),
    .reset(line_1147_reset),
    .valid(line_1147_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1148)) line_1148 (
    .clock(line_1148_clock),
    .reset(line_1148_reset),
    .valid(line_1148_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1149)) line_1149 (
    .clock(line_1149_clock),
    .reset(line_1149_reset),
    .valid(line_1149_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1150)) line_1150 (
    .clock(line_1150_clock),
    .reset(line_1150_reset),
    .valid(line_1150_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1151)) line_1151 (
    .clock(line_1151_clock),
    .reset(line_1151_reset),
    .valid(line_1151_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1152)) line_1152 (
    .clock(line_1152_clock),
    .reset(line_1152_reset),
    .valid(line_1152_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1153)) line_1153 (
    .clock(line_1153_clock),
    .reset(line_1153_reset),
    .valid(line_1153_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1154)) line_1154 (
    .clock(line_1154_clock),
    .reset(line_1154_reset),
    .valid(line_1154_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1155)) line_1155 (
    .clock(line_1155_clock),
    .reset(line_1155_reset),
    .valid(line_1155_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1156)) line_1156 (
    .clock(line_1156_clock),
    .reset(line_1156_reset),
    .valid(line_1156_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1157)) line_1157 (
    .clock(line_1157_clock),
    .reset(line_1157_reset),
    .valid(line_1157_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1158)) line_1158 (
    .clock(line_1158_clock),
    .reset(line_1158_reset),
    .valid(line_1158_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1159)) line_1159 (
    .clock(line_1159_clock),
    .reset(line_1159_reset),
    .valid(line_1159_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1160)) line_1160 (
    .clock(line_1160_clock),
    .reset(line_1160_reset),
    .valid(line_1160_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1161)) line_1161 (
    .clock(line_1161_clock),
    .reset(line_1161_reset),
    .valid(line_1161_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1162)) line_1162 (
    .clock(line_1162_clock),
    .reset(line_1162_reset),
    .valid(line_1162_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1163)) line_1163 (
    .clock(line_1163_clock),
    .reset(line_1163_reset),
    .valid(line_1163_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1164)) line_1164 (
    .clock(line_1164_clock),
    .reset(line_1164_reset),
    .valid(line_1164_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1165)) line_1165 (
    .clock(line_1165_clock),
    .reset(line_1165_reset),
    .valid(line_1165_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1166)) line_1166 (
    .clock(line_1166_clock),
    .reset(line_1166_reset),
    .valid(line_1166_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1167)) line_1167 (
    .clock(line_1167_clock),
    .reset(line_1167_reset),
    .valid(line_1167_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1168)) line_1168 (
    .clock(line_1168_clock),
    .reset(line_1168_reset),
    .valid(line_1168_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1169)) line_1169 (
    .clock(line_1169_clock),
    .reset(line_1169_reset),
    .valid(line_1169_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1170)) line_1170 (
    .clock(line_1170_clock),
    .reset(line_1170_reset),
    .valid(line_1170_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1171)) line_1171 (
    .clock(line_1171_clock),
    .reset(line_1171_reset),
    .valid(line_1171_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1172)) line_1172 (
    .clock(line_1172_clock),
    .reset(line_1172_reset),
    .valid(line_1172_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1173)) line_1173 (
    .clock(line_1173_clock),
    .reset(line_1173_reset),
    .valid(line_1173_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1174)) line_1174 (
    .clock(line_1174_clock),
    .reset(line_1174_reset),
    .valid(line_1174_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1175)) line_1175 (
    .clock(line_1175_clock),
    .reset(line_1175_reset),
    .valid(line_1175_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1176)) line_1176 (
    .clock(line_1176_clock),
    .reset(line_1176_reset),
    .valid(line_1176_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1177)) line_1177 (
    .clock(line_1177_clock),
    .reset(line_1177_reset),
    .valid(line_1177_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1178)) line_1178 (
    .clock(line_1178_clock),
    .reset(line_1178_reset),
    .valid(line_1178_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1179)) line_1179 (
    .clock(line_1179_clock),
    .reset(line_1179_reset),
    .valid(line_1179_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1180)) line_1180 (
    .clock(line_1180_clock),
    .reset(line_1180_reset),
    .valid(line_1180_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1181)) line_1181 (
    .clock(line_1181_clock),
    .reset(line_1181_reset),
    .valid(line_1181_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1182)) line_1182 (
    .clock(line_1182_clock),
    .reset(line_1182_reset),
    .valid(line_1182_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1183)) line_1183 (
    .clock(line_1183_clock),
    .reset(line_1183_reset),
    .valid(line_1183_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1184)) line_1184 (
    .clock(line_1184_clock),
    .reset(line_1184_reset),
    .valid(line_1184_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1185)) line_1185 (
    .clock(line_1185_clock),
    .reset(line_1185_reset),
    .valid(line_1185_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1186)) line_1186 (
    .clock(line_1186_clock),
    .reset(line_1186_reset),
    .valid(line_1186_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1187)) line_1187 (
    .clock(line_1187_clock),
    .reset(line_1187_reset),
    .valid(line_1187_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1188)) line_1188 (
    .clock(line_1188_clock),
    .reset(line_1188_reset),
    .valid(line_1188_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1189)) line_1189 (
    .clock(line_1189_clock),
    .reset(line_1189_reset),
    .valid(line_1189_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1190)) line_1190 (
    .clock(line_1190_clock),
    .reset(line_1190_reset),
    .valid(line_1190_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1191)) line_1191 (
    .clock(line_1191_clock),
    .reset(line_1191_reset),
    .valid(line_1191_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1192)) line_1192 (
    .clock(line_1192_clock),
    .reset(line_1192_reset),
    .valid(line_1192_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1193)) line_1193 (
    .clock(line_1193_clock),
    .reset(line_1193_reset),
    .valid(line_1193_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1194)) line_1194 (
    .clock(line_1194_clock),
    .reset(line_1194_reset),
    .valid(line_1194_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1195)) line_1195 (
    .clock(line_1195_clock),
    .reset(line_1195_reset),
    .valid(line_1195_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1196)) line_1196 (
    .clock(line_1196_clock),
    .reset(line_1196_reset),
    .valid(line_1196_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1197)) line_1197 (
    .clock(line_1197_clock),
    .reset(line_1197_reset),
    .valid(line_1197_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1198)) line_1198 (
    .clock(line_1198_clock),
    .reset(line_1198_reset),
    .valid(line_1198_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1199)) line_1199 (
    .clock(line_1199_clock),
    .reset(line_1199_reset),
    .valid(line_1199_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1200)) line_1200 (
    .clock(line_1200_clock),
    .reset(line_1200_reset),
    .valid(line_1200_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1201)) line_1201 (
    .clock(line_1201_clock),
    .reset(line_1201_reset),
    .valid(line_1201_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1202)) line_1202 (
    .clock(line_1202_clock),
    .reset(line_1202_reset),
    .valid(line_1202_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1203)) line_1203 (
    .clock(line_1203_clock),
    .reset(line_1203_reset),
    .valid(line_1203_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1204)) line_1204 (
    .clock(line_1204_clock),
    .reset(line_1204_reset),
    .valid(line_1204_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1205)) line_1205 (
    .clock(line_1205_clock),
    .reset(line_1205_reset),
    .valid(line_1205_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1206)) line_1206 (
    .clock(line_1206_clock),
    .reset(line_1206_reset),
    .valid(line_1206_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1207)) line_1207 (
    .clock(line_1207_clock),
    .reset(line_1207_reset),
    .valid(line_1207_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1208)) line_1208 (
    .clock(line_1208_clock),
    .reset(line_1208_reset),
    .valid(line_1208_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1209)) line_1209 (
    .clock(line_1209_clock),
    .reset(line_1209_reset),
    .valid(line_1209_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1210)) line_1210 (
    .clock(line_1210_clock),
    .reset(line_1210_reset),
    .valid(line_1210_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1211)) line_1211 (
    .clock(line_1211_clock),
    .reset(line_1211_reset),
    .valid(line_1211_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1212)) line_1212 (
    .clock(line_1212_clock),
    .reset(line_1212_reset),
    .valid(line_1212_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1213)) line_1213 (
    .clock(line_1213_clock),
    .reset(line_1213_reset),
    .valid(line_1213_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1214)) line_1214 (
    .clock(line_1214_clock),
    .reset(line_1214_reset),
    .valid(line_1214_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1215)) line_1215 (
    .clock(line_1215_clock),
    .reset(line_1215_reset),
    .valid(line_1215_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1216)) line_1216 (
    .clock(line_1216_clock),
    .reset(line_1216_reset),
    .valid(line_1216_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1217)) line_1217 (
    .clock(line_1217_clock),
    .reset(line_1217_reset),
    .valid(line_1217_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1218)) line_1218 (
    .clock(line_1218_clock),
    .reset(line_1218_reset),
    .valid(line_1218_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1219)) line_1219 (
    .clock(line_1219_clock),
    .reset(line_1219_reset),
    .valid(line_1219_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1220)) line_1220 (
    .clock(line_1220_clock),
    .reset(line_1220_reset),
    .valid(line_1220_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1221)) line_1221 (
    .clock(line_1221_clock),
    .reset(line_1221_reset),
    .valid(line_1221_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1222)) line_1222 (
    .clock(line_1222_clock),
    .reset(line_1222_reset),
    .valid(line_1222_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1223)) line_1223 (
    .clock(line_1223_clock),
    .reset(line_1223_reset),
    .valid(line_1223_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1224)) line_1224 (
    .clock(line_1224_clock),
    .reset(line_1224_reset),
    .valid(line_1224_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1225)) line_1225 (
    .clock(line_1225_clock),
    .reset(line_1225_reset),
    .valid(line_1225_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1226)) line_1226 (
    .clock(line_1226_clock),
    .reset(line_1226_reset),
    .valid(line_1226_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1227)) line_1227 (
    .clock(line_1227_clock),
    .reset(line_1227_reset),
    .valid(line_1227_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1228)) line_1228 (
    .clock(line_1228_clock),
    .reset(line_1228_reset),
    .valid(line_1228_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1229)) line_1229 (
    .clock(line_1229_clock),
    .reset(line_1229_reset),
    .valid(line_1229_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1230)) line_1230 (
    .clock(line_1230_clock),
    .reset(line_1230_reset),
    .valid(line_1230_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1231)) line_1231 (
    .clock(line_1231_clock),
    .reset(line_1231_reset),
    .valid(line_1231_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1232)) line_1232 (
    .clock(line_1232_clock),
    .reset(line_1232_reset),
    .valid(line_1232_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1233)) line_1233 (
    .clock(line_1233_clock),
    .reset(line_1233_reset),
    .valid(line_1233_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1234)) line_1234 (
    .clock(line_1234_clock),
    .reset(line_1234_reset),
    .valid(line_1234_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1235)) line_1235 (
    .clock(line_1235_clock),
    .reset(line_1235_reset),
    .valid(line_1235_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1236)) line_1236 (
    .clock(line_1236_clock),
    .reset(line_1236_reset),
    .valid(line_1236_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1237)) line_1237 (
    .clock(line_1237_clock),
    .reset(line_1237_reset),
    .valid(line_1237_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1238)) line_1238 (
    .clock(line_1238_clock),
    .reset(line_1238_reset),
    .valid(line_1238_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1239)) line_1239 (
    .clock(line_1239_clock),
    .reset(line_1239_reset),
    .valid(line_1239_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1240)) line_1240 (
    .clock(line_1240_clock),
    .reset(line_1240_reset),
    .valid(line_1240_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1241)) line_1241 (
    .clock(line_1241_clock),
    .reset(line_1241_reset),
    .valid(line_1241_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1242)) line_1242 (
    .clock(line_1242_clock),
    .reset(line_1242_reset),
    .valid(line_1242_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1243)) line_1243 (
    .clock(line_1243_clock),
    .reset(line_1243_reset),
    .valid(line_1243_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1244)) line_1244 (
    .clock(line_1244_clock),
    .reset(line_1244_reset),
    .valid(line_1244_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1245)) line_1245 (
    .clock(line_1245_clock),
    .reset(line_1245_reset),
    .valid(line_1245_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1246)) line_1246 (
    .clock(line_1246_clock),
    .reset(line_1246_reset),
    .valid(line_1246_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1247)) line_1247 (
    .clock(line_1247_clock),
    .reset(line_1247_reset),
    .valid(line_1247_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1248)) line_1248 (
    .clock(line_1248_clock),
    .reset(line_1248_reset),
    .valid(line_1248_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1249)) line_1249 (
    .clock(line_1249_clock),
    .reset(line_1249_reset),
    .valid(line_1249_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1250)) line_1250 (
    .clock(line_1250_clock),
    .reset(line_1250_reset),
    .valid(line_1250_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1251)) line_1251 (
    .clock(line_1251_clock),
    .reset(line_1251_reset),
    .valid(line_1251_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1252)) line_1252 (
    .clock(line_1252_clock),
    .reset(line_1252_reset),
    .valid(line_1252_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1253)) line_1253 (
    .clock(line_1253_clock),
    .reset(line_1253_reset),
    .valid(line_1253_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1254)) line_1254 (
    .clock(line_1254_clock),
    .reset(line_1254_reset),
    .valid(line_1254_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1255)) line_1255 (
    .clock(line_1255_clock),
    .reset(line_1255_reset),
    .valid(line_1255_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1256)) line_1256 (
    .clock(line_1256_clock),
    .reset(line_1256_reset),
    .valid(line_1256_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1257)) line_1257 (
    .clock(line_1257_clock),
    .reset(line_1257_reset),
    .valid(line_1257_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1258)) line_1258 (
    .clock(line_1258_clock),
    .reset(line_1258_reset),
    .valid(line_1258_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1259)) line_1259 (
    .clock(line_1259_clock),
    .reset(line_1259_reset),
    .valid(line_1259_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1260)) line_1260 (
    .clock(line_1260_clock),
    .reset(line_1260_reset),
    .valid(line_1260_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1261)) line_1261 (
    .clock(line_1261_clock),
    .reset(line_1261_reset),
    .valid(line_1261_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1262)) line_1262 (
    .clock(line_1262_clock),
    .reset(line_1262_reset),
    .valid(line_1262_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1263)) line_1263 (
    .clock(line_1263_clock),
    .reset(line_1263_reset),
    .valid(line_1263_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1264)) line_1264 (
    .clock(line_1264_clock),
    .reset(line_1264_reset),
    .valid(line_1264_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1265)) line_1265 (
    .clock(line_1265_clock),
    .reset(line_1265_reset),
    .valid(line_1265_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1266)) line_1266 (
    .clock(line_1266_clock),
    .reset(line_1266_reset),
    .valid(line_1266_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1267)) line_1267 (
    .clock(line_1267_clock),
    .reset(line_1267_reset),
    .valid(line_1267_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1268)) line_1268 (
    .clock(line_1268_clock),
    .reset(line_1268_reset),
    .valid(line_1268_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1269)) line_1269 (
    .clock(line_1269_clock),
    .reset(line_1269_reset),
    .valid(line_1269_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1270)) line_1270 (
    .clock(line_1270_clock),
    .reset(line_1270_reset),
    .valid(line_1270_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1271)) line_1271 (
    .clock(line_1271_clock),
    .reset(line_1271_reset),
    .valid(line_1271_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1272)) line_1272 (
    .clock(line_1272_clock),
    .reset(line_1272_reset),
    .valid(line_1272_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1273)) line_1273 (
    .clock(line_1273_clock),
    .reset(line_1273_reset),
    .valid(line_1273_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1274)) line_1274 (
    .clock(line_1274_clock),
    .reset(line_1274_reset),
    .valid(line_1274_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1275)) line_1275 (
    .clock(line_1275_clock),
    .reset(line_1275_reset),
    .valid(line_1275_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1276)) line_1276 (
    .clock(line_1276_clock),
    .reset(line_1276_reset),
    .valid(line_1276_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1277)) line_1277 (
    .clock(line_1277_clock),
    .reset(line_1277_reset),
    .valid(line_1277_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1278)) line_1278 (
    .clock(line_1278_clock),
    .reset(line_1278_reset),
    .valid(line_1278_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1279)) line_1279 (
    .clock(line_1279_clock),
    .reset(line_1279_reset),
    .valid(line_1279_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1280)) line_1280 (
    .clock(line_1280_clock),
    .reset(line_1280_reset),
    .valid(line_1280_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1281)) line_1281 (
    .clock(line_1281_clock),
    .reset(line_1281_reset),
    .valid(line_1281_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1282)) line_1282 (
    .clock(line_1282_clock),
    .reset(line_1282_reset),
    .valid(line_1282_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1283)) line_1283 (
    .clock(line_1283_clock),
    .reset(line_1283_reset),
    .valid(line_1283_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1284)) line_1284 (
    .clock(line_1284_clock),
    .reset(line_1284_reset),
    .valid(line_1284_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1285)) line_1285 (
    .clock(line_1285_clock),
    .reset(line_1285_reset),
    .valid(line_1285_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1286)) line_1286 (
    .clock(line_1286_clock),
    .reset(line_1286_reset),
    .valid(line_1286_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1287)) line_1287 (
    .clock(line_1287_clock),
    .reset(line_1287_reset),
    .valid(line_1287_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1288)) line_1288 (
    .clock(line_1288_clock),
    .reset(line_1288_reset),
    .valid(line_1288_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1289)) line_1289 (
    .clock(line_1289_clock),
    .reset(line_1289_reset),
    .valid(line_1289_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1290)) line_1290 (
    .clock(line_1290_clock),
    .reset(line_1290_reset),
    .valid(line_1290_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1291)) line_1291 (
    .clock(line_1291_clock),
    .reset(line_1291_reset),
    .valid(line_1291_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1292)) line_1292 (
    .clock(line_1292_clock),
    .reset(line_1292_reset),
    .valid(line_1292_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1293)) line_1293 (
    .clock(line_1293_clock),
    .reset(line_1293_reset),
    .valid(line_1293_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1294)) line_1294 (
    .clock(line_1294_clock),
    .reset(line_1294_reset),
    .valid(line_1294_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1295)) line_1295 (
    .clock(line_1295_clock),
    .reset(line_1295_reset),
    .valid(line_1295_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1296)) line_1296 (
    .clock(line_1296_clock),
    .reset(line_1296_reset),
    .valid(line_1296_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1297)) line_1297 (
    .clock(line_1297_clock),
    .reset(line_1297_reset),
    .valid(line_1297_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1298)) line_1298 (
    .clock(line_1298_clock),
    .reset(line_1298_reset),
    .valid(line_1298_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1299)) line_1299 (
    .clock(line_1299_clock),
    .reset(line_1299_reset),
    .valid(line_1299_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1300)) line_1300 (
    .clock(line_1300_clock),
    .reset(line_1300_reset),
    .valid(line_1300_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1301)) line_1301 (
    .clock(line_1301_clock),
    .reset(line_1301_reset),
    .valid(line_1301_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1302)) line_1302 (
    .clock(line_1302_clock),
    .reset(line_1302_reset),
    .valid(line_1302_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1303)) line_1303 (
    .clock(line_1303_clock),
    .reset(line_1303_reset),
    .valid(line_1303_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1304)) line_1304 (
    .clock(line_1304_clock),
    .reset(line_1304_reset),
    .valid(line_1304_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1305)) line_1305 (
    .clock(line_1305_clock),
    .reset(line_1305_reset),
    .valid(line_1305_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1306)) line_1306 (
    .clock(line_1306_clock),
    .reset(line_1306_reset),
    .valid(line_1306_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1307)) line_1307 (
    .clock(line_1307_clock),
    .reset(line_1307_reset),
    .valid(line_1307_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1308)) line_1308 (
    .clock(line_1308_clock),
    .reset(line_1308_reset),
    .valid(line_1308_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1309)) line_1309 (
    .clock(line_1309_clock),
    .reset(line_1309_reset),
    .valid(line_1309_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1310)) line_1310 (
    .clock(line_1310_clock),
    .reset(line_1310_reset),
    .valid(line_1310_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1311)) line_1311 (
    .clock(line_1311_clock),
    .reset(line_1311_reset),
    .valid(line_1311_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1312)) line_1312 (
    .clock(line_1312_clock),
    .reset(line_1312_reset),
    .valid(line_1312_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1313)) line_1313 (
    .clock(line_1313_clock),
    .reset(line_1313_reset),
    .valid(line_1313_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1314)) line_1314 (
    .clock(line_1314_clock),
    .reset(line_1314_reset),
    .valid(line_1314_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1315)) line_1315 (
    .clock(line_1315_clock),
    .reset(line_1315_reset),
    .valid(line_1315_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1316)) line_1316 (
    .clock(line_1316_clock),
    .reset(line_1316_reset),
    .valid(line_1316_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1317)) line_1317 (
    .clock(line_1317_clock),
    .reset(line_1317_reset),
    .valid(line_1317_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1318)) line_1318 (
    .clock(line_1318_clock),
    .reset(line_1318_reset),
    .valid(line_1318_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1319)) line_1319 (
    .clock(line_1319_clock),
    .reset(line_1319_reset),
    .valid(line_1319_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1320)) line_1320 (
    .clock(line_1320_clock),
    .reset(line_1320_reset),
    .valid(line_1320_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1321)) line_1321 (
    .clock(line_1321_clock),
    .reset(line_1321_reset),
    .valid(line_1321_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1322)) line_1322 (
    .clock(line_1322_clock),
    .reset(line_1322_reset),
    .valid(line_1322_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1323)) line_1323 (
    .clock(line_1323_clock),
    .reset(line_1323_reset),
    .valid(line_1323_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1324)) line_1324 (
    .clock(line_1324_clock),
    .reset(line_1324_reset),
    .valid(line_1324_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1325)) line_1325 (
    .clock(line_1325_clock),
    .reset(line_1325_reset),
    .valid(line_1325_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1326)) line_1326 (
    .clock(line_1326_clock),
    .reset(line_1326_reset),
    .valid(line_1326_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1327)) line_1327 (
    .clock(line_1327_clock),
    .reset(line_1327_reset),
    .valid(line_1327_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1328)) line_1328 (
    .clock(line_1328_clock),
    .reset(line_1328_reset),
    .valid(line_1328_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1329)) line_1329 (
    .clock(line_1329_clock),
    .reset(line_1329_reset),
    .valid(line_1329_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1330)) line_1330 (
    .clock(line_1330_clock),
    .reset(line_1330_reset),
    .valid(line_1330_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1331)) line_1331 (
    .clock(line_1331_clock),
    .reset(line_1331_reset),
    .valid(line_1331_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1332)) line_1332 (
    .clock(line_1332_clock),
    .reset(line_1332_reset),
    .valid(line_1332_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1333)) line_1333 (
    .clock(line_1333_clock),
    .reset(line_1333_reset),
    .valid(line_1333_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1334)) line_1334 (
    .clock(line_1334_clock),
    .reset(line_1334_reset),
    .valid(line_1334_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1335)) line_1335 (
    .clock(line_1335_clock),
    .reset(line_1335_reset),
    .valid(line_1335_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1336)) line_1336 (
    .clock(line_1336_clock),
    .reset(line_1336_reset),
    .valid(line_1336_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1337)) line_1337 (
    .clock(line_1337_clock),
    .reset(line_1337_reset),
    .valid(line_1337_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1338)) line_1338 (
    .clock(line_1338_clock),
    .reset(line_1338_reset),
    .valid(line_1338_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1339)) line_1339 (
    .clock(line_1339_clock),
    .reset(line_1339_reset),
    .valid(line_1339_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1340)) line_1340 (
    .clock(line_1340_clock),
    .reset(line_1340_reset),
    .valid(line_1340_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1341)) line_1341 (
    .clock(line_1341_clock),
    .reset(line_1341_reset),
    .valid(line_1341_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1342)) line_1342 (
    .clock(line_1342_clock),
    .reset(line_1342_reset),
    .valid(line_1342_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1343)) line_1343 (
    .clock(line_1343_clock),
    .reset(line_1343_reset),
    .valid(line_1343_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1344)) line_1344 (
    .clock(line_1344_clock),
    .reset(line_1344_reset),
    .valid(line_1344_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1345)) line_1345 (
    .clock(line_1345_clock),
    .reset(line_1345_reset),
    .valid(line_1345_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1346)) line_1346 (
    .clock(line_1346_clock),
    .reset(line_1346_reset),
    .valid(line_1346_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1347)) line_1347 (
    .clock(line_1347_clock),
    .reset(line_1347_reset),
    .valid(line_1347_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1348)) line_1348 (
    .clock(line_1348_clock),
    .reset(line_1348_reset),
    .valid(line_1348_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1349)) line_1349 (
    .clock(line_1349_clock),
    .reset(line_1349_reset),
    .valid(line_1349_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1350)) line_1350 (
    .clock(line_1350_clock),
    .reset(line_1350_reset),
    .valid(line_1350_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1351)) line_1351 (
    .clock(line_1351_clock),
    .reset(line_1351_reset),
    .valid(line_1351_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1352)) line_1352 (
    .clock(line_1352_clock),
    .reset(line_1352_reset),
    .valid(line_1352_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1353)) line_1353 (
    .clock(line_1353_clock),
    .reset(line_1353_reset),
    .valid(line_1353_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1354)) line_1354 (
    .clock(line_1354_clock),
    .reset(line_1354_reset),
    .valid(line_1354_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1355)) line_1355 (
    .clock(line_1355_clock),
    .reset(line_1355_reset),
    .valid(line_1355_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1356)) line_1356 (
    .clock(line_1356_clock),
    .reset(line_1356_reset),
    .valid(line_1356_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1357)) line_1357 (
    .clock(line_1357_clock),
    .reset(line_1357_reset),
    .valid(line_1357_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1358)) line_1358 (
    .clock(line_1358_clock),
    .reset(line_1358_reset),
    .valid(line_1358_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1359)) line_1359 (
    .clock(line_1359_clock),
    .reset(line_1359_reset),
    .valid(line_1359_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1360)) line_1360 (
    .clock(line_1360_clock),
    .reset(line_1360_reset),
    .valid(line_1360_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1361)) line_1361 (
    .clock(line_1361_clock),
    .reset(line_1361_reset),
    .valid(line_1361_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1362)) line_1362 (
    .clock(line_1362_clock),
    .reset(line_1362_reset),
    .valid(line_1362_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1363)) line_1363 (
    .clock(line_1363_clock),
    .reset(line_1363_reset),
    .valid(line_1363_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1364)) line_1364 (
    .clock(line_1364_clock),
    .reset(line_1364_reset),
    .valid(line_1364_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1365)) line_1365 (
    .clock(line_1365_clock),
    .reset(line_1365_reset),
    .valid(line_1365_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1366)) line_1366 (
    .clock(line_1366_clock),
    .reset(line_1366_reset),
    .valid(line_1366_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1367)) line_1367 (
    .clock(line_1367_clock),
    .reset(line_1367_reset),
    .valid(line_1367_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1368)) line_1368 (
    .clock(line_1368_clock),
    .reset(line_1368_reset),
    .valid(line_1368_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1369)) line_1369 (
    .clock(line_1369_clock),
    .reset(line_1369_reset),
    .valid(line_1369_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1370)) line_1370 (
    .clock(line_1370_clock),
    .reset(line_1370_reset),
    .valid(line_1370_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1371)) line_1371 (
    .clock(line_1371_clock),
    .reset(line_1371_reset),
    .valid(line_1371_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1372)) line_1372 (
    .clock(line_1372_clock),
    .reset(line_1372_reset),
    .valid(line_1372_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1373)) line_1373 (
    .clock(line_1373_clock),
    .reset(line_1373_reset),
    .valid(line_1373_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1374)) line_1374 (
    .clock(line_1374_clock),
    .reset(line_1374_reset),
    .valid(line_1374_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1375)) line_1375 (
    .clock(line_1375_clock),
    .reset(line_1375_reset),
    .valid(line_1375_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1376)) line_1376 (
    .clock(line_1376_clock),
    .reset(line_1376_reset),
    .valid(line_1376_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1377)) line_1377 (
    .clock(line_1377_clock),
    .reset(line_1377_reset),
    .valid(line_1377_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1378)) line_1378 (
    .clock(line_1378_clock),
    .reset(line_1378_reset),
    .valid(line_1378_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1379)) line_1379 (
    .clock(line_1379_clock),
    .reset(line_1379_reset),
    .valid(line_1379_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1380)) line_1380 (
    .clock(line_1380_clock),
    .reset(line_1380_reset),
    .valid(line_1380_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1381)) line_1381 (
    .clock(line_1381_clock),
    .reset(line_1381_reset),
    .valid(line_1381_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1382)) line_1382 (
    .clock(line_1382_clock),
    .reset(line_1382_reset),
    .valid(line_1382_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1383)) line_1383 (
    .clock(line_1383_clock),
    .reset(line_1383_reset),
    .valid(line_1383_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1384)) line_1384 (
    .clock(line_1384_clock),
    .reset(line_1384_reset),
    .valid(line_1384_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1385)) line_1385 (
    .clock(line_1385_clock),
    .reset(line_1385_reset),
    .valid(line_1385_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1386)) line_1386 (
    .clock(line_1386_clock),
    .reset(line_1386_reset),
    .valid(line_1386_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1387)) line_1387 (
    .clock(line_1387_clock),
    .reset(line_1387_reset),
    .valid(line_1387_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1388)) line_1388 (
    .clock(line_1388_clock),
    .reset(line_1388_reset),
    .valid(line_1388_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1389)) line_1389 (
    .clock(line_1389_clock),
    .reset(line_1389_reset),
    .valid(line_1389_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1390)) line_1390 (
    .clock(line_1390_clock),
    .reset(line_1390_reset),
    .valid(line_1390_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1391)) line_1391 (
    .clock(line_1391_clock),
    .reset(line_1391_reset),
    .valid(line_1391_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1392)) line_1392 (
    .clock(line_1392_clock),
    .reset(line_1392_reset),
    .valid(line_1392_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1393)) line_1393 (
    .clock(line_1393_clock),
    .reset(line_1393_reset),
    .valid(line_1393_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1394)) line_1394 (
    .clock(line_1394_clock),
    .reset(line_1394_reset),
    .valid(line_1394_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1395)) line_1395 (
    .clock(line_1395_clock),
    .reset(line_1395_reset),
    .valid(line_1395_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1396)) line_1396 (
    .clock(line_1396_clock),
    .reset(line_1396_reset),
    .valid(line_1396_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1397)) line_1397 (
    .clock(line_1397_clock),
    .reset(line_1397_reset),
    .valid(line_1397_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1398)) line_1398 (
    .clock(line_1398_clock),
    .reset(line_1398_reset),
    .valid(line_1398_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1399)) line_1399 (
    .clock(line_1399_clock),
    .reset(line_1399_reset),
    .valid(line_1399_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1400)) line_1400 (
    .clock(line_1400_clock),
    .reset(line_1400_reset),
    .valid(line_1400_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1401)) line_1401 (
    .clock(line_1401_clock),
    .reset(line_1401_reset),
    .valid(line_1401_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1402)) line_1402 (
    .clock(line_1402_clock),
    .reset(line_1402_reset),
    .valid(line_1402_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1403)) line_1403 (
    .clock(line_1403_clock),
    .reset(line_1403_reset),
    .valid(line_1403_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1404)) line_1404 (
    .clock(line_1404_clock),
    .reset(line_1404_reset),
    .valid(line_1404_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1405)) line_1405 (
    .clock(line_1405_clock),
    .reset(line_1405_reset),
    .valid(line_1405_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1406)) line_1406 (
    .clock(line_1406_clock),
    .reset(line_1406_reset),
    .valid(line_1406_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1407)) line_1407 (
    .clock(line_1407_clock),
    .reset(line_1407_reset),
    .valid(line_1407_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1408)) line_1408 (
    .clock(line_1408_clock),
    .reset(line_1408_reset),
    .valid(line_1408_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1409)) line_1409 (
    .clock(line_1409_clock),
    .reset(line_1409_reset),
    .valid(line_1409_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1410)) line_1410 (
    .clock(line_1410_clock),
    .reset(line_1410_reset),
    .valid(line_1410_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1411)) line_1411 (
    .clock(line_1411_clock),
    .reset(line_1411_reset),
    .valid(line_1411_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1412)) line_1412 (
    .clock(line_1412_clock),
    .reset(line_1412_reset),
    .valid(line_1412_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1413)) line_1413 (
    .clock(line_1413_clock),
    .reset(line_1413_reset),
    .valid(line_1413_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1414)) line_1414 (
    .clock(line_1414_clock),
    .reset(line_1414_reset),
    .valid(line_1414_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1415)) line_1415 (
    .clock(line_1415_clock),
    .reset(line_1415_reset),
    .valid(line_1415_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1416)) line_1416 (
    .clock(line_1416_clock),
    .reset(line_1416_reset),
    .valid(line_1416_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1417)) line_1417 (
    .clock(line_1417_clock),
    .reset(line_1417_reset),
    .valid(line_1417_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1418)) line_1418 (
    .clock(line_1418_clock),
    .reset(line_1418_reset),
    .valid(line_1418_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1419)) line_1419 (
    .clock(line_1419_clock),
    .reset(line_1419_reset),
    .valid(line_1419_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1420)) line_1420 (
    .clock(line_1420_clock),
    .reset(line_1420_reset),
    .valid(line_1420_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1421)) line_1421 (
    .clock(line_1421_clock),
    .reset(line_1421_reset),
    .valid(line_1421_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1422)) line_1422 (
    .clock(line_1422_clock),
    .reset(line_1422_reset),
    .valid(line_1422_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1423)) line_1423 (
    .clock(line_1423_clock),
    .reset(line_1423_reset),
    .valid(line_1423_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1424)) line_1424 (
    .clock(line_1424_clock),
    .reset(line_1424_reset),
    .valid(line_1424_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1425)) line_1425 (
    .clock(line_1425_clock),
    .reset(line_1425_reset),
    .valid(line_1425_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1426)) line_1426 (
    .clock(line_1426_clock),
    .reset(line_1426_reset),
    .valid(line_1426_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1427)) line_1427 (
    .clock(line_1427_clock),
    .reset(line_1427_reset),
    .valid(line_1427_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1428)) line_1428 (
    .clock(line_1428_clock),
    .reset(line_1428_reset),
    .valid(line_1428_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1429)) line_1429 (
    .clock(line_1429_clock),
    .reset(line_1429_reset),
    .valid(line_1429_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1430)) line_1430 (
    .clock(line_1430_clock),
    .reset(line_1430_reset),
    .valid(line_1430_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1431)) line_1431 (
    .clock(line_1431_clock),
    .reset(line_1431_reset),
    .valid(line_1431_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1432)) line_1432 (
    .clock(line_1432_clock),
    .reset(line_1432_reset),
    .valid(line_1432_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1433)) line_1433 (
    .clock(line_1433_clock),
    .reset(line_1433_reset),
    .valid(line_1433_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1434)) line_1434 (
    .clock(line_1434_clock),
    .reset(line_1434_reset),
    .valid(line_1434_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1435)) line_1435 (
    .clock(line_1435_clock),
    .reset(line_1435_reset),
    .valid(line_1435_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1436)) line_1436 (
    .clock(line_1436_clock),
    .reset(line_1436_reset),
    .valid(line_1436_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1437)) line_1437 (
    .clock(line_1437_clock),
    .reset(line_1437_reset),
    .valid(line_1437_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1438)) line_1438 (
    .clock(line_1438_clock),
    .reset(line_1438_reset),
    .valid(line_1438_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1439)) line_1439 (
    .clock(line_1439_clock),
    .reset(line_1439_reset),
    .valid(line_1439_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1440)) line_1440 (
    .clock(line_1440_clock),
    .reset(line_1440_reset),
    .valid(line_1440_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1441)) line_1441 (
    .clock(line_1441_clock),
    .reset(line_1441_reset),
    .valid(line_1441_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1442)) line_1442 (
    .clock(line_1442_clock),
    .reset(line_1442_reset),
    .valid(line_1442_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1443)) line_1443 (
    .clock(line_1443_clock),
    .reset(line_1443_reset),
    .valid(line_1443_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1444)) line_1444 (
    .clock(line_1444_clock),
    .reset(line_1444_reset),
    .valid(line_1444_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1445)) line_1445 (
    .clock(line_1445_clock),
    .reset(line_1445_reset),
    .valid(line_1445_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1446)) line_1446 (
    .clock(line_1446_clock),
    .reset(line_1446_reset),
    .valid(line_1446_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1447)) line_1447 (
    .clock(line_1447_clock),
    .reset(line_1447_reset),
    .valid(line_1447_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1448)) line_1448 (
    .clock(line_1448_clock),
    .reset(line_1448_reset),
    .valid(line_1448_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1449)) line_1449 (
    .clock(line_1449_clock),
    .reset(line_1449_reset),
    .valid(line_1449_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1450)) line_1450 (
    .clock(line_1450_clock),
    .reset(line_1450_reset),
    .valid(line_1450_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1451)) line_1451 (
    .clock(line_1451_clock),
    .reset(line_1451_reset),
    .valid(line_1451_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1452)) line_1452 (
    .clock(line_1452_clock),
    .reset(line_1452_reset),
    .valid(line_1452_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1453)) line_1453 (
    .clock(line_1453_clock),
    .reset(line_1453_reset),
    .valid(line_1453_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1454)) line_1454 (
    .clock(line_1454_clock),
    .reset(line_1454_reset),
    .valid(line_1454_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1455)) line_1455 (
    .clock(line_1455_clock),
    .reset(line_1455_reset),
    .valid(line_1455_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1456)) line_1456 (
    .clock(line_1456_clock),
    .reset(line_1456_reset),
    .valid(line_1456_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1457)) line_1457 (
    .clock(line_1457_clock),
    .reset(line_1457_reset),
    .valid(line_1457_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1458)) line_1458 (
    .clock(line_1458_clock),
    .reset(line_1458_reset),
    .valid(line_1458_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1459)) line_1459 (
    .clock(line_1459_clock),
    .reset(line_1459_reset),
    .valid(line_1459_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1460)) line_1460 (
    .clock(line_1460_clock),
    .reset(line_1460_reset),
    .valid(line_1460_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1461)) line_1461 (
    .clock(line_1461_clock),
    .reset(line_1461_reset),
    .valid(line_1461_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1462)) line_1462 (
    .clock(line_1462_clock),
    .reset(line_1462_reset),
    .valid(line_1462_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1463)) line_1463 (
    .clock(line_1463_clock),
    .reset(line_1463_reset),
    .valid(line_1463_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1464)) line_1464 (
    .clock(line_1464_clock),
    .reset(line_1464_reset),
    .valid(line_1464_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1465)) line_1465 (
    .clock(line_1465_clock),
    .reset(line_1465_reset),
    .valid(line_1465_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1466)) line_1466 (
    .clock(line_1466_clock),
    .reset(line_1466_reset),
    .valid(line_1466_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1467)) line_1467 (
    .clock(line_1467_clock),
    .reset(line_1467_reset),
    .valid(line_1467_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1468)) line_1468 (
    .clock(line_1468_clock),
    .reset(line_1468_reset),
    .valid(line_1468_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1469)) line_1469 (
    .clock(line_1469_clock),
    .reset(line_1469_reset),
    .valid(line_1469_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1470)) line_1470 (
    .clock(line_1470_clock),
    .reset(line_1470_reset),
    .valid(line_1470_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1471)) line_1471 (
    .clock(line_1471_clock),
    .reset(line_1471_reset),
    .valid(line_1471_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1472)) line_1472 (
    .clock(line_1472_clock),
    .reset(line_1472_reset),
    .valid(line_1472_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1473)) line_1473 (
    .clock(line_1473_clock),
    .reset(line_1473_reset),
    .valid(line_1473_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1474)) line_1474 (
    .clock(line_1474_clock),
    .reset(line_1474_reset),
    .valid(line_1474_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1475)) line_1475 (
    .clock(line_1475_clock),
    .reset(line_1475_reset),
    .valid(line_1475_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1476)) line_1476 (
    .clock(line_1476_clock),
    .reset(line_1476_reset),
    .valid(line_1476_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1477)) line_1477 (
    .clock(line_1477_clock),
    .reset(line_1477_reset),
    .valid(line_1477_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1478)) line_1478 (
    .clock(line_1478_clock),
    .reset(line_1478_reset),
    .valid(line_1478_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1479)) line_1479 (
    .clock(line_1479_clock),
    .reset(line_1479_reset),
    .valid(line_1479_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1480)) line_1480 (
    .clock(line_1480_clock),
    .reset(line_1480_reset),
    .valid(line_1480_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1481)) line_1481 (
    .clock(line_1481_clock),
    .reset(line_1481_reset),
    .valid(line_1481_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1482)) line_1482 (
    .clock(line_1482_clock),
    .reset(line_1482_reset),
    .valid(line_1482_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1483)) line_1483 (
    .clock(line_1483_clock),
    .reset(line_1483_reset),
    .valid(line_1483_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1484)) line_1484 (
    .clock(line_1484_clock),
    .reset(line_1484_reset),
    .valid(line_1484_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1485)) line_1485 (
    .clock(line_1485_clock),
    .reset(line_1485_reset),
    .valid(line_1485_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1486)) line_1486 (
    .clock(line_1486_clock),
    .reset(line_1486_reset),
    .valid(line_1486_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1487)) line_1487 (
    .clock(line_1487_clock),
    .reset(line_1487_reset),
    .valid(line_1487_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1488)) line_1488 (
    .clock(line_1488_clock),
    .reset(line_1488_reset),
    .valid(line_1488_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1489)) line_1489 (
    .clock(line_1489_clock),
    .reset(line_1489_reset),
    .valid(line_1489_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1490)) line_1490 (
    .clock(line_1490_clock),
    .reset(line_1490_reset),
    .valid(line_1490_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1491)) line_1491 (
    .clock(line_1491_clock),
    .reset(line_1491_reset),
    .valid(line_1491_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1492)) line_1492 (
    .clock(line_1492_clock),
    .reset(line_1492_reset),
    .valid(line_1492_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1493)) line_1493 (
    .clock(line_1493_clock),
    .reset(line_1493_reset),
    .valid(line_1493_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1494)) line_1494 (
    .clock(line_1494_clock),
    .reset(line_1494_reset),
    .valid(line_1494_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1495)) line_1495 (
    .clock(line_1495_clock),
    .reset(line_1495_reset),
    .valid(line_1495_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1496)) line_1496 (
    .clock(line_1496_clock),
    .reset(line_1496_reset),
    .valid(line_1496_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1497)) line_1497 (
    .clock(line_1497_clock),
    .reset(line_1497_reset),
    .valid(line_1497_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1498)) line_1498 (
    .clock(line_1498_clock),
    .reset(line_1498_reset),
    .valid(line_1498_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1499)) line_1499 (
    .clock(line_1499_clock),
    .reset(line_1499_reset),
    .valid(line_1499_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1500)) line_1500 (
    .clock(line_1500_clock),
    .reset(line_1500_reset),
    .valid(line_1500_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1501)) line_1501 (
    .clock(line_1501_clock),
    .reset(line_1501_reset),
    .valid(line_1501_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1502)) line_1502 (
    .clock(line_1502_clock),
    .reset(line_1502_reset),
    .valid(line_1502_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1503)) line_1503 (
    .clock(line_1503_clock),
    .reset(line_1503_reset),
    .valid(line_1503_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1504)) line_1504 (
    .clock(line_1504_clock),
    .reset(line_1504_reset),
    .valid(line_1504_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1505)) line_1505 (
    .clock(line_1505_clock),
    .reset(line_1505_reset),
    .valid(line_1505_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1506)) line_1506 (
    .clock(line_1506_clock),
    .reset(line_1506_reset),
    .valid(line_1506_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1507)) line_1507 (
    .clock(line_1507_clock),
    .reset(line_1507_reset),
    .valid(line_1507_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1508)) line_1508 (
    .clock(line_1508_clock),
    .reset(line_1508_reset),
    .valid(line_1508_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1509)) line_1509 (
    .clock(line_1509_clock),
    .reset(line_1509_reset),
    .valid(line_1509_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1510)) line_1510 (
    .clock(line_1510_clock),
    .reset(line_1510_reset),
    .valid(line_1510_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1511)) line_1511 (
    .clock(line_1511_clock),
    .reset(line_1511_reset),
    .valid(line_1511_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1512)) line_1512 (
    .clock(line_1512_clock),
    .reset(line_1512_reset),
    .valid(line_1512_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1513)) line_1513 (
    .clock(line_1513_clock),
    .reset(line_1513_reset),
    .valid(line_1513_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1514)) line_1514 (
    .clock(line_1514_clock),
    .reset(line_1514_reset),
    .valid(line_1514_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1515)) line_1515 (
    .clock(line_1515_clock),
    .reset(line_1515_reset),
    .valid(line_1515_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1516)) line_1516 (
    .clock(line_1516_clock),
    .reset(line_1516_reset),
    .valid(line_1516_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1517)) line_1517 (
    .clock(line_1517_clock),
    .reset(line_1517_reset),
    .valid(line_1517_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1518)) line_1518 (
    .clock(line_1518_clock),
    .reset(line_1518_reset),
    .valid(line_1518_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1519)) line_1519 (
    .clock(line_1519_clock),
    .reset(line_1519_reset),
    .valid(line_1519_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1520)) line_1520 (
    .clock(line_1520_clock),
    .reset(line_1520_reset),
    .valid(line_1520_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1521)) line_1521 (
    .clock(line_1521_clock),
    .reset(line_1521_reset),
    .valid(line_1521_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1522)) line_1522 (
    .clock(line_1522_clock),
    .reset(line_1522_reset),
    .valid(line_1522_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1523)) line_1523 (
    .clock(line_1523_clock),
    .reset(line_1523_reset),
    .valid(line_1523_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1524)) line_1524 (
    .clock(line_1524_clock),
    .reset(line_1524_reset),
    .valid(line_1524_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1525)) line_1525 (
    .clock(line_1525_clock),
    .reset(line_1525_reset),
    .valid(line_1525_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1526)) line_1526 (
    .clock(line_1526_clock),
    .reset(line_1526_reset),
    .valid(line_1526_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1527)) line_1527 (
    .clock(line_1527_clock),
    .reset(line_1527_reset),
    .valid(line_1527_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1528)) line_1528 (
    .clock(line_1528_clock),
    .reset(line_1528_reset),
    .valid(line_1528_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1529)) line_1529 (
    .clock(line_1529_clock),
    .reset(line_1529_reset),
    .valid(line_1529_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1530)) line_1530 (
    .clock(line_1530_clock),
    .reset(line_1530_reset),
    .valid(line_1530_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1531)) line_1531 (
    .clock(line_1531_clock),
    .reset(line_1531_reset),
    .valid(line_1531_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1532)) line_1532 (
    .clock(line_1532_clock),
    .reset(line_1532_reset),
    .valid(line_1532_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1533)) line_1533 (
    .clock(line_1533_clock),
    .reset(line_1533_reset),
    .valid(line_1533_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1534)) line_1534 (
    .clock(line_1534_clock),
    .reset(line_1534_reset),
    .valid(line_1534_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1535)) line_1535 (
    .clock(line_1535_clock),
    .reset(line_1535_reset),
    .valid(line_1535_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1536)) line_1536 (
    .clock(line_1536_clock),
    .reset(line_1536_reset),
    .valid(line_1536_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1537)) line_1537 (
    .clock(line_1537_clock),
    .reset(line_1537_reset),
    .valid(line_1537_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1538)) line_1538 (
    .clock(line_1538_clock),
    .reset(line_1538_reset),
    .valid(line_1538_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1539)) line_1539 (
    .clock(line_1539_clock),
    .reset(line_1539_reset),
    .valid(line_1539_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1540)) line_1540 (
    .clock(line_1540_clock),
    .reset(line_1540_reset),
    .valid(line_1540_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1541)) line_1541 (
    .clock(line_1541_clock),
    .reset(line_1541_reset),
    .valid(line_1541_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1542)) line_1542 (
    .clock(line_1542_clock),
    .reset(line_1542_reset),
    .valid(line_1542_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1543)) line_1543 (
    .clock(line_1543_clock),
    .reset(line_1543_reset),
    .valid(line_1543_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1544)) line_1544 (
    .clock(line_1544_clock),
    .reset(line_1544_reset),
    .valid(line_1544_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1545)) line_1545 (
    .clock(line_1545_clock),
    .reset(line_1545_reset),
    .valid(line_1545_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1546)) line_1546 (
    .clock(line_1546_clock),
    .reset(line_1546_reset),
    .valid(line_1546_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1547)) line_1547 (
    .clock(line_1547_clock),
    .reset(line_1547_reset),
    .valid(line_1547_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1548)) line_1548 (
    .clock(line_1548_clock),
    .reset(line_1548_reset),
    .valid(line_1548_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1549)) line_1549 (
    .clock(line_1549_clock),
    .reset(line_1549_reset),
    .valid(line_1549_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1550)) line_1550 (
    .clock(line_1550_clock),
    .reset(line_1550_reset),
    .valid(line_1550_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1551)) line_1551 (
    .clock(line_1551_clock),
    .reset(line_1551_reset),
    .valid(line_1551_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1552)) line_1552 (
    .clock(line_1552_clock),
    .reset(line_1552_reset),
    .valid(line_1552_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1553)) line_1553 (
    .clock(line_1553_clock),
    .reset(line_1553_reset),
    .valid(line_1553_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1554)) line_1554 (
    .clock(line_1554_clock),
    .reset(line_1554_reset),
    .valid(line_1554_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1555)) line_1555 (
    .clock(line_1555_clock),
    .reset(line_1555_reset),
    .valid(line_1555_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1556)) line_1556 (
    .clock(line_1556_clock),
    .reset(line_1556_reset),
    .valid(line_1556_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1557)) line_1557 (
    .clock(line_1557_clock),
    .reset(line_1557_reset),
    .valid(line_1557_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1558)) line_1558 (
    .clock(line_1558_clock),
    .reset(line_1558_reset),
    .valid(line_1558_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1559)) line_1559 (
    .clock(line_1559_clock),
    .reset(line_1559_reset),
    .valid(line_1559_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1560)) line_1560 (
    .clock(line_1560_clock),
    .reset(line_1560_reset),
    .valid(line_1560_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1561)) line_1561 (
    .clock(line_1561_clock),
    .reset(line_1561_reset),
    .valid(line_1561_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1562)) line_1562 (
    .clock(line_1562_clock),
    .reset(line_1562_reset),
    .valid(line_1562_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1563)) line_1563 (
    .clock(line_1563_clock),
    .reset(line_1563_reset),
    .valid(line_1563_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1564)) line_1564 (
    .clock(line_1564_clock),
    .reset(line_1564_reset),
    .valid(line_1564_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1565)) line_1565 (
    .clock(line_1565_clock),
    .reset(line_1565_reset),
    .valid(line_1565_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1566)) line_1566 (
    .clock(line_1566_clock),
    .reset(line_1566_reset),
    .valid(line_1566_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1567)) line_1567 (
    .clock(line_1567_clock),
    .reset(line_1567_reset),
    .valid(line_1567_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1568)) line_1568 (
    .clock(line_1568_clock),
    .reset(line_1568_reset),
    .valid(line_1568_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1569)) line_1569 (
    .clock(line_1569_clock),
    .reset(line_1569_reset),
    .valid(line_1569_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1570)) line_1570 (
    .clock(line_1570_clock),
    .reset(line_1570_reset),
    .valid(line_1570_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1571)) line_1571 (
    .clock(line_1571_clock),
    .reset(line_1571_reset),
    .valid(line_1571_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1572)) line_1572 (
    .clock(line_1572_clock),
    .reset(line_1572_reset),
    .valid(line_1572_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1573)) line_1573 (
    .clock(line_1573_clock),
    .reset(line_1573_reset),
    .valid(line_1573_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1574)) line_1574 (
    .clock(line_1574_clock),
    .reset(line_1574_reset),
    .valid(line_1574_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1575)) line_1575 (
    .clock(line_1575_clock),
    .reset(line_1575_reset),
    .valid(line_1575_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1576)) line_1576 (
    .clock(line_1576_clock),
    .reset(line_1576_reset),
    .valid(line_1576_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1577)) line_1577 (
    .clock(line_1577_clock),
    .reset(line_1577_reset),
    .valid(line_1577_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1578)) line_1578 (
    .clock(line_1578_clock),
    .reset(line_1578_reset),
    .valid(line_1578_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1579)) line_1579 (
    .clock(line_1579_clock),
    .reset(line_1579_reset),
    .valid(line_1579_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1580)) line_1580 (
    .clock(line_1580_clock),
    .reset(line_1580_reset),
    .valid(line_1580_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1581)) line_1581 (
    .clock(line_1581_clock),
    .reset(line_1581_reset),
    .valid(line_1581_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1582)) line_1582 (
    .clock(line_1582_clock),
    .reset(line_1582_reset),
    .valid(line_1582_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1583)) line_1583 (
    .clock(line_1583_clock),
    .reset(line_1583_reset),
    .valid(line_1583_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1584)) line_1584 (
    .clock(line_1584_clock),
    .reset(line_1584_reset),
    .valid(line_1584_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1585)) line_1585 (
    .clock(line_1585_clock),
    .reset(line_1585_reset),
    .valid(line_1585_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1586)) line_1586 (
    .clock(line_1586_clock),
    .reset(line_1586_reset),
    .valid(line_1586_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1587)) line_1587 (
    .clock(line_1587_clock),
    .reset(line_1587_reset),
    .valid(line_1587_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1588)) line_1588 (
    .clock(line_1588_clock),
    .reset(line_1588_reset),
    .valid(line_1588_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1589)) line_1589 (
    .clock(line_1589_clock),
    .reset(line_1589_reset),
    .valid(line_1589_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1590)) line_1590 (
    .clock(line_1590_clock),
    .reset(line_1590_reset),
    .valid(line_1590_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1591)) line_1591 (
    .clock(line_1591_clock),
    .reset(line_1591_reset),
    .valid(line_1591_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1592)) line_1592 (
    .clock(line_1592_clock),
    .reset(line_1592_reset),
    .valid(line_1592_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1593)) line_1593 (
    .clock(line_1593_clock),
    .reset(line_1593_reset),
    .valid(line_1593_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1594)) line_1594 (
    .clock(line_1594_clock),
    .reset(line_1594_reset),
    .valid(line_1594_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1595)) line_1595 (
    .clock(line_1595_clock),
    .reset(line_1595_reset),
    .valid(line_1595_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1596)) line_1596 (
    .clock(line_1596_clock),
    .reset(line_1596_reset),
    .valid(line_1596_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1597)) line_1597 (
    .clock(line_1597_clock),
    .reset(line_1597_reset),
    .valid(line_1597_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1598)) line_1598 (
    .clock(line_1598_clock),
    .reset(line_1598_reset),
    .valid(line_1598_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1599)) line_1599 (
    .clock(line_1599_clock),
    .reset(line_1599_reset),
    .valid(line_1599_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1600)) line_1600 (
    .clock(line_1600_clock),
    .reset(line_1600_reset),
    .valid(line_1600_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1601)) line_1601 (
    .clock(line_1601_clock),
    .reset(line_1601_reset),
    .valid(line_1601_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1602)) line_1602 (
    .clock(line_1602_clock),
    .reset(line_1602_reset),
    .valid(line_1602_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1603)) line_1603 (
    .clock(line_1603_clock),
    .reset(line_1603_reset),
    .valid(line_1603_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1604)) line_1604 (
    .clock(line_1604_clock),
    .reset(line_1604_reset),
    .valid(line_1604_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1605)) line_1605 (
    .clock(line_1605_clock),
    .reset(line_1605_reset),
    .valid(line_1605_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1606)) line_1606 (
    .clock(line_1606_clock),
    .reset(line_1606_reset),
    .valid(line_1606_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1607)) line_1607 (
    .clock(line_1607_clock),
    .reset(line_1607_reset),
    .valid(line_1607_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1608)) line_1608 (
    .clock(line_1608_clock),
    .reset(line_1608_reset),
    .valid(line_1608_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1609)) line_1609 (
    .clock(line_1609_clock),
    .reset(line_1609_reset),
    .valid(line_1609_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1610)) line_1610 (
    .clock(line_1610_clock),
    .reset(line_1610_reset),
    .valid(line_1610_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1611)) line_1611 (
    .clock(line_1611_clock),
    .reset(line_1611_reset),
    .valid(line_1611_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1612)) line_1612 (
    .clock(line_1612_clock),
    .reset(line_1612_reset),
    .valid(line_1612_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1613)) line_1613 (
    .clock(line_1613_clock),
    .reset(line_1613_reset),
    .valid(line_1613_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1614)) line_1614 (
    .clock(line_1614_clock),
    .reset(line_1614_reset),
    .valid(line_1614_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1615)) line_1615 (
    .clock(line_1615_clock),
    .reset(line_1615_reset),
    .valid(line_1615_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1616)) line_1616 (
    .clock(line_1616_clock),
    .reset(line_1616_reset),
    .valid(line_1616_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1617)) line_1617 (
    .clock(line_1617_clock),
    .reset(line_1617_reset),
    .valid(line_1617_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1618)) line_1618 (
    .clock(line_1618_clock),
    .reset(line_1618_reset),
    .valid(line_1618_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1619)) line_1619 (
    .clock(line_1619_clock),
    .reset(line_1619_reset),
    .valid(line_1619_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1620)) line_1620 (
    .clock(line_1620_clock),
    .reset(line_1620_reset),
    .valid(line_1620_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1621)) line_1621 (
    .clock(line_1621_clock),
    .reset(line_1621_reset),
    .valid(line_1621_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1622)) line_1622 (
    .clock(line_1622_clock),
    .reset(line_1622_reset),
    .valid(line_1622_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1623)) line_1623 (
    .clock(line_1623_clock),
    .reset(line_1623_reset),
    .valid(line_1623_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1624)) line_1624 (
    .clock(line_1624_clock),
    .reset(line_1624_reset),
    .valid(line_1624_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1625)) line_1625 (
    .clock(line_1625_clock),
    .reset(line_1625_reset),
    .valid(line_1625_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1626)) line_1626 (
    .clock(line_1626_clock),
    .reset(line_1626_reset),
    .valid(line_1626_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1627)) line_1627 (
    .clock(line_1627_clock),
    .reset(line_1627_reset),
    .valid(line_1627_valid)
  );
  assign line_727_clock = clock;
  assign line_727_reset = reset;
  assign line_727_valid = wen ^ line_727_valid_reg;
  assign line_728_clock = clock;
  assign line_728_reset = reset;
  assign line_728_valid = enqueueFire_0 ^ line_728_valid_reg;
  assign line_729_clock = clock;
  assign line_729_reset = reset;
  assign line_729_valid = 2'h0 == _T_1[1:0] ^ line_729_valid_reg;
  assign line_730_clock = clock;
  assign line_730_reset = reset;
  assign line_730_valid = 2'h1 == _T_1[1:0] ^ line_730_valid_reg;
  assign line_731_clock = clock;
  assign line_731_reset = reset;
  assign line_731_valid = 2'h2 == _T_1[1:0] ^ line_731_valid_reg;
  assign line_732_clock = clock;
  assign line_732_reset = reset;
  assign line_732_valid = 2'h3 == _T_1[1:0] ^ line_732_valid_reg;
  assign line_733_clock = clock;
  assign line_733_reset = reset;
  assign line_733_valid = 2'h0 == _T_1[1:0] ^ line_733_valid_reg;
  assign line_734_clock = clock;
  assign line_734_reset = reset;
  assign line_734_valid = 2'h1 == _T_1[1:0] ^ line_734_valid_reg;
  assign line_735_clock = clock;
  assign line_735_reset = reset;
  assign line_735_valid = 2'h2 == _T_1[1:0] ^ line_735_valid_reg;
  assign line_736_clock = clock;
  assign line_736_reset = reset;
  assign line_736_valid = 2'h3 == _T_1[1:0] ^ line_736_valid_reg;
  assign line_737_clock = clock;
  assign line_737_reset = reset;
  assign line_737_valid = 2'h0 == _T_1[1:0] ^ line_737_valid_reg;
  assign line_738_clock = clock;
  assign line_738_reset = reset;
  assign line_738_valid = 2'h1 == _T_1[1:0] ^ line_738_valid_reg;
  assign line_739_clock = clock;
  assign line_739_reset = reset;
  assign line_739_valid = 2'h2 == _T_1[1:0] ^ line_739_valid_reg;
  assign line_740_clock = clock;
  assign line_740_reset = reset;
  assign line_740_valid = 2'h3 == _T_1[1:0] ^ line_740_valid_reg;
  assign line_741_clock = clock;
  assign line_741_reset = reset;
  assign line_741_valid = 2'h0 == _T_1[1:0] ^ line_741_valid_reg;
  assign line_742_clock = clock;
  assign line_742_reset = reset;
  assign line_742_valid = 2'h1 == _T_1[1:0] ^ line_742_valid_reg;
  assign line_743_clock = clock;
  assign line_743_reset = reset;
  assign line_743_valid = 2'h2 == _T_1[1:0] ^ line_743_valid_reg;
  assign line_744_clock = clock;
  assign line_744_reset = reset;
  assign line_744_valid = 2'h3 == _T_1[1:0] ^ line_744_valid_reg;
  assign line_745_clock = clock;
  assign line_745_reset = reset;
  assign line_745_valid = 2'h0 == _T_1[1:0] ^ line_745_valid_reg;
  assign line_746_clock = clock;
  assign line_746_reset = reset;
  assign line_746_valid = 2'h1 == _T_1[1:0] ^ line_746_valid_reg;
  assign line_747_clock = clock;
  assign line_747_reset = reset;
  assign line_747_valid = 2'h2 == _T_1[1:0] ^ line_747_valid_reg;
  assign line_748_clock = clock;
  assign line_748_reset = reset;
  assign line_748_valid = 2'h3 == _T_1[1:0] ^ line_748_valid_reg;
  assign line_749_clock = clock;
  assign line_749_reset = reset;
  assign line_749_valid = 2'h0 == _T_1[1:0] ^ line_749_valid_reg;
  assign line_750_clock = clock;
  assign line_750_reset = reset;
  assign line_750_valid = 2'h1 == _T_1[1:0] ^ line_750_valid_reg;
  assign line_751_clock = clock;
  assign line_751_reset = reset;
  assign line_751_valid = 2'h2 == _T_1[1:0] ^ line_751_valid_reg;
  assign line_752_clock = clock;
  assign line_752_reset = reset;
  assign line_752_valid = 2'h3 == _T_1[1:0] ^ line_752_valid_reg;
  assign line_753_clock = clock;
  assign line_753_reset = reset;
  assign line_753_valid = 2'h0 == _T_1[1:0] ^ line_753_valid_reg;
  assign line_754_clock = clock;
  assign line_754_reset = reset;
  assign line_754_valid = 2'h1 == _T_1[1:0] ^ line_754_valid_reg;
  assign line_755_clock = clock;
  assign line_755_reset = reset;
  assign line_755_valid = 2'h2 == _T_1[1:0] ^ line_755_valid_reg;
  assign line_756_clock = clock;
  assign line_756_reset = reset;
  assign line_756_valid = 2'h3 == _T_1[1:0] ^ line_756_valid_reg;
  assign line_757_clock = clock;
  assign line_757_reset = reset;
  assign line_757_valid = 2'h0 == _T_1[1:0] ^ line_757_valid_reg;
  assign line_758_clock = clock;
  assign line_758_reset = reset;
  assign line_758_valid = 2'h1 == _T_1[1:0] ^ line_758_valid_reg;
  assign line_759_clock = clock;
  assign line_759_reset = reset;
  assign line_759_valid = 2'h2 == _T_1[1:0] ^ line_759_valid_reg;
  assign line_760_clock = clock;
  assign line_760_reset = reset;
  assign line_760_valid = 2'h3 == _T_1[1:0] ^ line_760_valid_reg;
  assign line_761_clock = clock;
  assign line_761_reset = reset;
  assign line_761_valid = 2'h0 == _T_1[1:0] ^ line_761_valid_reg;
  assign line_762_clock = clock;
  assign line_762_reset = reset;
  assign line_762_valid = 2'h1 == _T_1[1:0] ^ line_762_valid_reg;
  assign line_763_clock = clock;
  assign line_763_reset = reset;
  assign line_763_valid = 2'h2 == _T_1[1:0] ^ line_763_valid_reg;
  assign line_764_clock = clock;
  assign line_764_reset = reset;
  assign line_764_valid = 2'h3 == _T_1[1:0] ^ line_764_valid_reg;
  assign line_765_clock = clock;
  assign line_765_reset = reset;
  assign line_765_valid = 2'h0 == _T_1[1:0] ^ line_765_valid_reg;
  assign line_766_clock = clock;
  assign line_766_reset = reset;
  assign line_766_valid = 2'h1 == _T_1[1:0] ^ line_766_valid_reg;
  assign line_767_clock = clock;
  assign line_767_reset = reset;
  assign line_767_valid = 2'h2 == _T_1[1:0] ^ line_767_valid_reg;
  assign line_768_clock = clock;
  assign line_768_reset = reset;
  assign line_768_valid = 2'h3 == _T_1[1:0] ^ line_768_valid_reg;
  assign line_769_clock = clock;
  assign line_769_reset = reset;
  assign line_769_valid = 2'h0 == _T_1[1:0] ^ line_769_valid_reg;
  assign line_770_clock = clock;
  assign line_770_reset = reset;
  assign line_770_valid = 2'h1 == _T_1[1:0] ^ line_770_valid_reg;
  assign line_771_clock = clock;
  assign line_771_reset = reset;
  assign line_771_valid = 2'h2 == _T_1[1:0] ^ line_771_valid_reg;
  assign line_772_clock = clock;
  assign line_772_reset = reset;
  assign line_772_valid = 2'h3 == _T_1[1:0] ^ line_772_valid_reg;
  assign line_773_clock = clock;
  assign line_773_reset = reset;
  assign line_773_valid = 2'h0 == _T_1[1:0] ^ line_773_valid_reg;
  assign line_774_clock = clock;
  assign line_774_reset = reset;
  assign line_774_valid = 2'h1 == _T_1[1:0] ^ line_774_valid_reg;
  assign line_775_clock = clock;
  assign line_775_reset = reset;
  assign line_775_valid = 2'h2 == _T_1[1:0] ^ line_775_valid_reg;
  assign line_776_clock = clock;
  assign line_776_reset = reset;
  assign line_776_valid = 2'h3 == _T_1[1:0] ^ line_776_valid_reg;
  assign line_777_clock = clock;
  assign line_777_reset = reset;
  assign line_777_valid = 2'h0 == _T_1[1:0] ^ line_777_valid_reg;
  assign line_778_clock = clock;
  assign line_778_reset = reset;
  assign line_778_valid = 2'h1 == _T_1[1:0] ^ line_778_valid_reg;
  assign line_779_clock = clock;
  assign line_779_reset = reset;
  assign line_779_valid = 2'h2 == _T_1[1:0] ^ line_779_valid_reg;
  assign line_780_clock = clock;
  assign line_780_reset = reset;
  assign line_780_valid = 2'h3 == _T_1[1:0] ^ line_780_valid_reg;
  assign line_781_clock = clock;
  assign line_781_reset = reset;
  assign line_781_valid = 2'h0 == _T_1[1:0] ^ line_781_valid_reg;
  assign line_782_clock = clock;
  assign line_782_reset = reset;
  assign line_782_valid = 2'h1 == _T_1[1:0] ^ line_782_valid_reg;
  assign line_783_clock = clock;
  assign line_783_reset = reset;
  assign line_783_valid = 2'h2 == _T_1[1:0] ^ line_783_valid_reg;
  assign line_784_clock = clock;
  assign line_784_reset = reset;
  assign line_784_valid = 2'h3 == _T_1[1:0] ^ line_784_valid_reg;
  assign line_785_clock = clock;
  assign line_785_reset = reset;
  assign line_785_valid = 2'h0 == _T_1[1:0] ^ line_785_valid_reg;
  assign line_786_clock = clock;
  assign line_786_reset = reset;
  assign line_786_valid = 2'h1 == _T_1[1:0] ^ line_786_valid_reg;
  assign line_787_clock = clock;
  assign line_787_reset = reset;
  assign line_787_valid = 2'h2 == _T_1[1:0] ^ line_787_valid_reg;
  assign line_788_clock = clock;
  assign line_788_reset = reset;
  assign line_788_valid = 2'h3 == _T_1[1:0] ^ line_788_valid_reg;
  assign line_789_clock = clock;
  assign line_789_reset = reset;
  assign line_789_valid = 2'h0 == _T_1[1:0] ^ line_789_valid_reg;
  assign line_790_clock = clock;
  assign line_790_reset = reset;
  assign line_790_valid = 2'h1 == _T_1[1:0] ^ line_790_valid_reg;
  assign line_791_clock = clock;
  assign line_791_reset = reset;
  assign line_791_valid = 2'h2 == _T_1[1:0] ^ line_791_valid_reg;
  assign line_792_clock = clock;
  assign line_792_reset = reset;
  assign line_792_valid = 2'h3 == _T_1[1:0] ^ line_792_valid_reg;
  assign line_793_clock = clock;
  assign line_793_reset = reset;
  assign line_793_valid = 2'h0 == _T_1[1:0] ^ line_793_valid_reg;
  assign line_794_clock = clock;
  assign line_794_reset = reset;
  assign line_794_valid = 2'h1 == _T_1[1:0] ^ line_794_valid_reg;
  assign line_795_clock = clock;
  assign line_795_reset = reset;
  assign line_795_valid = 2'h2 == _T_1[1:0] ^ line_795_valid_reg;
  assign line_796_clock = clock;
  assign line_796_reset = reset;
  assign line_796_valid = 2'h3 == _T_1[1:0] ^ line_796_valid_reg;
  assign line_797_clock = clock;
  assign line_797_reset = reset;
  assign line_797_valid = 2'h0 == _T_1[1:0] ^ line_797_valid_reg;
  assign line_798_clock = clock;
  assign line_798_reset = reset;
  assign line_798_valid = 2'h1 == _T_1[1:0] ^ line_798_valid_reg;
  assign line_799_clock = clock;
  assign line_799_reset = reset;
  assign line_799_valid = 2'h2 == _T_1[1:0] ^ line_799_valid_reg;
  assign line_800_clock = clock;
  assign line_800_reset = reset;
  assign line_800_valid = 2'h3 == _T_1[1:0] ^ line_800_valid_reg;
  assign line_801_clock = clock;
  assign line_801_reset = reset;
  assign line_801_valid = 2'h0 == _T_1[1:0] ^ line_801_valid_reg;
  assign line_802_clock = clock;
  assign line_802_reset = reset;
  assign line_802_valid = 2'h1 == _T_1[1:0] ^ line_802_valid_reg;
  assign line_803_clock = clock;
  assign line_803_reset = reset;
  assign line_803_valid = 2'h2 == _T_1[1:0] ^ line_803_valid_reg;
  assign line_804_clock = clock;
  assign line_804_reset = reset;
  assign line_804_valid = 2'h3 == _T_1[1:0] ^ line_804_valid_reg;
  assign line_805_clock = clock;
  assign line_805_reset = reset;
  assign line_805_valid = 2'h0 == _T_1[1:0] ^ line_805_valid_reg;
  assign line_806_clock = clock;
  assign line_806_reset = reset;
  assign line_806_valid = 2'h1 == _T_1[1:0] ^ line_806_valid_reg;
  assign line_807_clock = clock;
  assign line_807_reset = reset;
  assign line_807_valid = 2'h2 == _T_1[1:0] ^ line_807_valid_reg;
  assign line_808_clock = clock;
  assign line_808_reset = reset;
  assign line_808_valid = 2'h3 == _T_1[1:0] ^ line_808_valid_reg;
  assign line_809_clock = clock;
  assign line_809_reset = reset;
  assign line_809_valid = 2'h0 == _T_1[1:0] ^ line_809_valid_reg;
  assign line_810_clock = clock;
  assign line_810_reset = reset;
  assign line_810_valid = 2'h1 == _T_1[1:0] ^ line_810_valid_reg;
  assign line_811_clock = clock;
  assign line_811_reset = reset;
  assign line_811_valid = 2'h2 == _T_1[1:0] ^ line_811_valid_reg;
  assign line_812_clock = clock;
  assign line_812_reset = reset;
  assign line_812_valid = 2'h3 == _T_1[1:0] ^ line_812_valid_reg;
  assign line_813_clock = clock;
  assign line_813_reset = reset;
  assign line_813_valid = 2'h0 == _T_1[1:0] ^ line_813_valid_reg;
  assign line_814_clock = clock;
  assign line_814_reset = reset;
  assign line_814_valid = 2'h1 == _T_1[1:0] ^ line_814_valid_reg;
  assign line_815_clock = clock;
  assign line_815_reset = reset;
  assign line_815_valid = 2'h2 == _T_1[1:0] ^ line_815_valid_reg;
  assign line_816_clock = clock;
  assign line_816_reset = reset;
  assign line_816_valid = 2'h3 == _T_1[1:0] ^ line_816_valid_reg;
  assign line_817_clock = clock;
  assign line_817_reset = reset;
  assign line_817_valid = 2'h0 == _T_1[1:0] ^ line_817_valid_reg;
  assign line_818_clock = clock;
  assign line_818_reset = reset;
  assign line_818_valid = 2'h1 == _T_1[1:0] ^ line_818_valid_reg;
  assign line_819_clock = clock;
  assign line_819_reset = reset;
  assign line_819_valid = 2'h2 == _T_1[1:0] ^ line_819_valid_reg;
  assign line_820_clock = clock;
  assign line_820_reset = reset;
  assign line_820_valid = 2'h3 == _T_1[1:0] ^ line_820_valid_reg;
  assign line_821_clock = clock;
  assign line_821_reset = reset;
  assign line_821_valid = 2'h0 == _T_1[1:0] ^ line_821_valid_reg;
  assign line_822_clock = clock;
  assign line_822_reset = reset;
  assign line_822_valid = 2'h1 == _T_1[1:0] ^ line_822_valid_reg;
  assign line_823_clock = clock;
  assign line_823_reset = reset;
  assign line_823_valid = 2'h2 == _T_1[1:0] ^ line_823_valid_reg;
  assign line_824_clock = clock;
  assign line_824_reset = reset;
  assign line_824_valid = 2'h3 == _T_1[1:0] ^ line_824_valid_reg;
  assign line_825_clock = clock;
  assign line_825_reset = reset;
  assign line_825_valid = 2'h0 == _T_1[1:0] ^ line_825_valid_reg;
  assign line_826_clock = clock;
  assign line_826_reset = reset;
  assign line_826_valid = 2'h1 == _T_1[1:0] ^ line_826_valid_reg;
  assign line_827_clock = clock;
  assign line_827_reset = reset;
  assign line_827_valid = 2'h2 == _T_1[1:0] ^ line_827_valid_reg;
  assign line_828_clock = clock;
  assign line_828_reset = reset;
  assign line_828_valid = 2'h3 == _T_1[1:0] ^ line_828_valid_reg;
  assign line_829_clock = clock;
  assign line_829_reset = reset;
  assign line_829_valid = 2'h0 == _T_1[1:0] ^ line_829_valid_reg;
  assign line_830_clock = clock;
  assign line_830_reset = reset;
  assign line_830_valid = 2'h1 == _T_1[1:0] ^ line_830_valid_reg;
  assign line_831_clock = clock;
  assign line_831_reset = reset;
  assign line_831_valid = 2'h2 == _T_1[1:0] ^ line_831_valid_reg;
  assign line_832_clock = clock;
  assign line_832_reset = reset;
  assign line_832_valid = 2'h3 == _T_1[1:0] ^ line_832_valid_reg;
  assign line_833_clock = clock;
  assign line_833_reset = reset;
  assign line_833_valid = 2'h0 == _T_1[1:0] ^ line_833_valid_reg;
  assign line_834_clock = clock;
  assign line_834_reset = reset;
  assign line_834_valid = 2'h1 == _T_1[1:0] ^ line_834_valid_reg;
  assign line_835_clock = clock;
  assign line_835_reset = reset;
  assign line_835_valid = 2'h2 == _T_1[1:0] ^ line_835_valid_reg;
  assign line_836_clock = clock;
  assign line_836_reset = reset;
  assign line_836_valid = 2'h3 == _T_1[1:0] ^ line_836_valid_reg;
  assign line_837_clock = clock;
  assign line_837_reset = reset;
  assign line_837_valid = 2'h0 == _T_1[1:0] ^ line_837_valid_reg;
  assign line_838_clock = clock;
  assign line_838_reset = reset;
  assign line_838_valid = 2'h1 == _T_1[1:0] ^ line_838_valid_reg;
  assign line_839_clock = clock;
  assign line_839_reset = reset;
  assign line_839_valid = 2'h2 == _T_1[1:0] ^ line_839_valid_reg;
  assign line_840_clock = clock;
  assign line_840_reset = reset;
  assign line_840_valid = 2'h3 == _T_1[1:0] ^ line_840_valid_reg;
  assign line_841_clock = clock;
  assign line_841_reset = reset;
  assign line_841_valid = 2'h0 == _T_1[1:0] ^ line_841_valid_reg;
  assign line_842_clock = clock;
  assign line_842_reset = reset;
  assign line_842_valid = 2'h1 == _T_1[1:0] ^ line_842_valid_reg;
  assign line_843_clock = clock;
  assign line_843_reset = reset;
  assign line_843_valid = 2'h2 == _T_1[1:0] ^ line_843_valid_reg;
  assign line_844_clock = clock;
  assign line_844_reset = reset;
  assign line_844_valid = 2'h3 == _T_1[1:0] ^ line_844_valid_reg;
  assign line_845_clock = clock;
  assign line_845_reset = reset;
  assign line_845_valid = 2'h0 == _T_1[1:0] ^ line_845_valid_reg;
  assign line_846_clock = clock;
  assign line_846_reset = reset;
  assign line_846_valid = 2'h1 == _T_1[1:0] ^ line_846_valid_reg;
  assign line_847_clock = clock;
  assign line_847_reset = reset;
  assign line_847_valid = 2'h2 == _T_1[1:0] ^ line_847_valid_reg;
  assign line_848_clock = clock;
  assign line_848_reset = reset;
  assign line_848_valid = 2'h3 == _T_1[1:0] ^ line_848_valid_reg;
  assign line_849_clock = clock;
  assign line_849_reset = reset;
  assign line_849_valid = 2'h0 == _T_1[1:0] ^ line_849_valid_reg;
  assign line_850_clock = clock;
  assign line_850_reset = reset;
  assign line_850_valid = 2'h1 == _T_1[1:0] ^ line_850_valid_reg;
  assign line_851_clock = clock;
  assign line_851_reset = reset;
  assign line_851_valid = 2'h2 == _T_1[1:0] ^ line_851_valid_reg;
  assign line_852_clock = clock;
  assign line_852_reset = reset;
  assign line_852_valid = 2'h3 == _T_1[1:0] ^ line_852_valid_reg;
  assign line_853_clock = clock;
  assign line_853_reset = reset;
  assign line_853_valid = 2'h0 == _T_1[1:0] ^ line_853_valid_reg;
  assign line_854_clock = clock;
  assign line_854_reset = reset;
  assign line_854_valid = 2'h1 == _T_1[1:0] ^ line_854_valid_reg;
  assign line_855_clock = clock;
  assign line_855_reset = reset;
  assign line_855_valid = 2'h2 == _T_1[1:0] ^ line_855_valid_reg;
  assign line_856_clock = clock;
  assign line_856_reset = reset;
  assign line_856_valid = 2'h3 == _T_1[1:0] ^ line_856_valid_reg;
  assign line_857_clock = clock;
  assign line_857_reset = reset;
  assign line_857_valid = 2'h0 == _T_1[1:0] ^ line_857_valid_reg;
  assign line_858_clock = clock;
  assign line_858_reset = reset;
  assign line_858_valid = 2'h1 == _T_1[1:0] ^ line_858_valid_reg;
  assign line_859_clock = clock;
  assign line_859_reset = reset;
  assign line_859_valid = 2'h2 == _T_1[1:0] ^ line_859_valid_reg;
  assign line_860_clock = clock;
  assign line_860_reset = reset;
  assign line_860_valid = 2'h3 == _T_1[1:0] ^ line_860_valid_reg;
  assign line_861_clock = clock;
  assign line_861_reset = reset;
  assign line_861_valid = 2'h0 == _T_1[1:0] ^ line_861_valid_reg;
  assign line_862_clock = clock;
  assign line_862_reset = reset;
  assign line_862_valid = 2'h1 == _T_1[1:0] ^ line_862_valid_reg;
  assign line_863_clock = clock;
  assign line_863_reset = reset;
  assign line_863_valid = 2'h2 == _T_1[1:0] ^ line_863_valid_reg;
  assign line_864_clock = clock;
  assign line_864_reset = reset;
  assign line_864_valid = 2'h3 == _T_1[1:0] ^ line_864_valid_reg;
  assign line_865_clock = clock;
  assign line_865_reset = reset;
  assign line_865_valid = 2'h0 == _T_1[1:0] ^ line_865_valid_reg;
  assign line_866_clock = clock;
  assign line_866_reset = reset;
  assign line_866_valid = 2'h1 == _T_1[1:0] ^ line_866_valid_reg;
  assign line_867_clock = clock;
  assign line_867_reset = reset;
  assign line_867_valid = 2'h2 == _T_1[1:0] ^ line_867_valid_reg;
  assign line_868_clock = clock;
  assign line_868_reset = reset;
  assign line_868_valid = 2'h3 == _T_1[1:0] ^ line_868_valid_reg;
  assign line_869_clock = clock;
  assign line_869_reset = reset;
  assign line_869_valid = 2'h0 == _T_1[1:0] ^ line_869_valid_reg;
  assign line_870_clock = clock;
  assign line_870_reset = reset;
  assign line_870_valid = 2'h1 == _T_1[1:0] ^ line_870_valid_reg;
  assign line_871_clock = clock;
  assign line_871_reset = reset;
  assign line_871_valid = 2'h2 == _T_1[1:0] ^ line_871_valid_reg;
  assign line_872_clock = clock;
  assign line_872_reset = reset;
  assign line_872_valid = 2'h3 == _T_1[1:0] ^ line_872_valid_reg;
  assign line_873_clock = clock;
  assign line_873_reset = reset;
  assign line_873_valid = 2'h0 == _T_1[1:0] ^ line_873_valid_reg;
  assign line_874_clock = clock;
  assign line_874_reset = reset;
  assign line_874_valid = 2'h1 == _T_1[1:0] ^ line_874_valid_reg;
  assign line_875_clock = clock;
  assign line_875_reset = reset;
  assign line_875_valid = 2'h2 == _T_1[1:0] ^ line_875_valid_reg;
  assign line_876_clock = clock;
  assign line_876_reset = reset;
  assign line_876_valid = 2'h3 == _T_1[1:0] ^ line_876_valid_reg;
  assign line_877_clock = clock;
  assign line_877_reset = reset;
  assign line_877_valid = 2'h0 == _T_1[1:0] ^ line_877_valid_reg;
  assign line_878_clock = clock;
  assign line_878_reset = reset;
  assign line_878_valid = 2'h1 == _T_1[1:0] ^ line_878_valid_reg;
  assign line_879_clock = clock;
  assign line_879_reset = reset;
  assign line_879_valid = 2'h2 == _T_1[1:0] ^ line_879_valid_reg;
  assign line_880_clock = clock;
  assign line_880_reset = reset;
  assign line_880_valid = 2'h3 == _T_1[1:0] ^ line_880_valid_reg;
  assign line_881_clock = clock;
  assign line_881_reset = reset;
  assign line_881_valid = 2'h0 == _T_1[1:0] ^ line_881_valid_reg;
  assign line_882_clock = clock;
  assign line_882_reset = reset;
  assign line_882_valid = 2'h1 == _T_1[1:0] ^ line_882_valid_reg;
  assign line_883_clock = clock;
  assign line_883_reset = reset;
  assign line_883_valid = 2'h2 == _T_1[1:0] ^ line_883_valid_reg;
  assign line_884_clock = clock;
  assign line_884_reset = reset;
  assign line_884_valid = 2'h3 == _T_1[1:0] ^ line_884_valid_reg;
  assign line_885_clock = clock;
  assign line_885_reset = reset;
  assign line_885_valid = 2'h0 == _T_1[1:0] ^ line_885_valid_reg;
  assign line_886_clock = clock;
  assign line_886_reset = reset;
  assign line_886_valid = 2'h1 == _T_1[1:0] ^ line_886_valid_reg;
  assign line_887_clock = clock;
  assign line_887_reset = reset;
  assign line_887_valid = 2'h2 == _T_1[1:0] ^ line_887_valid_reg;
  assign line_888_clock = clock;
  assign line_888_reset = reset;
  assign line_888_valid = 2'h3 == _T_1[1:0] ^ line_888_valid_reg;
  assign line_889_clock = clock;
  assign line_889_reset = reset;
  assign line_889_valid = 2'h0 == _T_1[1:0] ^ line_889_valid_reg;
  assign line_890_clock = clock;
  assign line_890_reset = reset;
  assign line_890_valid = 2'h1 == _T_1[1:0] ^ line_890_valid_reg;
  assign line_891_clock = clock;
  assign line_891_reset = reset;
  assign line_891_valid = 2'h2 == _T_1[1:0] ^ line_891_valid_reg;
  assign line_892_clock = clock;
  assign line_892_reset = reset;
  assign line_892_valid = 2'h3 == _T_1[1:0] ^ line_892_valid_reg;
  assign line_893_clock = clock;
  assign line_893_reset = reset;
  assign line_893_valid = 2'h0 == _T_1[1:0] ^ line_893_valid_reg;
  assign line_894_clock = clock;
  assign line_894_reset = reset;
  assign line_894_valid = 2'h1 == _T_1[1:0] ^ line_894_valid_reg;
  assign line_895_clock = clock;
  assign line_895_reset = reset;
  assign line_895_valid = 2'h2 == _T_1[1:0] ^ line_895_valid_reg;
  assign line_896_clock = clock;
  assign line_896_reset = reset;
  assign line_896_valid = 2'h3 == _T_1[1:0] ^ line_896_valid_reg;
  assign line_897_clock = clock;
  assign line_897_reset = reset;
  assign line_897_valid = 2'h0 == _T_1[1:0] ^ line_897_valid_reg;
  assign line_898_clock = clock;
  assign line_898_reset = reset;
  assign line_898_valid = 2'h1 == _T_1[1:0] ^ line_898_valid_reg;
  assign line_899_clock = clock;
  assign line_899_reset = reset;
  assign line_899_valid = 2'h2 == _T_1[1:0] ^ line_899_valid_reg;
  assign line_900_clock = clock;
  assign line_900_reset = reset;
  assign line_900_valid = 2'h3 == _T_1[1:0] ^ line_900_valid_reg;
  assign line_901_clock = clock;
  assign line_901_reset = reset;
  assign line_901_valid = 2'h0 == _T_1[1:0] ^ line_901_valid_reg;
  assign line_902_clock = clock;
  assign line_902_reset = reset;
  assign line_902_valid = 2'h1 == _T_1[1:0] ^ line_902_valid_reg;
  assign line_903_clock = clock;
  assign line_903_reset = reset;
  assign line_903_valid = 2'h2 == _T_1[1:0] ^ line_903_valid_reg;
  assign line_904_clock = clock;
  assign line_904_reset = reset;
  assign line_904_valid = 2'h3 == _T_1[1:0] ^ line_904_valid_reg;
  assign line_905_clock = clock;
  assign line_905_reset = reset;
  assign line_905_valid = 2'h0 == _T_1[1:0] ^ line_905_valid_reg;
  assign line_906_clock = clock;
  assign line_906_reset = reset;
  assign line_906_valid = 2'h1 == _T_1[1:0] ^ line_906_valid_reg;
  assign line_907_clock = clock;
  assign line_907_reset = reset;
  assign line_907_valid = 2'h2 == _T_1[1:0] ^ line_907_valid_reg;
  assign line_908_clock = clock;
  assign line_908_reset = reset;
  assign line_908_valid = 2'h3 == _T_1[1:0] ^ line_908_valid_reg;
  assign line_909_clock = clock;
  assign line_909_reset = reset;
  assign line_909_valid = 2'h0 == _T_1[1:0] ^ line_909_valid_reg;
  assign line_910_clock = clock;
  assign line_910_reset = reset;
  assign line_910_valid = 2'h1 == _T_1[1:0] ^ line_910_valid_reg;
  assign line_911_clock = clock;
  assign line_911_reset = reset;
  assign line_911_valid = 2'h2 == _T_1[1:0] ^ line_911_valid_reg;
  assign line_912_clock = clock;
  assign line_912_reset = reset;
  assign line_912_valid = 2'h3 == _T_1[1:0] ^ line_912_valid_reg;
  assign line_913_clock = clock;
  assign line_913_reset = reset;
  assign line_913_valid = 2'h0 == _T_1[1:0] ^ line_913_valid_reg;
  assign line_914_clock = clock;
  assign line_914_reset = reset;
  assign line_914_valid = 2'h1 == _T_1[1:0] ^ line_914_valid_reg;
  assign line_915_clock = clock;
  assign line_915_reset = reset;
  assign line_915_valid = 2'h2 == _T_1[1:0] ^ line_915_valid_reg;
  assign line_916_clock = clock;
  assign line_916_reset = reset;
  assign line_916_valid = 2'h3 == _T_1[1:0] ^ line_916_valid_reg;
  assign line_917_clock = clock;
  assign line_917_reset = reset;
  assign line_917_valid = 2'h0 == _T_1[1:0] ^ line_917_valid_reg;
  assign line_918_clock = clock;
  assign line_918_reset = reset;
  assign line_918_valid = 2'h1 == _T_1[1:0] ^ line_918_valid_reg;
  assign line_919_clock = clock;
  assign line_919_reset = reset;
  assign line_919_valid = 2'h2 == _T_1[1:0] ^ line_919_valid_reg;
  assign line_920_clock = clock;
  assign line_920_reset = reset;
  assign line_920_valid = 2'h3 == _T_1[1:0] ^ line_920_valid_reg;
  assign line_921_clock = clock;
  assign line_921_reset = reset;
  assign line_921_valid = 2'h0 == _T_1[1:0] ^ line_921_valid_reg;
  assign line_922_clock = clock;
  assign line_922_reset = reset;
  assign line_922_valid = 2'h1 == _T_1[1:0] ^ line_922_valid_reg;
  assign line_923_clock = clock;
  assign line_923_reset = reset;
  assign line_923_valid = 2'h2 == _T_1[1:0] ^ line_923_valid_reg;
  assign line_924_clock = clock;
  assign line_924_reset = reset;
  assign line_924_valid = 2'h3 == _T_1[1:0] ^ line_924_valid_reg;
  assign line_925_clock = clock;
  assign line_925_reset = reset;
  assign line_925_valid = 2'h0 == _T_1[1:0] ^ line_925_valid_reg;
  assign line_926_clock = clock;
  assign line_926_reset = reset;
  assign line_926_valid = 2'h1 == _T_1[1:0] ^ line_926_valid_reg;
  assign line_927_clock = clock;
  assign line_927_reset = reset;
  assign line_927_valid = 2'h2 == _T_1[1:0] ^ line_927_valid_reg;
  assign line_928_clock = clock;
  assign line_928_reset = reset;
  assign line_928_valid = 2'h3 == _T_1[1:0] ^ line_928_valid_reg;
  assign line_929_clock = clock;
  assign line_929_reset = reset;
  assign line_929_valid = 2'h0 == _T_1[1:0] ^ line_929_valid_reg;
  assign line_930_clock = clock;
  assign line_930_reset = reset;
  assign line_930_valid = 2'h1 == _T_1[1:0] ^ line_930_valid_reg;
  assign line_931_clock = clock;
  assign line_931_reset = reset;
  assign line_931_valid = 2'h2 == _T_1[1:0] ^ line_931_valid_reg;
  assign line_932_clock = clock;
  assign line_932_reset = reset;
  assign line_932_valid = 2'h3 == _T_1[1:0] ^ line_932_valid_reg;
  assign line_933_clock = clock;
  assign line_933_reset = reset;
  assign line_933_valid = 2'h0 == _T_1[1:0] ^ line_933_valid_reg;
  assign line_934_clock = clock;
  assign line_934_reset = reset;
  assign line_934_valid = 2'h1 == _T_1[1:0] ^ line_934_valid_reg;
  assign line_935_clock = clock;
  assign line_935_reset = reset;
  assign line_935_valid = 2'h2 == _T_1[1:0] ^ line_935_valid_reg;
  assign line_936_clock = clock;
  assign line_936_reset = reset;
  assign line_936_valid = 2'h3 == _T_1[1:0] ^ line_936_valid_reg;
  assign line_937_clock = clock;
  assign line_937_reset = reset;
  assign line_937_valid = 2'h0 == _T_1[1:0] ^ line_937_valid_reg;
  assign line_938_clock = clock;
  assign line_938_reset = reset;
  assign line_938_valid = 2'h1 == _T_1[1:0] ^ line_938_valid_reg;
  assign line_939_clock = clock;
  assign line_939_reset = reset;
  assign line_939_valid = 2'h2 == _T_1[1:0] ^ line_939_valid_reg;
  assign line_940_clock = clock;
  assign line_940_reset = reset;
  assign line_940_valid = 2'h3 == _T_1[1:0] ^ line_940_valid_reg;
  assign line_941_clock = clock;
  assign line_941_reset = reset;
  assign line_941_valid = 2'h0 == _T_1[1:0] ^ line_941_valid_reg;
  assign line_942_clock = clock;
  assign line_942_reset = reset;
  assign line_942_valid = 2'h1 == _T_1[1:0] ^ line_942_valid_reg;
  assign line_943_clock = clock;
  assign line_943_reset = reset;
  assign line_943_valid = 2'h2 == _T_1[1:0] ^ line_943_valid_reg;
  assign line_944_clock = clock;
  assign line_944_reset = reset;
  assign line_944_valid = 2'h3 == _T_1[1:0] ^ line_944_valid_reg;
  assign line_945_clock = clock;
  assign line_945_reset = reset;
  assign line_945_valid = 2'h0 == _T_1[1:0] ^ line_945_valid_reg;
  assign line_946_clock = clock;
  assign line_946_reset = reset;
  assign line_946_valid = 2'h1 == _T_1[1:0] ^ line_946_valid_reg;
  assign line_947_clock = clock;
  assign line_947_reset = reset;
  assign line_947_valid = 2'h2 == _T_1[1:0] ^ line_947_valid_reg;
  assign line_948_clock = clock;
  assign line_948_reset = reset;
  assign line_948_valid = 2'h3 == _T_1[1:0] ^ line_948_valid_reg;
  assign line_949_clock = clock;
  assign line_949_reset = reset;
  assign line_949_valid = 2'h0 == _T_1[1:0] ^ line_949_valid_reg;
  assign line_950_clock = clock;
  assign line_950_reset = reset;
  assign line_950_valid = 2'h1 == _T_1[1:0] ^ line_950_valid_reg;
  assign line_951_clock = clock;
  assign line_951_reset = reset;
  assign line_951_valid = 2'h2 == _T_1[1:0] ^ line_951_valid_reg;
  assign line_952_clock = clock;
  assign line_952_reset = reset;
  assign line_952_valid = 2'h3 == _T_1[1:0] ^ line_952_valid_reg;
  assign line_953_clock = clock;
  assign line_953_reset = reset;
  assign line_953_valid = enqueueFire_1 ^ line_953_valid_reg;
  assign line_954_clock = clock;
  assign line_954_reset = reset;
  assign line_954_valid = 2'h0 == _T_4 ^ line_954_valid_reg;
  assign line_955_clock = clock;
  assign line_955_reset = reset;
  assign line_955_valid = 2'h1 == _T_4 ^ line_955_valid_reg;
  assign line_956_clock = clock;
  assign line_956_reset = reset;
  assign line_956_valid = 2'h2 == _T_4 ^ line_956_valid_reg;
  assign line_957_clock = clock;
  assign line_957_reset = reset;
  assign line_957_valid = 2'h3 == _T_4 ^ line_957_valid_reg;
  assign line_958_clock = clock;
  assign line_958_reset = reset;
  assign line_958_valid = 2'h0 == _T_4 ^ line_958_valid_reg;
  assign line_959_clock = clock;
  assign line_959_reset = reset;
  assign line_959_valid = 2'h1 == _T_4 ^ line_959_valid_reg;
  assign line_960_clock = clock;
  assign line_960_reset = reset;
  assign line_960_valid = 2'h2 == _T_4 ^ line_960_valid_reg;
  assign line_961_clock = clock;
  assign line_961_reset = reset;
  assign line_961_valid = 2'h3 == _T_4 ^ line_961_valid_reg;
  assign line_962_clock = clock;
  assign line_962_reset = reset;
  assign line_962_valid = 2'h0 == _T_4 ^ line_962_valid_reg;
  assign line_963_clock = clock;
  assign line_963_reset = reset;
  assign line_963_valid = 2'h1 == _T_4 ^ line_963_valid_reg;
  assign line_964_clock = clock;
  assign line_964_reset = reset;
  assign line_964_valid = 2'h2 == _T_4 ^ line_964_valid_reg;
  assign line_965_clock = clock;
  assign line_965_reset = reset;
  assign line_965_valid = 2'h3 == _T_4 ^ line_965_valid_reg;
  assign line_966_clock = clock;
  assign line_966_reset = reset;
  assign line_966_valid = 2'h0 == _T_4 ^ line_966_valid_reg;
  assign line_967_clock = clock;
  assign line_967_reset = reset;
  assign line_967_valid = 2'h1 == _T_4 ^ line_967_valid_reg;
  assign line_968_clock = clock;
  assign line_968_reset = reset;
  assign line_968_valid = 2'h2 == _T_4 ^ line_968_valid_reg;
  assign line_969_clock = clock;
  assign line_969_reset = reset;
  assign line_969_valid = 2'h3 == _T_4 ^ line_969_valid_reg;
  assign line_970_clock = clock;
  assign line_970_reset = reset;
  assign line_970_valid = 2'h0 == _T_4 ^ line_970_valid_reg;
  assign line_971_clock = clock;
  assign line_971_reset = reset;
  assign line_971_valid = 2'h1 == _T_4 ^ line_971_valid_reg;
  assign line_972_clock = clock;
  assign line_972_reset = reset;
  assign line_972_valid = 2'h2 == _T_4 ^ line_972_valid_reg;
  assign line_973_clock = clock;
  assign line_973_reset = reset;
  assign line_973_valid = 2'h3 == _T_4 ^ line_973_valid_reg;
  assign line_974_clock = clock;
  assign line_974_reset = reset;
  assign line_974_valid = 2'h0 == _T_4 ^ line_974_valid_reg;
  assign line_975_clock = clock;
  assign line_975_reset = reset;
  assign line_975_valid = 2'h1 == _T_4 ^ line_975_valid_reg;
  assign line_976_clock = clock;
  assign line_976_reset = reset;
  assign line_976_valid = 2'h2 == _T_4 ^ line_976_valid_reg;
  assign line_977_clock = clock;
  assign line_977_reset = reset;
  assign line_977_valid = 2'h3 == _T_4 ^ line_977_valid_reg;
  assign line_978_clock = clock;
  assign line_978_reset = reset;
  assign line_978_valid = 2'h0 == _T_4 ^ line_978_valid_reg;
  assign line_979_clock = clock;
  assign line_979_reset = reset;
  assign line_979_valid = 2'h1 == _T_4 ^ line_979_valid_reg;
  assign line_980_clock = clock;
  assign line_980_reset = reset;
  assign line_980_valid = 2'h2 == _T_4 ^ line_980_valid_reg;
  assign line_981_clock = clock;
  assign line_981_reset = reset;
  assign line_981_valid = 2'h3 == _T_4 ^ line_981_valid_reg;
  assign line_982_clock = clock;
  assign line_982_reset = reset;
  assign line_982_valid = 2'h0 == _T_4 ^ line_982_valid_reg;
  assign line_983_clock = clock;
  assign line_983_reset = reset;
  assign line_983_valid = 2'h1 == _T_4 ^ line_983_valid_reg;
  assign line_984_clock = clock;
  assign line_984_reset = reset;
  assign line_984_valid = 2'h2 == _T_4 ^ line_984_valid_reg;
  assign line_985_clock = clock;
  assign line_985_reset = reset;
  assign line_985_valid = 2'h3 == _T_4 ^ line_985_valid_reg;
  assign line_986_clock = clock;
  assign line_986_reset = reset;
  assign line_986_valid = 2'h0 == _T_4 ^ line_986_valid_reg;
  assign line_987_clock = clock;
  assign line_987_reset = reset;
  assign line_987_valid = 2'h1 == _T_4 ^ line_987_valid_reg;
  assign line_988_clock = clock;
  assign line_988_reset = reset;
  assign line_988_valid = 2'h2 == _T_4 ^ line_988_valid_reg;
  assign line_989_clock = clock;
  assign line_989_reset = reset;
  assign line_989_valid = 2'h3 == _T_4 ^ line_989_valid_reg;
  assign line_990_clock = clock;
  assign line_990_reset = reset;
  assign line_990_valid = 2'h0 == _T_4 ^ line_990_valid_reg;
  assign line_991_clock = clock;
  assign line_991_reset = reset;
  assign line_991_valid = 2'h1 == _T_4 ^ line_991_valid_reg;
  assign line_992_clock = clock;
  assign line_992_reset = reset;
  assign line_992_valid = 2'h2 == _T_4 ^ line_992_valid_reg;
  assign line_993_clock = clock;
  assign line_993_reset = reset;
  assign line_993_valid = 2'h3 == _T_4 ^ line_993_valid_reg;
  assign line_994_clock = clock;
  assign line_994_reset = reset;
  assign line_994_valid = 2'h0 == _T_4 ^ line_994_valid_reg;
  assign line_995_clock = clock;
  assign line_995_reset = reset;
  assign line_995_valid = 2'h1 == _T_4 ^ line_995_valid_reg;
  assign line_996_clock = clock;
  assign line_996_reset = reset;
  assign line_996_valid = 2'h2 == _T_4 ^ line_996_valid_reg;
  assign line_997_clock = clock;
  assign line_997_reset = reset;
  assign line_997_valid = 2'h3 == _T_4 ^ line_997_valid_reg;
  assign line_998_clock = clock;
  assign line_998_reset = reset;
  assign line_998_valid = 2'h0 == _T_4 ^ line_998_valid_reg;
  assign line_999_clock = clock;
  assign line_999_reset = reset;
  assign line_999_valid = 2'h1 == _T_4 ^ line_999_valid_reg;
  assign line_1000_clock = clock;
  assign line_1000_reset = reset;
  assign line_1000_valid = 2'h2 == _T_4 ^ line_1000_valid_reg;
  assign line_1001_clock = clock;
  assign line_1001_reset = reset;
  assign line_1001_valid = 2'h3 == _T_4 ^ line_1001_valid_reg;
  assign line_1002_clock = clock;
  assign line_1002_reset = reset;
  assign line_1002_valid = 2'h0 == _T_4 ^ line_1002_valid_reg;
  assign line_1003_clock = clock;
  assign line_1003_reset = reset;
  assign line_1003_valid = 2'h1 == _T_4 ^ line_1003_valid_reg;
  assign line_1004_clock = clock;
  assign line_1004_reset = reset;
  assign line_1004_valid = 2'h2 == _T_4 ^ line_1004_valid_reg;
  assign line_1005_clock = clock;
  assign line_1005_reset = reset;
  assign line_1005_valid = 2'h3 == _T_4 ^ line_1005_valid_reg;
  assign line_1006_clock = clock;
  assign line_1006_reset = reset;
  assign line_1006_valid = 2'h0 == _T_4 ^ line_1006_valid_reg;
  assign line_1007_clock = clock;
  assign line_1007_reset = reset;
  assign line_1007_valid = 2'h1 == _T_4 ^ line_1007_valid_reg;
  assign line_1008_clock = clock;
  assign line_1008_reset = reset;
  assign line_1008_valid = 2'h2 == _T_4 ^ line_1008_valid_reg;
  assign line_1009_clock = clock;
  assign line_1009_reset = reset;
  assign line_1009_valid = 2'h3 == _T_4 ^ line_1009_valid_reg;
  assign line_1010_clock = clock;
  assign line_1010_reset = reset;
  assign line_1010_valid = 2'h0 == _T_4 ^ line_1010_valid_reg;
  assign line_1011_clock = clock;
  assign line_1011_reset = reset;
  assign line_1011_valid = 2'h1 == _T_4 ^ line_1011_valid_reg;
  assign line_1012_clock = clock;
  assign line_1012_reset = reset;
  assign line_1012_valid = 2'h2 == _T_4 ^ line_1012_valid_reg;
  assign line_1013_clock = clock;
  assign line_1013_reset = reset;
  assign line_1013_valid = 2'h3 == _T_4 ^ line_1013_valid_reg;
  assign line_1014_clock = clock;
  assign line_1014_reset = reset;
  assign line_1014_valid = 2'h0 == _T_4 ^ line_1014_valid_reg;
  assign line_1015_clock = clock;
  assign line_1015_reset = reset;
  assign line_1015_valid = 2'h1 == _T_4 ^ line_1015_valid_reg;
  assign line_1016_clock = clock;
  assign line_1016_reset = reset;
  assign line_1016_valid = 2'h2 == _T_4 ^ line_1016_valid_reg;
  assign line_1017_clock = clock;
  assign line_1017_reset = reset;
  assign line_1017_valid = 2'h3 == _T_4 ^ line_1017_valid_reg;
  assign line_1018_clock = clock;
  assign line_1018_reset = reset;
  assign line_1018_valid = 2'h0 == _T_4 ^ line_1018_valid_reg;
  assign line_1019_clock = clock;
  assign line_1019_reset = reset;
  assign line_1019_valid = 2'h1 == _T_4 ^ line_1019_valid_reg;
  assign line_1020_clock = clock;
  assign line_1020_reset = reset;
  assign line_1020_valid = 2'h2 == _T_4 ^ line_1020_valid_reg;
  assign line_1021_clock = clock;
  assign line_1021_reset = reset;
  assign line_1021_valid = 2'h3 == _T_4 ^ line_1021_valid_reg;
  assign line_1022_clock = clock;
  assign line_1022_reset = reset;
  assign line_1022_valid = 2'h0 == _T_4 ^ line_1022_valid_reg;
  assign line_1023_clock = clock;
  assign line_1023_reset = reset;
  assign line_1023_valid = 2'h1 == _T_4 ^ line_1023_valid_reg;
  assign line_1024_clock = clock;
  assign line_1024_reset = reset;
  assign line_1024_valid = 2'h2 == _T_4 ^ line_1024_valid_reg;
  assign line_1025_clock = clock;
  assign line_1025_reset = reset;
  assign line_1025_valid = 2'h3 == _T_4 ^ line_1025_valid_reg;
  assign line_1026_clock = clock;
  assign line_1026_reset = reset;
  assign line_1026_valid = 2'h0 == _T_4 ^ line_1026_valid_reg;
  assign line_1027_clock = clock;
  assign line_1027_reset = reset;
  assign line_1027_valid = 2'h1 == _T_4 ^ line_1027_valid_reg;
  assign line_1028_clock = clock;
  assign line_1028_reset = reset;
  assign line_1028_valid = 2'h2 == _T_4 ^ line_1028_valid_reg;
  assign line_1029_clock = clock;
  assign line_1029_reset = reset;
  assign line_1029_valid = 2'h3 == _T_4 ^ line_1029_valid_reg;
  assign line_1030_clock = clock;
  assign line_1030_reset = reset;
  assign line_1030_valid = 2'h0 == _T_4 ^ line_1030_valid_reg;
  assign line_1031_clock = clock;
  assign line_1031_reset = reset;
  assign line_1031_valid = 2'h1 == _T_4 ^ line_1031_valid_reg;
  assign line_1032_clock = clock;
  assign line_1032_reset = reset;
  assign line_1032_valid = 2'h2 == _T_4 ^ line_1032_valid_reg;
  assign line_1033_clock = clock;
  assign line_1033_reset = reset;
  assign line_1033_valid = 2'h3 == _T_4 ^ line_1033_valid_reg;
  assign line_1034_clock = clock;
  assign line_1034_reset = reset;
  assign line_1034_valid = 2'h0 == _T_4 ^ line_1034_valid_reg;
  assign line_1035_clock = clock;
  assign line_1035_reset = reset;
  assign line_1035_valid = 2'h1 == _T_4 ^ line_1035_valid_reg;
  assign line_1036_clock = clock;
  assign line_1036_reset = reset;
  assign line_1036_valid = 2'h2 == _T_4 ^ line_1036_valid_reg;
  assign line_1037_clock = clock;
  assign line_1037_reset = reset;
  assign line_1037_valid = 2'h3 == _T_4 ^ line_1037_valid_reg;
  assign line_1038_clock = clock;
  assign line_1038_reset = reset;
  assign line_1038_valid = 2'h0 == _T_4 ^ line_1038_valid_reg;
  assign line_1039_clock = clock;
  assign line_1039_reset = reset;
  assign line_1039_valid = 2'h1 == _T_4 ^ line_1039_valid_reg;
  assign line_1040_clock = clock;
  assign line_1040_reset = reset;
  assign line_1040_valid = 2'h2 == _T_4 ^ line_1040_valid_reg;
  assign line_1041_clock = clock;
  assign line_1041_reset = reset;
  assign line_1041_valid = 2'h3 == _T_4 ^ line_1041_valid_reg;
  assign line_1042_clock = clock;
  assign line_1042_reset = reset;
  assign line_1042_valid = 2'h0 == _T_4 ^ line_1042_valid_reg;
  assign line_1043_clock = clock;
  assign line_1043_reset = reset;
  assign line_1043_valid = 2'h1 == _T_4 ^ line_1043_valid_reg;
  assign line_1044_clock = clock;
  assign line_1044_reset = reset;
  assign line_1044_valid = 2'h2 == _T_4 ^ line_1044_valid_reg;
  assign line_1045_clock = clock;
  assign line_1045_reset = reset;
  assign line_1045_valid = 2'h3 == _T_4 ^ line_1045_valid_reg;
  assign line_1046_clock = clock;
  assign line_1046_reset = reset;
  assign line_1046_valid = 2'h0 == _T_4 ^ line_1046_valid_reg;
  assign line_1047_clock = clock;
  assign line_1047_reset = reset;
  assign line_1047_valid = 2'h1 == _T_4 ^ line_1047_valid_reg;
  assign line_1048_clock = clock;
  assign line_1048_reset = reset;
  assign line_1048_valid = 2'h2 == _T_4 ^ line_1048_valid_reg;
  assign line_1049_clock = clock;
  assign line_1049_reset = reset;
  assign line_1049_valid = 2'h3 == _T_4 ^ line_1049_valid_reg;
  assign line_1050_clock = clock;
  assign line_1050_reset = reset;
  assign line_1050_valid = 2'h0 == _T_4 ^ line_1050_valid_reg;
  assign line_1051_clock = clock;
  assign line_1051_reset = reset;
  assign line_1051_valid = 2'h1 == _T_4 ^ line_1051_valid_reg;
  assign line_1052_clock = clock;
  assign line_1052_reset = reset;
  assign line_1052_valid = 2'h2 == _T_4 ^ line_1052_valid_reg;
  assign line_1053_clock = clock;
  assign line_1053_reset = reset;
  assign line_1053_valid = 2'h3 == _T_4 ^ line_1053_valid_reg;
  assign line_1054_clock = clock;
  assign line_1054_reset = reset;
  assign line_1054_valid = 2'h0 == _T_4 ^ line_1054_valid_reg;
  assign line_1055_clock = clock;
  assign line_1055_reset = reset;
  assign line_1055_valid = 2'h1 == _T_4 ^ line_1055_valid_reg;
  assign line_1056_clock = clock;
  assign line_1056_reset = reset;
  assign line_1056_valid = 2'h2 == _T_4 ^ line_1056_valid_reg;
  assign line_1057_clock = clock;
  assign line_1057_reset = reset;
  assign line_1057_valid = 2'h3 == _T_4 ^ line_1057_valid_reg;
  assign line_1058_clock = clock;
  assign line_1058_reset = reset;
  assign line_1058_valid = 2'h0 == _T_4 ^ line_1058_valid_reg;
  assign line_1059_clock = clock;
  assign line_1059_reset = reset;
  assign line_1059_valid = 2'h1 == _T_4 ^ line_1059_valid_reg;
  assign line_1060_clock = clock;
  assign line_1060_reset = reset;
  assign line_1060_valid = 2'h2 == _T_4 ^ line_1060_valid_reg;
  assign line_1061_clock = clock;
  assign line_1061_reset = reset;
  assign line_1061_valid = 2'h3 == _T_4 ^ line_1061_valid_reg;
  assign line_1062_clock = clock;
  assign line_1062_reset = reset;
  assign line_1062_valid = 2'h0 == _T_4 ^ line_1062_valid_reg;
  assign line_1063_clock = clock;
  assign line_1063_reset = reset;
  assign line_1063_valid = 2'h1 == _T_4 ^ line_1063_valid_reg;
  assign line_1064_clock = clock;
  assign line_1064_reset = reset;
  assign line_1064_valid = 2'h2 == _T_4 ^ line_1064_valid_reg;
  assign line_1065_clock = clock;
  assign line_1065_reset = reset;
  assign line_1065_valid = 2'h3 == _T_4 ^ line_1065_valid_reg;
  assign line_1066_clock = clock;
  assign line_1066_reset = reset;
  assign line_1066_valid = 2'h0 == _T_4 ^ line_1066_valid_reg;
  assign line_1067_clock = clock;
  assign line_1067_reset = reset;
  assign line_1067_valid = 2'h1 == _T_4 ^ line_1067_valid_reg;
  assign line_1068_clock = clock;
  assign line_1068_reset = reset;
  assign line_1068_valid = 2'h2 == _T_4 ^ line_1068_valid_reg;
  assign line_1069_clock = clock;
  assign line_1069_reset = reset;
  assign line_1069_valid = 2'h3 == _T_4 ^ line_1069_valid_reg;
  assign line_1070_clock = clock;
  assign line_1070_reset = reset;
  assign line_1070_valid = 2'h0 == _T_4 ^ line_1070_valid_reg;
  assign line_1071_clock = clock;
  assign line_1071_reset = reset;
  assign line_1071_valid = 2'h1 == _T_4 ^ line_1071_valid_reg;
  assign line_1072_clock = clock;
  assign line_1072_reset = reset;
  assign line_1072_valid = 2'h2 == _T_4 ^ line_1072_valid_reg;
  assign line_1073_clock = clock;
  assign line_1073_reset = reset;
  assign line_1073_valid = 2'h3 == _T_4 ^ line_1073_valid_reg;
  assign line_1074_clock = clock;
  assign line_1074_reset = reset;
  assign line_1074_valid = 2'h0 == _T_4 ^ line_1074_valid_reg;
  assign line_1075_clock = clock;
  assign line_1075_reset = reset;
  assign line_1075_valid = 2'h1 == _T_4 ^ line_1075_valid_reg;
  assign line_1076_clock = clock;
  assign line_1076_reset = reset;
  assign line_1076_valid = 2'h2 == _T_4 ^ line_1076_valid_reg;
  assign line_1077_clock = clock;
  assign line_1077_reset = reset;
  assign line_1077_valid = 2'h3 == _T_4 ^ line_1077_valid_reg;
  assign line_1078_clock = clock;
  assign line_1078_reset = reset;
  assign line_1078_valid = 2'h0 == _T_4 ^ line_1078_valid_reg;
  assign line_1079_clock = clock;
  assign line_1079_reset = reset;
  assign line_1079_valid = 2'h1 == _T_4 ^ line_1079_valid_reg;
  assign line_1080_clock = clock;
  assign line_1080_reset = reset;
  assign line_1080_valid = 2'h2 == _T_4 ^ line_1080_valid_reg;
  assign line_1081_clock = clock;
  assign line_1081_reset = reset;
  assign line_1081_valid = 2'h3 == _T_4 ^ line_1081_valid_reg;
  assign line_1082_clock = clock;
  assign line_1082_reset = reset;
  assign line_1082_valid = 2'h0 == _T_4 ^ line_1082_valid_reg;
  assign line_1083_clock = clock;
  assign line_1083_reset = reset;
  assign line_1083_valid = 2'h1 == _T_4 ^ line_1083_valid_reg;
  assign line_1084_clock = clock;
  assign line_1084_reset = reset;
  assign line_1084_valid = 2'h2 == _T_4 ^ line_1084_valid_reg;
  assign line_1085_clock = clock;
  assign line_1085_reset = reset;
  assign line_1085_valid = 2'h3 == _T_4 ^ line_1085_valid_reg;
  assign line_1086_clock = clock;
  assign line_1086_reset = reset;
  assign line_1086_valid = 2'h0 == _T_4 ^ line_1086_valid_reg;
  assign line_1087_clock = clock;
  assign line_1087_reset = reset;
  assign line_1087_valid = 2'h1 == _T_4 ^ line_1087_valid_reg;
  assign line_1088_clock = clock;
  assign line_1088_reset = reset;
  assign line_1088_valid = 2'h2 == _T_4 ^ line_1088_valid_reg;
  assign line_1089_clock = clock;
  assign line_1089_reset = reset;
  assign line_1089_valid = 2'h3 == _T_4 ^ line_1089_valid_reg;
  assign line_1090_clock = clock;
  assign line_1090_reset = reset;
  assign line_1090_valid = 2'h0 == _T_4 ^ line_1090_valid_reg;
  assign line_1091_clock = clock;
  assign line_1091_reset = reset;
  assign line_1091_valid = 2'h1 == _T_4 ^ line_1091_valid_reg;
  assign line_1092_clock = clock;
  assign line_1092_reset = reset;
  assign line_1092_valid = 2'h2 == _T_4 ^ line_1092_valid_reg;
  assign line_1093_clock = clock;
  assign line_1093_reset = reset;
  assign line_1093_valid = 2'h3 == _T_4 ^ line_1093_valid_reg;
  assign line_1094_clock = clock;
  assign line_1094_reset = reset;
  assign line_1094_valid = 2'h0 == _T_4 ^ line_1094_valid_reg;
  assign line_1095_clock = clock;
  assign line_1095_reset = reset;
  assign line_1095_valid = 2'h1 == _T_4 ^ line_1095_valid_reg;
  assign line_1096_clock = clock;
  assign line_1096_reset = reset;
  assign line_1096_valid = 2'h2 == _T_4 ^ line_1096_valid_reg;
  assign line_1097_clock = clock;
  assign line_1097_reset = reset;
  assign line_1097_valid = 2'h3 == _T_4 ^ line_1097_valid_reg;
  assign line_1098_clock = clock;
  assign line_1098_reset = reset;
  assign line_1098_valid = 2'h0 == _T_4 ^ line_1098_valid_reg;
  assign line_1099_clock = clock;
  assign line_1099_reset = reset;
  assign line_1099_valid = 2'h1 == _T_4 ^ line_1099_valid_reg;
  assign line_1100_clock = clock;
  assign line_1100_reset = reset;
  assign line_1100_valid = 2'h2 == _T_4 ^ line_1100_valid_reg;
  assign line_1101_clock = clock;
  assign line_1101_reset = reset;
  assign line_1101_valid = 2'h3 == _T_4 ^ line_1101_valid_reg;
  assign line_1102_clock = clock;
  assign line_1102_reset = reset;
  assign line_1102_valid = 2'h0 == _T_4 ^ line_1102_valid_reg;
  assign line_1103_clock = clock;
  assign line_1103_reset = reset;
  assign line_1103_valid = 2'h1 == _T_4 ^ line_1103_valid_reg;
  assign line_1104_clock = clock;
  assign line_1104_reset = reset;
  assign line_1104_valid = 2'h2 == _T_4 ^ line_1104_valid_reg;
  assign line_1105_clock = clock;
  assign line_1105_reset = reset;
  assign line_1105_valid = 2'h3 == _T_4 ^ line_1105_valid_reg;
  assign line_1106_clock = clock;
  assign line_1106_reset = reset;
  assign line_1106_valid = 2'h0 == _T_4 ^ line_1106_valid_reg;
  assign line_1107_clock = clock;
  assign line_1107_reset = reset;
  assign line_1107_valid = 2'h1 == _T_4 ^ line_1107_valid_reg;
  assign line_1108_clock = clock;
  assign line_1108_reset = reset;
  assign line_1108_valid = 2'h2 == _T_4 ^ line_1108_valid_reg;
  assign line_1109_clock = clock;
  assign line_1109_reset = reset;
  assign line_1109_valid = 2'h3 == _T_4 ^ line_1109_valid_reg;
  assign line_1110_clock = clock;
  assign line_1110_reset = reset;
  assign line_1110_valid = 2'h0 == _T_4 ^ line_1110_valid_reg;
  assign line_1111_clock = clock;
  assign line_1111_reset = reset;
  assign line_1111_valid = 2'h1 == _T_4 ^ line_1111_valid_reg;
  assign line_1112_clock = clock;
  assign line_1112_reset = reset;
  assign line_1112_valid = 2'h2 == _T_4 ^ line_1112_valid_reg;
  assign line_1113_clock = clock;
  assign line_1113_reset = reset;
  assign line_1113_valid = 2'h3 == _T_4 ^ line_1113_valid_reg;
  assign line_1114_clock = clock;
  assign line_1114_reset = reset;
  assign line_1114_valid = 2'h0 == _T_4 ^ line_1114_valid_reg;
  assign line_1115_clock = clock;
  assign line_1115_reset = reset;
  assign line_1115_valid = 2'h1 == _T_4 ^ line_1115_valid_reg;
  assign line_1116_clock = clock;
  assign line_1116_reset = reset;
  assign line_1116_valid = 2'h2 == _T_4 ^ line_1116_valid_reg;
  assign line_1117_clock = clock;
  assign line_1117_reset = reset;
  assign line_1117_valid = 2'h3 == _T_4 ^ line_1117_valid_reg;
  assign line_1118_clock = clock;
  assign line_1118_reset = reset;
  assign line_1118_valid = 2'h0 == _T_4 ^ line_1118_valid_reg;
  assign line_1119_clock = clock;
  assign line_1119_reset = reset;
  assign line_1119_valid = 2'h1 == _T_4 ^ line_1119_valid_reg;
  assign line_1120_clock = clock;
  assign line_1120_reset = reset;
  assign line_1120_valid = 2'h2 == _T_4 ^ line_1120_valid_reg;
  assign line_1121_clock = clock;
  assign line_1121_reset = reset;
  assign line_1121_valid = 2'h3 == _T_4 ^ line_1121_valid_reg;
  assign line_1122_clock = clock;
  assign line_1122_reset = reset;
  assign line_1122_valid = 2'h0 == _T_4 ^ line_1122_valid_reg;
  assign line_1123_clock = clock;
  assign line_1123_reset = reset;
  assign line_1123_valid = 2'h1 == _T_4 ^ line_1123_valid_reg;
  assign line_1124_clock = clock;
  assign line_1124_reset = reset;
  assign line_1124_valid = 2'h2 == _T_4 ^ line_1124_valid_reg;
  assign line_1125_clock = clock;
  assign line_1125_reset = reset;
  assign line_1125_valid = 2'h3 == _T_4 ^ line_1125_valid_reg;
  assign line_1126_clock = clock;
  assign line_1126_reset = reset;
  assign line_1126_valid = 2'h0 == _T_4 ^ line_1126_valid_reg;
  assign line_1127_clock = clock;
  assign line_1127_reset = reset;
  assign line_1127_valid = 2'h1 == _T_4 ^ line_1127_valid_reg;
  assign line_1128_clock = clock;
  assign line_1128_reset = reset;
  assign line_1128_valid = 2'h2 == _T_4 ^ line_1128_valid_reg;
  assign line_1129_clock = clock;
  assign line_1129_reset = reset;
  assign line_1129_valid = 2'h3 == _T_4 ^ line_1129_valid_reg;
  assign line_1130_clock = clock;
  assign line_1130_reset = reset;
  assign line_1130_valid = 2'h0 == _T_4 ^ line_1130_valid_reg;
  assign line_1131_clock = clock;
  assign line_1131_reset = reset;
  assign line_1131_valid = 2'h1 == _T_4 ^ line_1131_valid_reg;
  assign line_1132_clock = clock;
  assign line_1132_reset = reset;
  assign line_1132_valid = 2'h2 == _T_4 ^ line_1132_valid_reg;
  assign line_1133_clock = clock;
  assign line_1133_reset = reset;
  assign line_1133_valid = 2'h3 == _T_4 ^ line_1133_valid_reg;
  assign line_1134_clock = clock;
  assign line_1134_reset = reset;
  assign line_1134_valid = 2'h0 == _T_4 ^ line_1134_valid_reg;
  assign line_1135_clock = clock;
  assign line_1135_reset = reset;
  assign line_1135_valid = 2'h1 == _T_4 ^ line_1135_valid_reg;
  assign line_1136_clock = clock;
  assign line_1136_reset = reset;
  assign line_1136_valid = 2'h2 == _T_4 ^ line_1136_valid_reg;
  assign line_1137_clock = clock;
  assign line_1137_reset = reset;
  assign line_1137_valid = 2'h3 == _T_4 ^ line_1137_valid_reg;
  assign line_1138_clock = clock;
  assign line_1138_reset = reset;
  assign line_1138_valid = 2'h0 == _T_4 ^ line_1138_valid_reg;
  assign line_1139_clock = clock;
  assign line_1139_reset = reset;
  assign line_1139_valid = 2'h1 == _T_4 ^ line_1139_valid_reg;
  assign line_1140_clock = clock;
  assign line_1140_reset = reset;
  assign line_1140_valid = 2'h2 == _T_4 ^ line_1140_valid_reg;
  assign line_1141_clock = clock;
  assign line_1141_reset = reset;
  assign line_1141_valid = 2'h3 == _T_4 ^ line_1141_valid_reg;
  assign line_1142_clock = clock;
  assign line_1142_reset = reset;
  assign line_1142_valid = 2'h0 == _T_4 ^ line_1142_valid_reg;
  assign line_1143_clock = clock;
  assign line_1143_reset = reset;
  assign line_1143_valid = 2'h1 == _T_4 ^ line_1143_valid_reg;
  assign line_1144_clock = clock;
  assign line_1144_reset = reset;
  assign line_1144_valid = 2'h2 == _T_4 ^ line_1144_valid_reg;
  assign line_1145_clock = clock;
  assign line_1145_reset = reset;
  assign line_1145_valid = 2'h3 == _T_4 ^ line_1145_valid_reg;
  assign line_1146_clock = clock;
  assign line_1146_reset = reset;
  assign line_1146_valid = 2'h0 == _T_4 ^ line_1146_valid_reg;
  assign line_1147_clock = clock;
  assign line_1147_reset = reset;
  assign line_1147_valid = 2'h1 == _T_4 ^ line_1147_valid_reg;
  assign line_1148_clock = clock;
  assign line_1148_reset = reset;
  assign line_1148_valid = 2'h2 == _T_4 ^ line_1148_valid_reg;
  assign line_1149_clock = clock;
  assign line_1149_reset = reset;
  assign line_1149_valid = 2'h3 == _T_4 ^ line_1149_valid_reg;
  assign line_1150_clock = clock;
  assign line_1150_reset = reset;
  assign line_1150_valid = 2'h0 == _T_4 ^ line_1150_valid_reg;
  assign line_1151_clock = clock;
  assign line_1151_reset = reset;
  assign line_1151_valid = 2'h1 == _T_4 ^ line_1151_valid_reg;
  assign line_1152_clock = clock;
  assign line_1152_reset = reset;
  assign line_1152_valid = 2'h2 == _T_4 ^ line_1152_valid_reg;
  assign line_1153_clock = clock;
  assign line_1153_reset = reset;
  assign line_1153_valid = 2'h3 == _T_4 ^ line_1153_valid_reg;
  assign line_1154_clock = clock;
  assign line_1154_reset = reset;
  assign line_1154_valid = 2'h0 == _T_4 ^ line_1154_valid_reg;
  assign line_1155_clock = clock;
  assign line_1155_reset = reset;
  assign line_1155_valid = 2'h1 == _T_4 ^ line_1155_valid_reg;
  assign line_1156_clock = clock;
  assign line_1156_reset = reset;
  assign line_1156_valid = 2'h2 == _T_4 ^ line_1156_valid_reg;
  assign line_1157_clock = clock;
  assign line_1157_reset = reset;
  assign line_1157_valid = 2'h3 == _T_4 ^ line_1157_valid_reg;
  assign line_1158_clock = clock;
  assign line_1158_reset = reset;
  assign line_1158_valid = 2'h0 == _T_4 ^ line_1158_valid_reg;
  assign line_1159_clock = clock;
  assign line_1159_reset = reset;
  assign line_1159_valid = 2'h1 == _T_4 ^ line_1159_valid_reg;
  assign line_1160_clock = clock;
  assign line_1160_reset = reset;
  assign line_1160_valid = 2'h2 == _T_4 ^ line_1160_valid_reg;
  assign line_1161_clock = clock;
  assign line_1161_reset = reset;
  assign line_1161_valid = 2'h3 == _T_4 ^ line_1161_valid_reg;
  assign line_1162_clock = clock;
  assign line_1162_reset = reset;
  assign line_1162_valid = 2'h0 == _T_4 ^ line_1162_valid_reg;
  assign line_1163_clock = clock;
  assign line_1163_reset = reset;
  assign line_1163_valid = 2'h1 == _T_4 ^ line_1163_valid_reg;
  assign line_1164_clock = clock;
  assign line_1164_reset = reset;
  assign line_1164_valid = 2'h2 == _T_4 ^ line_1164_valid_reg;
  assign line_1165_clock = clock;
  assign line_1165_reset = reset;
  assign line_1165_valid = 2'h3 == _T_4 ^ line_1165_valid_reg;
  assign line_1166_clock = clock;
  assign line_1166_reset = reset;
  assign line_1166_valid = 2'h0 == _T_4 ^ line_1166_valid_reg;
  assign line_1167_clock = clock;
  assign line_1167_reset = reset;
  assign line_1167_valid = 2'h1 == _T_4 ^ line_1167_valid_reg;
  assign line_1168_clock = clock;
  assign line_1168_reset = reset;
  assign line_1168_valid = 2'h2 == _T_4 ^ line_1168_valid_reg;
  assign line_1169_clock = clock;
  assign line_1169_reset = reset;
  assign line_1169_valid = 2'h3 == _T_4 ^ line_1169_valid_reg;
  assign line_1170_clock = clock;
  assign line_1170_reset = reset;
  assign line_1170_valid = 2'h0 == _T_4 ^ line_1170_valid_reg;
  assign line_1171_clock = clock;
  assign line_1171_reset = reset;
  assign line_1171_valid = 2'h1 == _T_4 ^ line_1171_valid_reg;
  assign line_1172_clock = clock;
  assign line_1172_reset = reset;
  assign line_1172_valid = 2'h2 == _T_4 ^ line_1172_valid_reg;
  assign line_1173_clock = clock;
  assign line_1173_reset = reset;
  assign line_1173_valid = 2'h3 == _T_4 ^ line_1173_valid_reg;
  assign line_1174_clock = clock;
  assign line_1174_reset = reset;
  assign line_1174_valid = 2'h0 == _T_4 ^ line_1174_valid_reg;
  assign line_1175_clock = clock;
  assign line_1175_reset = reset;
  assign line_1175_valid = 2'h1 == _T_4 ^ line_1175_valid_reg;
  assign line_1176_clock = clock;
  assign line_1176_reset = reset;
  assign line_1176_valid = 2'h2 == _T_4 ^ line_1176_valid_reg;
  assign line_1177_clock = clock;
  assign line_1177_reset = reset;
  assign line_1177_valid = 2'h3 == _T_4 ^ line_1177_valid_reg;
  assign line_1178_clock = clock;
  assign line_1178_reset = reset;
  assign line_1178_valid = 2'h0 == ringBufferTail ^ line_1178_valid_reg;
  assign line_1179_clock = clock;
  assign line_1179_reset = reset;
  assign line_1179_valid = 2'h1 == ringBufferTail ^ line_1179_valid_reg;
  assign line_1180_clock = clock;
  assign line_1180_reset = reset;
  assign line_1180_valid = 2'h2 == ringBufferTail ^ line_1180_valid_reg;
  assign line_1181_clock = clock;
  assign line_1181_reset = reset;
  assign line_1181_valid = 2'h3 == ringBufferTail ^ line_1181_valid_reg;
  assign line_1182_clock = clock;
  assign line_1182_reset = reset;
  assign line_1182_valid = 2'h0 == ringBufferTail ^ line_1182_valid_reg;
  assign line_1183_clock = clock;
  assign line_1183_reset = reset;
  assign line_1183_valid = 2'h1 == ringBufferTail ^ line_1183_valid_reg;
  assign line_1184_clock = clock;
  assign line_1184_reset = reset;
  assign line_1184_valid = 2'h2 == ringBufferTail ^ line_1184_valid_reg;
  assign line_1185_clock = clock;
  assign line_1185_reset = reset;
  assign line_1185_valid = 2'h3 == ringBufferTail ^ line_1185_valid_reg;
  assign line_1186_clock = clock;
  assign line_1186_reset = reset;
  assign line_1186_valid = 2'h0 == ringBufferTail ^ line_1186_valid_reg;
  assign line_1187_clock = clock;
  assign line_1187_reset = reset;
  assign line_1187_valid = 2'h1 == ringBufferTail ^ line_1187_valid_reg;
  assign line_1188_clock = clock;
  assign line_1188_reset = reset;
  assign line_1188_valid = 2'h2 == ringBufferTail ^ line_1188_valid_reg;
  assign line_1189_clock = clock;
  assign line_1189_reset = reset;
  assign line_1189_valid = 2'h3 == ringBufferTail ^ line_1189_valid_reg;
  assign line_1190_clock = clock;
  assign line_1190_reset = reset;
  assign line_1190_valid = 2'h0 == ringBufferTail ^ line_1190_valid_reg;
  assign line_1191_clock = clock;
  assign line_1191_reset = reset;
  assign line_1191_valid = 2'h1 == ringBufferTail ^ line_1191_valid_reg;
  assign line_1192_clock = clock;
  assign line_1192_reset = reset;
  assign line_1192_valid = 2'h2 == ringBufferTail ^ line_1192_valid_reg;
  assign line_1193_clock = clock;
  assign line_1193_reset = reset;
  assign line_1193_valid = 2'h3 == ringBufferTail ^ line_1193_valid_reg;
  assign line_1194_clock = clock;
  assign line_1194_reset = reset;
  assign line_1194_valid = 2'h0 == ringBufferTail ^ line_1194_valid_reg;
  assign line_1195_clock = clock;
  assign line_1195_reset = reset;
  assign line_1195_valid = 2'h1 == ringBufferTail ^ line_1195_valid_reg;
  assign line_1196_clock = clock;
  assign line_1196_reset = reset;
  assign line_1196_valid = 2'h2 == ringBufferTail ^ line_1196_valid_reg;
  assign line_1197_clock = clock;
  assign line_1197_reset = reset;
  assign line_1197_valid = 2'h3 == ringBufferTail ^ line_1197_valid_reg;
  assign line_1198_clock = clock;
  assign line_1198_reset = reset;
  assign line_1198_valid = 2'h0 == ringBufferTail ^ line_1198_valid_reg;
  assign line_1199_clock = clock;
  assign line_1199_reset = reset;
  assign line_1199_valid = 2'h1 == ringBufferTail ^ line_1199_valid_reg;
  assign line_1200_clock = clock;
  assign line_1200_reset = reset;
  assign line_1200_valid = 2'h2 == ringBufferTail ^ line_1200_valid_reg;
  assign line_1201_clock = clock;
  assign line_1201_reset = reset;
  assign line_1201_valid = 2'h3 == ringBufferTail ^ line_1201_valid_reg;
  assign line_1202_clock = clock;
  assign line_1202_reset = reset;
  assign line_1202_valid = 2'h0 == ringBufferTail ^ line_1202_valid_reg;
  assign line_1203_clock = clock;
  assign line_1203_reset = reset;
  assign line_1203_valid = 2'h1 == ringBufferTail ^ line_1203_valid_reg;
  assign line_1204_clock = clock;
  assign line_1204_reset = reset;
  assign line_1204_valid = 2'h2 == ringBufferTail ^ line_1204_valid_reg;
  assign line_1205_clock = clock;
  assign line_1205_reset = reset;
  assign line_1205_valid = 2'h3 == ringBufferTail ^ line_1205_valid_reg;
  assign line_1206_clock = clock;
  assign line_1206_reset = reset;
  assign line_1206_valid = 2'h0 == ringBufferTail ^ line_1206_valid_reg;
  assign line_1207_clock = clock;
  assign line_1207_reset = reset;
  assign line_1207_valid = 2'h1 == ringBufferTail ^ line_1207_valid_reg;
  assign line_1208_clock = clock;
  assign line_1208_reset = reset;
  assign line_1208_valid = 2'h2 == ringBufferTail ^ line_1208_valid_reg;
  assign line_1209_clock = clock;
  assign line_1209_reset = reset;
  assign line_1209_valid = 2'h3 == ringBufferTail ^ line_1209_valid_reg;
  assign line_1210_clock = clock;
  assign line_1210_reset = reset;
  assign line_1210_valid = 2'h0 == ringBufferTail ^ line_1210_valid_reg;
  assign line_1211_clock = clock;
  assign line_1211_reset = reset;
  assign line_1211_valid = 2'h1 == ringBufferTail ^ line_1211_valid_reg;
  assign line_1212_clock = clock;
  assign line_1212_reset = reset;
  assign line_1212_valid = 2'h2 == ringBufferTail ^ line_1212_valid_reg;
  assign line_1213_clock = clock;
  assign line_1213_reset = reset;
  assign line_1213_valid = 2'h3 == ringBufferTail ^ line_1213_valid_reg;
  assign line_1214_clock = clock;
  assign line_1214_reset = reset;
  assign line_1214_valid = 2'h0 == ringBufferTail ^ line_1214_valid_reg;
  assign line_1215_clock = clock;
  assign line_1215_reset = reset;
  assign line_1215_valid = 2'h1 == ringBufferTail ^ line_1215_valid_reg;
  assign line_1216_clock = clock;
  assign line_1216_reset = reset;
  assign line_1216_valid = 2'h2 == ringBufferTail ^ line_1216_valid_reg;
  assign line_1217_clock = clock;
  assign line_1217_reset = reset;
  assign line_1217_valid = 2'h3 == ringBufferTail ^ line_1217_valid_reg;
  assign line_1218_clock = clock;
  assign line_1218_reset = reset;
  assign line_1218_valid = 2'h0 == ringBufferTail ^ line_1218_valid_reg;
  assign line_1219_clock = clock;
  assign line_1219_reset = reset;
  assign line_1219_valid = 2'h1 == ringBufferTail ^ line_1219_valid_reg;
  assign line_1220_clock = clock;
  assign line_1220_reset = reset;
  assign line_1220_valid = 2'h2 == ringBufferTail ^ line_1220_valid_reg;
  assign line_1221_clock = clock;
  assign line_1221_reset = reset;
  assign line_1221_valid = 2'h3 == ringBufferTail ^ line_1221_valid_reg;
  assign line_1222_clock = clock;
  assign line_1222_reset = reset;
  assign line_1222_valid = 2'h0 == ringBufferTail ^ line_1222_valid_reg;
  assign line_1223_clock = clock;
  assign line_1223_reset = reset;
  assign line_1223_valid = 2'h1 == ringBufferTail ^ line_1223_valid_reg;
  assign line_1224_clock = clock;
  assign line_1224_reset = reset;
  assign line_1224_valid = 2'h2 == ringBufferTail ^ line_1224_valid_reg;
  assign line_1225_clock = clock;
  assign line_1225_reset = reset;
  assign line_1225_valid = 2'h3 == ringBufferTail ^ line_1225_valid_reg;
  assign line_1226_clock = clock;
  assign line_1226_reset = reset;
  assign line_1226_valid = 2'h0 == ringBufferTail ^ line_1226_valid_reg;
  assign line_1227_clock = clock;
  assign line_1227_reset = reset;
  assign line_1227_valid = 2'h1 == ringBufferTail ^ line_1227_valid_reg;
  assign line_1228_clock = clock;
  assign line_1228_reset = reset;
  assign line_1228_valid = 2'h2 == ringBufferTail ^ line_1228_valid_reg;
  assign line_1229_clock = clock;
  assign line_1229_reset = reset;
  assign line_1229_valid = 2'h3 == ringBufferTail ^ line_1229_valid_reg;
  assign line_1230_clock = clock;
  assign line_1230_reset = reset;
  assign line_1230_valid = 2'h0 == ringBufferTail ^ line_1230_valid_reg;
  assign line_1231_clock = clock;
  assign line_1231_reset = reset;
  assign line_1231_valid = 2'h1 == ringBufferTail ^ line_1231_valid_reg;
  assign line_1232_clock = clock;
  assign line_1232_reset = reset;
  assign line_1232_valid = 2'h2 == ringBufferTail ^ line_1232_valid_reg;
  assign line_1233_clock = clock;
  assign line_1233_reset = reset;
  assign line_1233_valid = 2'h3 == ringBufferTail ^ line_1233_valid_reg;
  assign line_1234_clock = clock;
  assign line_1234_reset = reset;
  assign line_1234_valid = 2'h0 == ringBufferTail ^ line_1234_valid_reg;
  assign line_1235_clock = clock;
  assign line_1235_reset = reset;
  assign line_1235_valid = 2'h1 == ringBufferTail ^ line_1235_valid_reg;
  assign line_1236_clock = clock;
  assign line_1236_reset = reset;
  assign line_1236_valid = 2'h2 == ringBufferTail ^ line_1236_valid_reg;
  assign line_1237_clock = clock;
  assign line_1237_reset = reset;
  assign line_1237_valid = 2'h3 == ringBufferTail ^ line_1237_valid_reg;
  assign line_1238_clock = clock;
  assign line_1238_reset = reset;
  assign line_1238_valid = 2'h0 == ringBufferTail ^ line_1238_valid_reg;
  assign line_1239_clock = clock;
  assign line_1239_reset = reset;
  assign line_1239_valid = 2'h1 == ringBufferTail ^ line_1239_valid_reg;
  assign line_1240_clock = clock;
  assign line_1240_reset = reset;
  assign line_1240_valid = 2'h2 == ringBufferTail ^ line_1240_valid_reg;
  assign line_1241_clock = clock;
  assign line_1241_reset = reset;
  assign line_1241_valid = 2'h3 == ringBufferTail ^ line_1241_valid_reg;
  assign line_1242_clock = clock;
  assign line_1242_reset = reset;
  assign line_1242_valid = 2'h0 == ringBufferTail ^ line_1242_valid_reg;
  assign line_1243_clock = clock;
  assign line_1243_reset = reset;
  assign line_1243_valid = 2'h1 == ringBufferTail ^ line_1243_valid_reg;
  assign line_1244_clock = clock;
  assign line_1244_reset = reset;
  assign line_1244_valid = 2'h2 == ringBufferTail ^ line_1244_valid_reg;
  assign line_1245_clock = clock;
  assign line_1245_reset = reset;
  assign line_1245_valid = 2'h3 == ringBufferTail ^ line_1245_valid_reg;
  assign line_1246_clock = clock;
  assign line_1246_reset = reset;
  assign line_1246_valid = 2'h0 == ringBufferTail ^ line_1246_valid_reg;
  assign line_1247_clock = clock;
  assign line_1247_reset = reset;
  assign line_1247_valid = 2'h1 == ringBufferTail ^ line_1247_valid_reg;
  assign line_1248_clock = clock;
  assign line_1248_reset = reset;
  assign line_1248_valid = 2'h2 == ringBufferTail ^ line_1248_valid_reg;
  assign line_1249_clock = clock;
  assign line_1249_reset = reset;
  assign line_1249_valid = 2'h3 == ringBufferTail ^ line_1249_valid_reg;
  assign line_1250_clock = clock;
  assign line_1250_reset = reset;
  assign line_1250_valid = 2'h0 == ringBufferTail ^ line_1250_valid_reg;
  assign line_1251_clock = clock;
  assign line_1251_reset = reset;
  assign line_1251_valid = 2'h1 == ringBufferTail ^ line_1251_valid_reg;
  assign line_1252_clock = clock;
  assign line_1252_reset = reset;
  assign line_1252_valid = 2'h2 == ringBufferTail ^ line_1252_valid_reg;
  assign line_1253_clock = clock;
  assign line_1253_reset = reset;
  assign line_1253_valid = 2'h3 == ringBufferTail ^ line_1253_valid_reg;
  assign line_1254_clock = clock;
  assign line_1254_reset = reset;
  assign line_1254_valid = 2'h0 == ringBufferTail ^ line_1254_valid_reg;
  assign line_1255_clock = clock;
  assign line_1255_reset = reset;
  assign line_1255_valid = 2'h1 == ringBufferTail ^ line_1255_valid_reg;
  assign line_1256_clock = clock;
  assign line_1256_reset = reset;
  assign line_1256_valid = 2'h2 == ringBufferTail ^ line_1256_valid_reg;
  assign line_1257_clock = clock;
  assign line_1257_reset = reset;
  assign line_1257_valid = 2'h3 == ringBufferTail ^ line_1257_valid_reg;
  assign line_1258_clock = clock;
  assign line_1258_reset = reset;
  assign line_1258_valid = 2'h0 == ringBufferTail ^ line_1258_valid_reg;
  assign line_1259_clock = clock;
  assign line_1259_reset = reset;
  assign line_1259_valid = 2'h1 == ringBufferTail ^ line_1259_valid_reg;
  assign line_1260_clock = clock;
  assign line_1260_reset = reset;
  assign line_1260_valid = 2'h2 == ringBufferTail ^ line_1260_valid_reg;
  assign line_1261_clock = clock;
  assign line_1261_reset = reset;
  assign line_1261_valid = 2'h3 == ringBufferTail ^ line_1261_valid_reg;
  assign line_1262_clock = clock;
  assign line_1262_reset = reset;
  assign line_1262_valid = 2'h0 == ringBufferTail ^ line_1262_valid_reg;
  assign line_1263_clock = clock;
  assign line_1263_reset = reset;
  assign line_1263_valid = 2'h1 == ringBufferTail ^ line_1263_valid_reg;
  assign line_1264_clock = clock;
  assign line_1264_reset = reset;
  assign line_1264_valid = 2'h2 == ringBufferTail ^ line_1264_valid_reg;
  assign line_1265_clock = clock;
  assign line_1265_reset = reset;
  assign line_1265_valid = 2'h3 == ringBufferTail ^ line_1265_valid_reg;
  assign line_1266_clock = clock;
  assign line_1266_reset = reset;
  assign line_1266_valid = 2'h0 == ringBufferTail ^ line_1266_valid_reg;
  assign line_1267_clock = clock;
  assign line_1267_reset = reset;
  assign line_1267_valid = 2'h1 == ringBufferTail ^ line_1267_valid_reg;
  assign line_1268_clock = clock;
  assign line_1268_reset = reset;
  assign line_1268_valid = 2'h2 == ringBufferTail ^ line_1268_valid_reg;
  assign line_1269_clock = clock;
  assign line_1269_reset = reset;
  assign line_1269_valid = 2'h3 == ringBufferTail ^ line_1269_valid_reg;
  assign line_1270_clock = clock;
  assign line_1270_reset = reset;
  assign line_1270_valid = 2'h0 == ringBufferTail ^ line_1270_valid_reg;
  assign line_1271_clock = clock;
  assign line_1271_reset = reset;
  assign line_1271_valid = 2'h1 == ringBufferTail ^ line_1271_valid_reg;
  assign line_1272_clock = clock;
  assign line_1272_reset = reset;
  assign line_1272_valid = 2'h2 == ringBufferTail ^ line_1272_valid_reg;
  assign line_1273_clock = clock;
  assign line_1273_reset = reset;
  assign line_1273_valid = 2'h3 == ringBufferTail ^ line_1273_valid_reg;
  assign line_1274_clock = clock;
  assign line_1274_reset = reset;
  assign line_1274_valid = 2'h0 == ringBufferTail ^ line_1274_valid_reg;
  assign line_1275_clock = clock;
  assign line_1275_reset = reset;
  assign line_1275_valid = 2'h1 == ringBufferTail ^ line_1275_valid_reg;
  assign line_1276_clock = clock;
  assign line_1276_reset = reset;
  assign line_1276_valid = 2'h2 == ringBufferTail ^ line_1276_valid_reg;
  assign line_1277_clock = clock;
  assign line_1277_reset = reset;
  assign line_1277_valid = 2'h3 == ringBufferTail ^ line_1277_valid_reg;
  assign line_1278_clock = clock;
  assign line_1278_reset = reset;
  assign line_1278_valid = 2'h0 == ringBufferTail ^ line_1278_valid_reg;
  assign line_1279_clock = clock;
  assign line_1279_reset = reset;
  assign line_1279_valid = 2'h1 == ringBufferTail ^ line_1279_valid_reg;
  assign line_1280_clock = clock;
  assign line_1280_reset = reset;
  assign line_1280_valid = 2'h2 == ringBufferTail ^ line_1280_valid_reg;
  assign line_1281_clock = clock;
  assign line_1281_reset = reset;
  assign line_1281_valid = 2'h3 == ringBufferTail ^ line_1281_valid_reg;
  assign line_1282_clock = clock;
  assign line_1282_reset = reset;
  assign line_1282_valid = 2'h0 == ringBufferTail ^ line_1282_valid_reg;
  assign line_1283_clock = clock;
  assign line_1283_reset = reset;
  assign line_1283_valid = 2'h1 == ringBufferTail ^ line_1283_valid_reg;
  assign line_1284_clock = clock;
  assign line_1284_reset = reset;
  assign line_1284_valid = 2'h2 == ringBufferTail ^ line_1284_valid_reg;
  assign line_1285_clock = clock;
  assign line_1285_reset = reset;
  assign line_1285_valid = 2'h3 == ringBufferTail ^ line_1285_valid_reg;
  assign line_1286_clock = clock;
  assign line_1286_reset = reset;
  assign line_1286_valid = 2'h0 == ringBufferTail ^ line_1286_valid_reg;
  assign line_1287_clock = clock;
  assign line_1287_reset = reset;
  assign line_1287_valid = 2'h1 == ringBufferTail ^ line_1287_valid_reg;
  assign line_1288_clock = clock;
  assign line_1288_reset = reset;
  assign line_1288_valid = 2'h2 == ringBufferTail ^ line_1288_valid_reg;
  assign line_1289_clock = clock;
  assign line_1289_reset = reset;
  assign line_1289_valid = 2'h3 == ringBufferTail ^ line_1289_valid_reg;
  assign line_1290_clock = clock;
  assign line_1290_reset = reset;
  assign line_1290_valid = 2'h0 == ringBufferTail ^ line_1290_valid_reg;
  assign line_1291_clock = clock;
  assign line_1291_reset = reset;
  assign line_1291_valid = 2'h1 == ringBufferTail ^ line_1291_valid_reg;
  assign line_1292_clock = clock;
  assign line_1292_reset = reset;
  assign line_1292_valid = 2'h2 == ringBufferTail ^ line_1292_valid_reg;
  assign line_1293_clock = clock;
  assign line_1293_reset = reset;
  assign line_1293_valid = 2'h3 == ringBufferTail ^ line_1293_valid_reg;
  assign line_1294_clock = clock;
  assign line_1294_reset = reset;
  assign line_1294_valid = 2'h0 == ringBufferTail ^ line_1294_valid_reg;
  assign line_1295_clock = clock;
  assign line_1295_reset = reset;
  assign line_1295_valid = 2'h1 == ringBufferTail ^ line_1295_valid_reg;
  assign line_1296_clock = clock;
  assign line_1296_reset = reset;
  assign line_1296_valid = 2'h2 == ringBufferTail ^ line_1296_valid_reg;
  assign line_1297_clock = clock;
  assign line_1297_reset = reset;
  assign line_1297_valid = 2'h3 == ringBufferTail ^ line_1297_valid_reg;
  assign line_1298_clock = clock;
  assign line_1298_reset = reset;
  assign line_1298_valid = 2'h0 == ringBufferTail ^ line_1298_valid_reg;
  assign line_1299_clock = clock;
  assign line_1299_reset = reset;
  assign line_1299_valid = 2'h1 == ringBufferTail ^ line_1299_valid_reg;
  assign line_1300_clock = clock;
  assign line_1300_reset = reset;
  assign line_1300_valid = 2'h2 == ringBufferTail ^ line_1300_valid_reg;
  assign line_1301_clock = clock;
  assign line_1301_reset = reset;
  assign line_1301_valid = 2'h3 == ringBufferTail ^ line_1301_valid_reg;
  assign line_1302_clock = clock;
  assign line_1302_reset = reset;
  assign line_1302_valid = 2'h0 == ringBufferTail ^ line_1302_valid_reg;
  assign line_1303_clock = clock;
  assign line_1303_reset = reset;
  assign line_1303_valid = 2'h1 == ringBufferTail ^ line_1303_valid_reg;
  assign line_1304_clock = clock;
  assign line_1304_reset = reset;
  assign line_1304_valid = 2'h2 == ringBufferTail ^ line_1304_valid_reg;
  assign line_1305_clock = clock;
  assign line_1305_reset = reset;
  assign line_1305_valid = 2'h3 == ringBufferTail ^ line_1305_valid_reg;
  assign line_1306_clock = clock;
  assign line_1306_reset = reset;
  assign line_1306_valid = 2'h0 == ringBufferTail ^ line_1306_valid_reg;
  assign line_1307_clock = clock;
  assign line_1307_reset = reset;
  assign line_1307_valid = 2'h1 == ringBufferTail ^ line_1307_valid_reg;
  assign line_1308_clock = clock;
  assign line_1308_reset = reset;
  assign line_1308_valid = 2'h2 == ringBufferTail ^ line_1308_valid_reg;
  assign line_1309_clock = clock;
  assign line_1309_reset = reset;
  assign line_1309_valid = 2'h3 == ringBufferTail ^ line_1309_valid_reg;
  assign line_1310_clock = clock;
  assign line_1310_reset = reset;
  assign line_1310_valid = 2'h0 == ringBufferTail ^ line_1310_valid_reg;
  assign line_1311_clock = clock;
  assign line_1311_reset = reset;
  assign line_1311_valid = 2'h1 == ringBufferTail ^ line_1311_valid_reg;
  assign line_1312_clock = clock;
  assign line_1312_reset = reset;
  assign line_1312_valid = 2'h2 == ringBufferTail ^ line_1312_valid_reg;
  assign line_1313_clock = clock;
  assign line_1313_reset = reset;
  assign line_1313_valid = 2'h3 == ringBufferTail ^ line_1313_valid_reg;
  assign line_1314_clock = clock;
  assign line_1314_reset = reset;
  assign line_1314_valid = 2'h0 == ringBufferTail ^ line_1314_valid_reg;
  assign line_1315_clock = clock;
  assign line_1315_reset = reset;
  assign line_1315_valid = 2'h1 == ringBufferTail ^ line_1315_valid_reg;
  assign line_1316_clock = clock;
  assign line_1316_reset = reset;
  assign line_1316_valid = 2'h2 == ringBufferTail ^ line_1316_valid_reg;
  assign line_1317_clock = clock;
  assign line_1317_reset = reset;
  assign line_1317_valid = 2'h3 == ringBufferTail ^ line_1317_valid_reg;
  assign line_1318_clock = clock;
  assign line_1318_reset = reset;
  assign line_1318_valid = 2'h0 == ringBufferTail ^ line_1318_valid_reg;
  assign line_1319_clock = clock;
  assign line_1319_reset = reset;
  assign line_1319_valid = 2'h1 == ringBufferTail ^ line_1319_valid_reg;
  assign line_1320_clock = clock;
  assign line_1320_reset = reset;
  assign line_1320_valid = 2'h2 == ringBufferTail ^ line_1320_valid_reg;
  assign line_1321_clock = clock;
  assign line_1321_reset = reset;
  assign line_1321_valid = 2'h3 == ringBufferTail ^ line_1321_valid_reg;
  assign line_1322_clock = clock;
  assign line_1322_reset = reset;
  assign line_1322_valid = 2'h0 == ringBufferTail ^ line_1322_valid_reg;
  assign line_1323_clock = clock;
  assign line_1323_reset = reset;
  assign line_1323_valid = 2'h1 == ringBufferTail ^ line_1323_valid_reg;
  assign line_1324_clock = clock;
  assign line_1324_reset = reset;
  assign line_1324_valid = 2'h2 == ringBufferTail ^ line_1324_valid_reg;
  assign line_1325_clock = clock;
  assign line_1325_reset = reset;
  assign line_1325_valid = 2'h3 == ringBufferTail ^ line_1325_valid_reg;
  assign line_1326_clock = clock;
  assign line_1326_reset = reset;
  assign line_1326_valid = 2'h0 == ringBufferTail ^ line_1326_valid_reg;
  assign line_1327_clock = clock;
  assign line_1327_reset = reset;
  assign line_1327_valid = 2'h1 == ringBufferTail ^ line_1327_valid_reg;
  assign line_1328_clock = clock;
  assign line_1328_reset = reset;
  assign line_1328_valid = 2'h2 == ringBufferTail ^ line_1328_valid_reg;
  assign line_1329_clock = clock;
  assign line_1329_reset = reset;
  assign line_1329_valid = 2'h3 == ringBufferTail ^ line_1329_valid_reg;
  assign line_1330_clock = clock;
  assign line_1330_reset = reset;
  assign line_1330_valid = 2'h0 == ringBufferTail ^ line_1330_valid_reg;
  assign line_1331_clock = clock;
  assign line_1331_reset = reset;
  assign line_1331_valid = 2'h1 == ringBufferTail ^ line_1331_valid_reg;
  assign line_1332_clock = clock;
  assign line_1332_reset = reset;
  assign line_1332_valid = 2'h2 == ringBufferTail ^ line_1332_valid_reg;
  assign line_1333_clock = clock;
  assign line_1333_reset = reset;
  assign line_1333_valid = 2'h3 == ringBufferTail ^ line_1333_valid_reg;
  assign line_1334_clock = clock;
  assign line_1334_reset = reset;
  assign line_1334_valid = 2'h0 == ringBufferTail ^ line_1334_valid_reg;
  assign line_1335_clock = clock;
  assign line_1335_reset = reset;
  assign line_1335_valid = 2'h1 == ringBufferTail ^ line_1335_valid_reg;
  assign line_1336_clock = clock;
  assign line_1336_reset = reset;
  assign line_1336_valid = 2'h2 == ringBufferTail ^ line_1336_valid_reg;
  assign line_1337_clock = clock;
  assign line_1337_reset = reset;
  assign line_1337_valid = 2'h3 == ringBufferTail ^ line_1337_valid_reg;
  assign line_1338_clock = clock;
  assign line_1338_reset = reset;
  assign line_1338_valid = 2'h0 == ringBufferTail ^ line_1338_valid_reg;
  assign line_1339_clock = clock;
  assign line_1339_reset = reset;
  assign line_1339_valid = 2'h1 == ringBufferTail ^ line_1339_valid_reg;
  assign line_1340_clock = clock;
  assign line_1340_reset = reset;
  assign line_1340_valid = 2'h2 == ringBufferTail ^ line_1340_valid_reg;
  assign line_1341_clock = clock;
  assign line_1341_reset = reset;
  assign line_1341_valid = 2'h3 == ringBufferTail ^ line_1341_valid_reg;
  assign line_1342_clock = clock;
  assign line_1342_reset = reset;
  assign line_1342_valid = 2'h0 == ringBufferTail ^ line_1342_valid_reg;
  assign line_1343_clock = clock;
  assign line_1343_reset = reset;
  assign line_1343_valid = 2'h1 == ringBufferTail ^ line_1343_valid_reg;
  assign line_1344_clock = clock;
  assign line_1344_reset = reset;
  assign line_1344_valid = 2'h2 == ringBufferTail ^ line_1344_valid_reg;
  assign line_1345_clock = clock;
  assign line_1345_reset = reset;
  assign line_1345_valid = 2'h3 == ringBufferTail ^ line_1345_valid_reg;
  assign line_1346_clock = clock;
  assign line_1346_reset = reset;
  assign line_1346_valid = 2'h0 == ringBufferTail ^ line_1346_valid_reg;
  assign line_1347_clock = clock;
  assign line_1347_reset = reset;
  assign line_1347_valid = 2'h1 == ringBufferTail ^ line_1347_valid_reg;
  assign line_1348_clock = clock;
  assign line_1348_reset = reset;
  assign line_1348_valid = 2'h2 == ringBufferTail ^ line_1348_valid_reg;
  assign line_1349_clock = clock;
  assign line_1349_reset = reset;
  assign line_1349_valid = 2'h3 == ringBufferTail ^ line_1349_valid_reg;
  assign line_1350_clock = clock;
  assign line_1350_reset = reset;
  assign line_1350_valid = 2'h0 == ringBufferTail ^ line_1350_valid_reg;
  assign line_1351_clock = clock;
  assign line_1351_reset = reset;
  assign line_1351_valid = 2'h1 == ringBufferTail ^ line_1351_valid_reg;
  assign line_1352_clock = clock;
  assign line_1352_reset = reset;
  assign line_1352_valid = 2'h2 == ringBufferTail ^ line_1352_valid_reg;
  assign line_1353_clock = clock;
  assign line_1353_reset = reset;
  assign line_1353_valid = 2'h3 == ringBufferTail ^ line_1353_valid_reg;
  assign line_1354_clock = clock;
  assign line_1354_reset = reset;
  assign line_1354_valid = 2'h0 == ringBufferTail ^ line_1354_valid_reg;
  assign line_1355_clock = clock;
  assign line_1355_reset = reset;
  assign line_1355_valid = 2'h1 == ringBufferTail ^ line_1355_valid_reg;
  assign line_1356_clock = clock;
  assign line_1356_reset = reset;
  assign line_1356_valid = 2'h2 == ringBufferTail ^ line_1356_valid_reg;
  assign line_1357_clock = clock;
  assign line_1357_reset = reset;
  assign line_1357_valid = 2'h3 == ringBufferTail ^ line_1357_valid_reg;
  assign line_1358_clock = clock;
  assign line_1358_reset = reset;
  assign line_1358_valid = 2'h0 == ringBufferTail ^ line_1358_valid_reg;
  assign line_1359_clock = clock;
  assign line_1359_reset = reset;
  assign line_1359_valid = 2'h1 == ringBufferTail ^ line_1359_valid_reg;
  assign line_1360_clock = clock;
  assign line_1360_reset = reset;
  assign line_1360_valid = 2'h2 == ringBufferTail ^ line_1360_valid_reg;
  assign line_1361_clock = clock;
  assign line_1361_reset = reset;
  assign line_1361_valid = 2'h3 == ringBufferTail ^ line_1361_valid_reg;
  assign line_1362_clock = clock;
  assign line_1362_reset = reset;
  assign line_1362_valid = 2'h0 == ringBufferTail ^ line_1362_valid_reg;
  assign line_1363_clock = clock;
  assign line_1363_reset = reset;
  assign line_1363_valid = 2'h1 == ringBufferTail ^ line_1363_valid_reg;
  assign line_1364_clock = clock;
  assign line_1364_reset = reset;
  assign line_1364_valid = 2'h2 == ringBufferTail ^ line_1364_valid_reg;
  assign line_1365_clock = clock;
  assign line_1365_reset = reset;
  assign line_1365_valid = 2'h3 == ringBufferTail ^ line_1365_valid_reg;
  assign line_1366_clock = clock;
  assign line_1366_reset = reset;
  assign line_1366_valid = 2'h0 == ringBufferTail ^ line_1366_valid_reg;
  assign line_1367_clock = clock;
  assign line_1367_reset = reset;
  assign line_1367_valid = 2'h1 == ringBufferTail ^ line_1367_valid_reg;
  assign line_1368_clock = clock;
  assign line_1368_reset = reset;
  assign line_1368_valid = 2'h2 == ringBufferTail ^ line_1368_valid_reg;
  assign line_1369_clock = clock;
  assign line_1369_reset = reset;
  assign line_1369_valid = 2'h3 == ringBufferTail ^ line_1369_valid_reg;
  assign line_1370_clock = clock;
  assign line_1370_reset = reset;
  assign line_1370_valid = 2'h0 == ringBufferTail ^ line_1370_valid_reg;
  assign line_1371_clock = clock;
  assign line_1371_reset = reset;
  assign line_1371_valid = 2'h1 == ringBufferTail ^ line_1371_valid_reg;
  assign line_1372_clock = clock;
  assign line_1372_reset = reset;
  assign line_1372_valid = 2'h2 == ringBufferTail ^ line_1372_valid_reg;
  assign line_1373_clock = clock;
  assign line_1373_reset = reset;
  assign line_1373_valid = 2'h3 == ringBufferTail ^ line_1373_valid_reg;
  assign line_1374_clock = clock;
  assign line_1374_reset = reset;
  assign line_1374_valid = 2'h0 == ringBufferTail ^ line_1374_valid_reg;
  assign line_1375_clock = clock;
  assign line_1375_reset = reset;
  assign line_1375_valid = 2'h1 == ringBufferTail ^ line_1375_valid_reg;
  assign line_1376_clock = clock;
  assign line_1376_reset = reset;
  assign line_1376_valid = 2'h2 == ringBufferTail ^ line_1376_valid_reg;
  assign line_1377_clock = clock;
  assign line_1377_reset = reset;
  assign line_1377_valid = 2'h3 == ringBufferTail ^ line_1377_valid_reg;
  assign line_1378_clock = clock;
  assign line_1378_reset = reset;
  assign line_1378_valid = 2'h0 == ringBufferTail ^ line_1378_valid_reg;
  assign line_1379_clock = clock;
  assign line_1379_reset = reset;
  assign line_1379_valid = 2'h1 == ringBufferTail ^ line_1379_valid_reg;
  assign line_1380_clock = clock;
  assign line_1380_reset = reset;
  assign line_1380_valid = 2'h2 == ringBufferTail ^ line_1380_valid_reg;
  assign line_1381_clock = clock;
  assign line_1381_reset = reset;
  assign line_1381_valid = 2'h3 == ringBufferTail ^ line_1381_valid_reg;
  assign line_1382_clock = clock;
  assign line_1382_reset = reset;
  assign line_1382_valid = 2'h0 == ringBufferTail ^ line_1382_valid_reg;
  assign line_1383_clock = clock;
  assign line_1383_reset = reset;
  assign line_1383_valid = 2'h1 == ringBufferTail ^ line_1383_valid_reg;
  assign line_1384_clock = clock;
  assign line_1384_reset = reset;
  assign line_1384_valid = 2'h2 == ringBufferTail ^ line_1384_valid_reg;
  assign line_1385_clock = clock;
  assign line_1385_reset = reset;
  assign line_1385_valid = 2'h3 == ringBufferTail ^ line_1385_valid_reg;
  assign line_1386_clock = clock;
  assign line_1386_reset = reset;
  assign line_1386_valid = 2'h0 == ringBufferTail ^ line_1386_valid_reg;
  assign line_1387_clock = clock;
  assign line_1387_reset = reset;
  assign line_1387_valid = 2'h1 == ringBufferTail ^ line_1387_valid_reg;
  assign line_1388_clock = clock;
  assign line_1388_reset = reset;
  assign line_1388_valid = 2'h2 == ringBufferTail ^ line_1388_valid_reg;
  assign line_1389_clock = clock;
  assign line_1389_reset = reset;
  assign line_1389_valid = 2'h3 == ringBufferTail ^ line_1389_valid_reg;
  assign line_1390_clock = clock;
  assign line_1390_reset = reset;
  assign line_1390_valid = 2'h0 == ringBufferTail ^ line_1390_valid_reg;
  assign line_1391_clock = clock;
  assign line_1391_reset = reset;
  assign line_1391_valid = 2'h1 == ringBufferTail ^ line_1391_valid_reg;
  assign line_1392_clock = clock;
  assign line_1392_reset = reset;
  assign line_1392_valid = 2'h2 == ringBufferTail ^ line_1392_valid_reg;
  assign line_1393_clock = clock;
  assign line_1393_reset = reset;
  assign line_1393_valid = 2'h3 == ringBufferTail ^ line_1393_valid_reg;
  assign line_1394_clock = clock;
  assign line_1394_reset = reset;
  assign line_1394_valid = 2'h0 == ringBufferTail ^ line_1394_valid_reg;
  assign line_1395_clock = clock;
  assign line_1395_reset = reset;
  assign line_1395_valid = 2'h1 == ringBufferTail ^ line_1395_valid_reg;
  assign line_1396_clock = clock;
  assign line_1396_reset = reset;
  assign line_1396_valid = 2'h2 == ringBufferTail ^ line_1396_valid_reg;
  assign line_1397_clock = clock;
  assign line_1397_reset = reset;
  assign line_1397_valid = 2'h3 == ringBufferTail ^ line_1397_valid_reg;
  assign line_1398_clock = clock;
  assign line_1398_reset = reset;
  assign line_1398_valid = 2'h0 == ringBufferTail ^ line_1398_valid_reg;
  assign line_1399_clock = clock;
  assign line_1399_reset = reset;
  assign line_1399_valid = 2'h1 == ringBufferTail ^ line_1399_valid_reg;
  assign line_1400_clock = clock;
  assign line_1400_reset = reset;
  assign line_1400_valid = 2'h2 == ringBufferTail ^ line_1400_valid_reg;
  assign line_1401_clock = clock;
  assign line_1401_reset = reset;
  assign line_1401_valid = 2'h3 == ringBufferTail ^ line_1401_valid_reg;
  assign line_1402_clock = clock;
  assign line_1402_reset = reset;
  assign line_1402_valid = 2'h0 == deq2_StartIndex ^ line_1402_valid_reg;
  assign line_1403_clock = clock;
  assign line_1403_reset = reset;
  assign line_1403_valid = 2'h1 == deq2_StartIndex ^ line_1403_valid_reg;
  assign line_1404_clock = clock;
  assign line_1404_reset = reset;
  assign line_1404_valid = 2'h2 == deq2_StartIndex ^ line_1404_valid_reg;
  assign line_1405_clock = clock;
  assign line_1405_reset = reset;
  assign line_1405_valid = 2'h3 == deq2_StartIndex ^ line_1405_valid_reg;
  assign line_1406_clock = clock;
  assign line_1406_reset = reset;
  assign line_1406_valid = 2'h0 == deq2_StartIndex ^ line_1406_valid_reg;
  assign line_1407_clock = clock;
  assign line_1407_reset = reset;
  assign line_1407_valid = 2'h1 == deq2_StartIndex ^ line_1407_valid_reg;
  assign line_1408_clock = clock;
  assign line_1408_reset = reset;
  assign line_1408_valid = 2'h2 == deq2_StartIndex ^ line_1408_valid_reg;
  assign line_1409_clock = clock;
  assign line_1409_reset = reset;
  assign line_1409_valid = 2'h3 == deq2_StartIndex ^ line_1409_valid_reg;
  assign line_1410_clock = clock;
  assign line_1410_reset = reset;
  assign line_1410_valid = 2'h0 == deq2_StartIndex ^ line_1410_valid_reg;
  assign line_1411_clock = clock;
  assign line_1411_reset = reset;
  assign line_1411_valid = 2'h1 == deq2_StartIndex ^ line_1411_valid_reg;
  assign line_1412_clock = clock;
  assign line_1412_reset = reset;
  assign line_1412_valid = 2'h2 == deq2_StartIndex ^ line_1412_valid_reg;
  assign line_1413_clock = clock;
  assign line_1413_reset = reset;
  assign line_1413_valid = 2'h3 == deq2_StartIndex ^ line_1413_valid_reg;
  assign line_1414_clock = clock;
  assign line_1414_reset = reset;
  assign line_1414_valid = 2'h0 == deq2_StartIndex ^ line_1414_valid_reg;
  assign line_1415_clock = clock;
  assign line_1415_reset = reset;
  assign line_1415_valid = 2'h1 == deq2_StartIndex ^ line_1415_valid_reg;
  assign line_1416_clock = clock;
  assign line_1416_reset = reset;
  assign line_1416_valid = 2'h2 == deq2_StartIndex ^ line_1416_valid_reg;
  assign line_1417_clock = clock;
  assign line_1417_reset = reset;
  assign line_1417_valid = 2'h3 == deq2_StartIndex ^ line_1417_valid_reg;
  assign line_1418_clock = clock;
  assign line_1418_reset = reset;
  assign line_1418_valid = 2'h0 == deq2_StartIndex ^ line_1418_valid_reg;
  assign line_1419_clock = clock;
  assign line_1419_reset = reset;
  assign line_1419_valid = 2'h1 == deq2_StartIndex ^ line_1419_valid_reg;
  assign line_1420_clock = clock;
  assign line_1420_reset = reset;
  assign line_1420_valid = 2'h2 == deq2_StartIndex ^ line_1420_valid_reg;
  assign line_1421_clock = clock;
  assign line_1421_reset = reset;
  assign line_1421_valid = 2'h3 == deq2_StartIndex ^ line_1421_valid_reg;
  assign line_1422_clock = clock;
  assign line_1422_reset = reset;
  assign line_1422_valid = 2'h0 == deq2_StartIndex ^ line_1422_valid_reg;
  assign line_1423_clock = clock;
  assign line_1423_reset = reset;
  assign line_1423_valid = 2'h1 == deq2_StartIndex ^ line_1423_valid_reg;
  assign line_1424_clock = clock;
  assign line_1424_reset = reset;
  assign line_1424_valid = 2'h2 == deq2_StartIndex ^ line_1424_valid_reg;
  assign line_1425_clock = clock;
  assign line_1425_reset = reset;
  assign line_1425_valid = 2'h3 == deq2_StartIndex ^ line_1425_valid_reg;
  assign line_1426_clock = clock;
  assign line_1426_reset = reset;
  assign line_1426_valid = 2'h0 == deq2_StartIndex ^ line_1426_valid_reg;
  assign line_1427_clock = clock;
  assign line_1427_reset = reset;
  assign line_1427_valid = 2'h1 == deq2_StartIndex ^ line_1427_valid_reg;
  assign line_1428_clock = clock;
  assign line_1428_reset = reset;
  assign line_1428_valid = 2'h2 == deq2_StartIndex ^ line_1428_valid_reg;
  assign line_1429_clock = clock;
  assign line_1429_reset = reset;
  assign line_1429_valid = 2'h3 == deq2_StartIndex ^ line_1429_valid_reg;
  assign line_1430_clock = clock;
  assign line_1430_reset = reset;
  assign line_1430_valid = 2'h0 == deq2_StartIndex ^ line_1430_valid_reg;
  assign line_1431_clock = clock;
  assign line_1431_reset = reset;
  assign line_1431_valid = 2'h1 == deq2_StartIndex ^ line_1431_valid_reg;
  assign line_1432_clock = clock;
  assign line_1432_reset = reset;
  assign line_1432_valid = 2'h2 == deq2_StartIndex ^ line_1432_valid_reg;
  assign line_1433_clock = clock;
  assign line_1433_reset = reset;
  assign line_1433_valid = 2'h3 == deq2_StartIndex ^ line_1433_valid_reg;
  assign line_1434_clock = clock;
  assign line_1434_reset = reset;
  assign line_1434_valid = 2'h0 == deq2_StartIndex ^ line_1434_valid_reg;
  assign line_1435_clock = clock;
  assign line_1435_reset = reset;
  assign line_1435_valid = 2'h1 == deq2_StartIndex ^ line_1435_valid_reg;
  assign line_1436_clock = clock;
  assign line_1436_reset = reset;
  assign line_1436_valid = 2'h2 == deq2_StartIndex ^ line_1436_valid_reg;
  assign line_1437_clock = clock;
  assign line_1437_reset = reset;
  assign line_1437_valid = 2'h3 == deq2_StartIndex ^ line_1437_valid_reg;
  assign line_1438_clock = clock;
  assign line_1438_reset = reset;
  assign line_1438_valid = 2'h0 == deq2_StartIndex ^ line_1438_valid_reg;
  assign line_1439_clock = clock;
  assign line_1439_reset = reset;
  assign line_1439_valid = 2'h1 == deq2_StartIndex ^ line_1439_valid_reg;
  assign line_1440_clock = clock;
  assign line_1440_reset = reset;
  assign line_1440_valid = 2'h2 == deq2_StartIndex ^ line_1440_valid_reg;
  assign line_1441_clock = clock;
  assign line_1441_reset = reset;
  assign line_1441_valid = 2'h3 == deq2_StartIndex ^ line_1441_valid_reg;
  assign line_1442_clock = clock;
  assign line_1442_reset = reset;
  assign line_1442_valid = 2'h0 == deq2_StartIndex ^ line_1442_valid_reg;
  assign line_1443_clock = clock;
  assign line_1443_reset = reset;
  assign line_1443_valid = 2'h1 == deq2_StartIndex ^ line_1443_valid_reg;
  assign line_1444_clock = clock;
  assign line_1444_reset = reset;
  assign line_1444_valid = 2'h2 == deq2_StartIndex ^ line_1444_valid_reg;
  assign line_1445_clock = clock;
  assign line_1445_reset = reset;
  assign line_1445_valid = 2'h3 == deq2_StartIndex ^ line_1445_valid_reg;
  assign line_1446_clock = clock;
  assign line_1446_reset = reset;
  assign line_1446_valid = 2'h0 == deq2_StartIndex ^ line_1446_valid_reg;
  assign line_1447_clock = clock;
  assign line_1447_reset = reset;
  assign line_1447_valid = 2'h1 == deq2_StartIndex ^ line_1447_valid_reg;
  assign line_1448_clock = clock;
  assign line_1448_reset = reset;
  assign line_1448_valid = 2'h2 == deq2_StartIndex ^ line_1448_valid_reg;
  assign line_1449_clock = clock;
  assign line_1449_reset = reset;
  assign line_1449_valid = 2'h3 == deq2_StartIndex ^ line_1449_valid_reg;
  assign line_1450_clock = clock;
  assign line_1450_reset = reset;
  assign line_1450_valid = 2'h0 == deq2_StartIndex ^ line_1450_valid_reg;
  assign line_1451_clock = clock;
  assign line_1451_reset = reset;
  assign line_1451_valid = 2'h1 == deq2_StartIndex ^ line_1451_valid_reg;
  assign line_1452_clock = clock;
  assign line_1452_reset = reset;
  assign line_1452_valid = 2'h2 == deq2_StartIndex ^ line_1452_valid_reg;
  assign line_1453_clock = clock;
  assign line_1453_reset = reset;
  assign line_1453_valid = 2'h3 == deq2_StartIndex ^ line_1453_valid_reg;
  assign line_1454_clock = clock;
  assign line_1454_reset = reset;
  assign line_1454_valid = 2'h0 == deq2_StartIndex ^ line_1454_valid_reg;
  assign line_1455_clock = clock;
  assign line_1455_reset = reset;
  assign line_1455_valid = 2'h1 == deq2_StartIndex ^ line_1455_valid_reg;
  assign line_1456_clock = clock;
  assign line_1456_reset = reset;
  assign line_1456_valid = 2'h2 == deq2_StartIndex ^ line_1456_valid_reg;
  assign line_1457_clock = clock;
  assign line_1457_reset = reset;
  assign line_1457_valid = 2'h3 == deq2_StartIndex ^ line_1457_valid_reg;
  assign line_1458_clock = clock;
  assign line_1458_reset = reset;
  assign line_1458_valid = 2'h0 == deq2_StartIndex ^ line_1458_valid_reg;
  assign line_1459_clock = clock;
  assign line_1459_reset = reset;
  assign line_1459_valid = 2'h1 == deq2_StartIndex ^ line_1459_valid_reg;
  assign line_1460_clock = clock;
  assign line_1460_reset = reset;
  assign line_1460_valid = 2'h2 == deq2_StartIndex ^ line_1460_valid_reg;
  assign line_1461_clock = clock;
  assign line_1461_reset = reset;
  assign line_1461_valid = 2'h3 == deq2_StartIndex ^ line_1461_valid_reg;
  assign line_1462_clock = clock;
  assign line_1462_reset = reset;
  assign line_1462_valid = 2'h0 == deq2_StartIndex ^ line_1462_valid_reg;
  assign line_1463_clock = clock;
  assign line_1463_reset = reset;
  assign line_1463_valid = 2'h1 == deq2_StartIndex ^ line_1463_valid_reg;
  assign line_1464_clock = clock;
  assign line_1464_reset = reset;
  assign line_1464_valid = 2'h2 == deq2_StartIndex ^ line_1464_valid_reg;
  assign line_1465_clock = clock;
  assign line_1465_reset = reset;
  assign line_1465_valid = 2'h3 == deq2_StartIndex ^ line_1465_valid_reg;
  assign line_1466_clock = clock;
  assign line_1466_reset = reset;
  assign line_1466_valid = 2'h0 == deq2_StartIndex ^ line_1466_valid_reg;
  assign line_1467_clock = clock;
  assign line_1467_reset = reset;
  assign line_1467_valid = 2'h1 == deq2_StartIndex ^ line_1467_valid_reg;
  assign line_1468_clock = clock;
  assign line_1468_reset = reset;
  assign line_1468_valid = 2'h2 == deq2_StartIndex ^ line_1468_valid_reg;
  assign line_1469_clock = clock;
  assign line_1469_reset = reset;
  assign line_1469_valid = 2'h3 == deq2_StartIndex ^ line_1469_valid_reg;
  assign line_1470_clock = clock;
  assign line_1470_reset = reset;
  assign line_1470_valid = 2'h0 == deq2_StartIndex ^ line_1470_valid_reg;
  assign line_1471_clock = clock;
  assign line_1471_reset = reset;
  assign line_1471_valid = 2'h1 == deq2_StartIndex ^ line_1471_valid_reg;
  assign line_1472_clock = clock;
  assign line_1472_reset = reset;
  assign line_1472_valid = 2'h2 == deq2_StartIndex ^ line_1472_valid_reg;
  assign line_1473_clock = clock;
  assign line_1473_reset = reset;
  assign line_1473_valid = 2'h3 == deq2_StartIndex ^ line_1473_valid_reg;
  assign line_1474_clock = clock;
  assign line_1474_reset = reset;
  assign line_1474_valid = 2'h0 == deq2_StartIndex ^ line_1474_valid_reg;
  assign line_1475_clock = clock;
  assign line_1475_reset = reset;
  assign line_1475_valid = 2'h1 == deq2_StartIndex ^ line_1475_valid_reg;
  assign line_1476_clock = clock;
  assign line_1476_reset = reset;
  assign line_1476_valid = 2'h2 == deq2_StartIndex ^ line_1476_valid_reg;
  assign line_1477_clock = clock;
  assign line_1477_reset = reset;
  assign line_1477_valid = 2'h3 == deq2_StartIndex ^ line_1477_valid_reg;
  assign line_1478_clock = clock;
  assign line_1478_reset = reset;
  assign line_1478_valid = 2'h0 == deq2_StartIndex ^ line_1478_valid_reg;
  assign line_1479_clock = clock;
  assign line_1479_reset = reset;
  assign line_1479_valid = 2'h1 == deq2_StartIndex ^ line_1479_valid_reg;
  assign line_1480_clock = clock;
  assign line_1480_reset = reset;
  assign line_1480_valid = 2'h2 == deq2_StartIndex ^ line_1480_valid_reg;
  assign line_1481_clock = clock;
  assign line_1481_reset = reset;
  assign line_1481_valid = 2'h3 == deq2_StartIndex ^ line_1481_valid_reg;
  assign line_1482_clock = clock;
  assign line_1482_reset = reset;
  assign line_1482_valid = 2'h0 == deq2_StartIndex ^ line_1482_valid_reg;
  assign line_1483_clock = clock;
  assign line_1483_reset = reset;
  assign line_1483_valid = 2'h1 == deq2_StartIndex ^ line_1483_valid_reg;
  assign line_1484_clock = clock;
  assign line_1484_reset = reset;
  assign line_1484_valid = 2'h2 == deq2_StartIndex ^ line_1484_valid_reg;
  assign line_1485_clock = clock;
  assign line_1485_reset = reset;
  assign line_1485_valid = 2'h3 == deq2_StartIndex ^ line_1485_valid_reg;
  assign line_1486_clock = clock;
  assign line_1486_reset = reset;
  assign line_1486_valid = 2'h0 == deq2_StartIndex ^ line_1486_valid_reg;
  assign line_1487_clock = clock;
  assign line_1487_reset = reset;
  assign line_1487_valid = 2'h1 == deq2_StartIndex ^ line_1487_valid_reg;
  assign line_1488_clock = clock;
  assign line_1488_reset = reset;
  assign line_1488_valid = 2'h2 == deq2_StartIndex ^ line_1488_valid_reg;
  assign line_1489_clock = clock;
  assign line_1489_reset = reset;
  assign line_1489_valid = 2'h3 == deq2_StartIndex ^ line_1489_valid_reg;
  assign line_1490_clock = clock;
  assign line_1490_reset = reset;
  assign line_1490_valid = 2'h0 == deq2_StartIndex ^ line_1490_valid_reg;
  assign line_1491_clock = clock;
  assign line_1491_reset = reset;
  assign line_1491_valid = 2'h1 == deq2_StartIndex ^ line_1491_valid_reg;
  assign line_1492_clock = clock;
  assign line_1492_reset = reset;
  assign line_1492_valid = 2'h2 == deq2_StartIndex ^ line_1492_valid_reg;
  assign line_1493_clock = clock;
  assign line_1493_reset = reset;
  assign line_1493_valid = 2'h3 == deq2_StartIndex ^ line_1493_valid_reg;
  assign line_1494_clock = clock;
  assign line_1494_reset = reset;
  assign line_1494_valid = 2'h0 == deq2_StartIndex ^ line_1494_valid_reg;
  assign line_1495_clock = clock;
  assign line_1495_reset = reset;
  assign line_1495_valid = 2'h1 == deq2_StartIndex ^ line_1495_valid_reg;
  assign line_1496_clock = clock;
  assign line_1496_reset = reset;
  assign line_1496_valid = 2'h2 == deq2_StartIndex ^ line_1496_valid_reg;
  assign line_1497_clock = clock;
  assign line_1497_reset = reset;
  assign line_1497_valid = 2'h3 == deq2_StartIndex ^ line_1497_valid_reg;
  assign line_1498_clock = clock;
  assign line_1498_reset = reset;
  assign line_1498_valid = 2'h0 == deq2_StartIndex ^ line_1498_valid_reg;
  assign line_1499_clock = clock;
  assign line_1499_reset = reset;
  assign line_1499_valid = 2'h1 == deq2_StartIndex ^ line_1499_valid_reg;
  assign line_1500_clock = clock;
  assign line_1500_reset = reset;
  assign line_1500_valid = 2'h2 == deq2_StartIndex ^ line_1500_valid_reg;
  assign line_1501_clock = clock;
  assign line_1501_reset = reset;
  assign line_1501_valid = 2'h3 == deq2_StartIndex ^ line_1501_valid_reg;
  assign line_1502_clock = clock;
  assign line_1502_reset = reset;
  assign line_1502_valid = 2'h0 == deq2_StartIndex ^ line_1502_valid_reg;
  assign line_1503_clock = clock;
  assign line_1503_reset = reset;
  assign line_1503_valid = 2'h1 == deq2_StartIndex ^ line_1503_valid_reg;
  assign line_1504_clock = clock;
  assign line_1504_reset = reset;
  assign line_1504_valid = 2'h2 == deq2_StartIndex ^ line_1504_valid_reg;
  assign line_1505_clock = clock;
  assign line_1505_reset = reset;
  assign line_1505_valid = 2'h3 == deq2_StartIndex ^ line_1505_valid_reg;
  assign line_1506_clock = clock;
  assign line_1506_reset = reset;
  assign line_1506_valid = 2'h0 == deq2_StartIndex ^ line_1506_valid_reg;
  assign line_1507_clock = clock;
  assign line_1507_reset = reset;
  assign line_1507_valid = 2'h1 == deq2_StartIndex ^ line_1507_valid_reg;
  assign line_1508_clock = clock;
  assign line_1508_reset = reset;
  assign line_1508_valid = 2'h2 == deq2_StartIndex ^ line_1508_valid_reg;
  assign line_1509_clock = clock;
  assign line_1509_reset = reset;
  assign line_1509_valid = 2'h3 == deq2_StartIndex ^ line_1509_valid_reg;
  assign line_1510_clock = clock;
  assign line_1510_reset = reset;
  assign line_1510_valid = 2'h0 == deq2_StartIndex ^ line_1510_valid_reg;
  assign line_1511_clock = clock;
  assign line_1511_reset = reset;
  assign line_1511_valid = 2'h1 == deq2_StartIndex ^ line_1511_valid_reg;
  assign line_1512_clock = clock;
  assign line_1512_reset = reset;
  assign line_1512_valid = 2'h2 == deq2_StartIndex ^ line_1512_valid_reg;
  assign line_1513_clock = clock;
  assign line_1513_reset = reset;
  assign line_1513_valid = 2'h3 == deq2_StartIndex ^ line_1513_valid_reg;
  assign line_1514_clock = clock;
  assign line_1514_reset = reset;
  assign line_1514_valid = 2'h0 == deq2_StartIndex ^ line_1514_valid_reg;
  assign line_1515_clock = clock;
  assign line_1515_reset = reset;
  assign line_1515_valid = 2'h1 == deq2_StartIndex ^ line_1515_valid_reg;
  assign line_1516_clock = clock;
  assign line_1516_reset = reset;
  assign line_1516_valid = 2'h2 == deq2_StartIndex ^ line_1516_valid_reg;
  assign line_1517_clock = clock;
  assign line_1517_reset = reset;
  assign line_1517_valid = 2'h3 == deq2_StartIndex ^ line_1517_valid_reg;
  assign line_1518_clock = clock;
  assign line_1518_reset = reset;
  assign line_1518_valid = 2'h0 == deq2_StartIndex ^ line_1518_valid_reg;
  assign line_1519_clock = clock;
  assign line_1519_reset = reset;
  assign line_1519_valid = 2'h1 == deq2_StartIndex ^ line_1519_valid_reg;
  assign line_1520_clock = clock;
  assign line_1520_reset = reset;
  assign line_1520_valid = 2'h2 == deq2_StartIndex ^ line_1520_valid_reg;
  assign line_1521_clock = clock;
  assign line_1521_reset = reset;
  assign line_1521_valid = 2'h3 == deq2_StartIndex ^ line_1521_valid_reg;
  assign line_1522_clock = clock;
  assign line_1522_reset = reset;
  assign line_1522_valid = 2'h0 == deq2_StartIndex ^ line_1522_valid_reg;
  assign line_1523_clock = clock;
  assign line_1523_reset = reset;
  assign line_1523_valid = 2'h1 == deq2_StartIndex ^ line_1523_valid_reg;
  assign line_1524_clock = clock;
  assign line_1524_reset = reset;
  assign line_1524_valid = 2'h2 == deq2_StartIndex ^ line_1524_valid_reg;
  assign line_1525_clock = clock;
  assign line_1525_reset = reset;
  assign line_1525_valid = 2'h3 == deq2_StartIndex ^ line_1525_valid_reg;
  assign line_1526_clock = clock;
  assign line_1526_reset = reset;
  assign line_1526_valid = 2'h0 == deq2_StartIndex ^ line_1526_valid_reg;
  assign line_1527_clock = clock;
  assign line_1527_reset = reset;
  assign line_1527_valid = 2'h1 == deq2_StartIndex ^ line_1527_valid_reg;
  assign line_1528_clock = clock;
  assign line_1528_reset = reset;
  assign line_1528_valid = 2'h2 == deq2_StartIndex ^ line_1528_valid_reg;
  assign line_1529_clock = clock;
  assign line_1529_reset = reset;
  assign line_1529_valid = 2'h3 == deq2_StartIndex ^ line_1529_valid_reg;
  assign line_1530_clock = clock;
  assign line_1530_reset = reset;
  assign line_1530_valid = 2'h0 == deq2_StartIndex ^ line_1530_valid_reg;
  assign line_1531_clock = clock;
  assign line_1531_reset = reset;
  assign line_1531_valid = 2'h1 == deq2_StartIndex ^ line_1531_valid_reg;
  assign line_1532_clock = clock;
  assign line_1532_reset = reset;
  assign line_1532_valid = 2'h2 == deq2_StartIndex ^ line_1532_valid_reg;
  assign line_1533_clock = clock;
  assign line_1533_reset = reset;
  assign line_1533_valid = 2'h3 == deq2_StartIndex ^ line_1533_valid_reg;
  assign line_1534_clock = clock;
  assign line_1534_reset = reset;
  assign line_1534_valid = 2'h0 == deq2_StartIndex ^ line_1534_valid_reg;
  assign line_1535_clock = clock;
  assign line_1535_reset = reset;
  assign line_1535_valid = 2'h1 == deq2_StartIndex ^ line_1535_valid_reg;
  assign line_1536_clock = clock;
  assign line_1536_reset = reset;
  assign line_1536_valid = 2'h2 == deq2_StartIndex ^ line_1536_valid_reg;
  assign line_1537_clock = clock;
  assign line_1537_reset = reset;
  assign line_1537_valid = 2'h3 == deq2_StartIndex ^ line_1537_valid_reg;
  assign line_1538_clock = clock;
  assign line_1538_reset = reset;
  assign line_1538_valid = 2'h0 == deq2_StartIndex ^ line_1538_valid_reg;
  assign line_1539_clock = clock;
  assign line_1539_reset = reset;
  assign line_1539_valid = 2'h1 == deq2_StartIndex ^ line_1539_valid_reg;
  assign line_1540_clock = clock;
  assign line_1540_reset = reset;
  assign line_1540_valid = 2'h2 == deq2_StartIndex ^ line_1540_valid_reg;
  assign line_1541_clock = clock;
  assign line_1541_reset = reset;
  assign line_1541_valid = 2'h3 == deq2_StartIndex ^ line_1541_valid_reg;
  assign line_1542_clock = clock;
  assign line_1542_reset = reset;
  assign line_1542_valid = 2'h0 == deq2_StartIndex ^ line_1542_valid_reg;
  assign line_1543_clock = clock;
  assign line_1543_reset = reset;
  assign line_1543_valid = 2'h1 == deq2_StartIndex ^ line_1543_valid_reg;
  assign line_1544_clock = clock;
  assign line_1544_reset = reset;
  assign line_1544_valid = 2'h2 == deq2_StartIndex ^ line_1544_valid_reg;
  assign line_1545_clock = clock;
  assign line_1545_reset = reset;
  assign line_1545_valid = 2'h3 == deq2_StartIndex ^ line_1545_valid_reg;
  assign line_1546_clock = clock;
  assign line_1546_reset = reset;
  assign line_1546_valid = 2'h0 == deq2_StartIndex ^ line_1546_valid_reg;
  assign line_1547_clock = clock;
  assign line_1547_reset = reset;
  assign line_1547_valid = 2'h1 == deq2_StartIndex ^ line_1547_valid_reg;
  assign line_1548_clock = clock;
  assign line_1548_reset = reset;
  assign line_1548_valid = 2'h2 == deq2_StartIndex ^ line_1548_valid_reg;
  assign line_1549_clock = clock;
  assign line_1549_reset = reset;
  assign line_1549_valid = 2'h3 == deq2_StartIndex ^ line_1549_valid_reg;
  assign line_1550_clock = clock;
  assign line_1550_reset = reset;
  assign line_1550_valid = 2'h0 == deq2_StartIndex ^ line_1550_valid_reg;
  assign line_1551_clock = clock;
  assign line_1551_reset = reset;
  assign line_1551_valid = 2'h1 == deq2_StartIndex ^ line_1551_valid_reg;
  assign line_1552_clock = clock;
  assign line_1552_reset = reset;
  assign line_1552_valid = 2'h2 == deq2_StartIndex ^ line_1552_valid_reg;
  assign line_1553_clock = clock;
  assign line_1553_reset = reset;
  assign line_1553_valid = 2'h3 == deq2_StartIndex ^ line_1553_valid_reg;
  assign line_1554_clock = clock;
  assign line_1554_reset = reset;
  assign line_1554_valid = 2'h0 == deq2_StartIndex ^ line_1554_valid_reg;
  assign line_1555_clock = clock;
  assign line_1555_reset = reset;
  assign line_1555_valid = 2'h1 == deq2_StartIndex ^ line_1555_valid_reg;
  assign line_1556_clock = clock;
  assign line_1556_reset = reset;
  assign line_1556_valid = 2'h2 == deq2_StartIndex ^ line_1556_valid_reg;
  assign line_1557_clock = clock;
  assign line_1557_reset = reset;
  assign line_1557_valid = 2'h3 == deq2_StartIndex ^ line_1557_valid_reg;
  assign line_1558_clock = clock;
  assign line_1558_reset = reset;
  assign line_1558_valid = 2'h0 == deq2_StartIndex ^ line_1558_valid_reg;
  assign line_1559_clock = clock;
  assign line_1559_reset = reset;
  assign line_1559_valid = 2'h1 == deq2_StartIndex ^ line_1559_valid_reg;
  assign line_1560_clock = clock;
  assign line_1560_reset = reset;
  assign line_1560_valid = 2'h2 == deq2_StartIndex ^ line_1560_valid_reg;
  assign line_1561_clock = clock;
  assign line_1561_reset = reset;
  assign line_1561_valid = 2'h3 == deq2_StartIndex ^ line_1561_valid_reg;
  assign line_1562_clock = clock;
  assign line_1562_reset = reset;
  assign line_1562_valid = 2'h0 == deq2_StartIndex ^ line_1562_valid_reg;
  assign line_1563_clock = clock;
  assign line_1563_reset = reset;
  assign line_1563_valid = 2'h1 == deq2_StartIndex ^ line_1563_valid_reg;
  assign line_1564_clock = clock;
  assign line_1564_reset = reset;
  assign line_1564_valid = 2'h2 == deq2_StartIndex ^ line_1564_valid_reg;
  assign line_1565_clock = clock;
  assign line_1565_reset = reset;
  assign line_1565_valid = 2'h3 == deq2_StartIndex ^ line_1565_valid_reg;
  assign line_1566_clock = clock;
  assign line_1566_reset = reset;
  assign line_1566_valid = 2'h0 == deq2_StartIndex ^ line_1566_valid_reg;
  assign line_1567_clock = clock;
  assign line_1567_reset = reset;
  assign line_1567_valid = 2'h1 == deq2_StartIndex ^ line_1567_valid_reg;
  assign line_1568_clock = clock;
  assign line_1568_reset = reset;
  assign line_1568_valid = 2'h2 == deq2_StartIndex ^ line_1568_valid_reg;
  assign line_1569_clock = clock;
  assign line_1569_reset = reset;
  assign line_1569_valid = 2'h3 == deq2_StartIndex ^ line_1569_valid_reg;
  assign line_1570_clock = clock;
  assign line_1570_reset = reset;
  assign line_1570_valid = 2'h0 == deq2_StartIndex ^ line_1570_valid_reg;
  assign line_1571_clock = clock;
  assign line_1571_reset = reset;
  assign line_1571_valid = 2'h1 == deq2_StartIndex ^ line_1571_valid_reg;
  assign line_1572_clock = clock;
  assign line_1572_reset = reset;
  assign line_1572_valid = 2'h2 == deq2_StartIndex ^ line_1572_valid_reg;
  assign line_1573_clock = clock;
  assign line_1573_reset = reset;
  assign line_1573_valid = 2'h3 == deq2_StartIndex ^ line_1573_valid_reg;
  assign line_1574_clock = clock;
  assign line_1574_reset = reset;
  assign line_1574_valid = 2'h0 == deq2_StartIndex ^ line_1574_valid_reg;
  assign line_1575_clock = clock;
  assign line_1575_reset = reset;
  assign line_1575_valid = 2'h1 == deq2_StartIndex ^ line_1575_valid_reg;
  assign line_1576_clock = clock;
  assign line_1576_reset = reset;
  assign line_1576_valid = 2'h2 == deq2_StartIndex ^ line_1576_valid_reg;
  assign line_1577_clock = clock;
  assign line_1577_reset = reset;
  assign line_1577_valid = 2'h3 == deq2_StartIndex ^ line_1577_valid_reg;
  assign line_1578_clock = clock;
  assign line_1578_reset = reset;
  assign line_1578_valid = 2'h0 == deq2_StartIndex ^ line_1578_valid_reg;
  assign line_1579_clock = clock;
  assign line_1579_reset = reset;
  assign line_1579_valid = 2'h1 == deq2_StartIndex ^ line_1579_valid_reg;
  assign line_1580_clock = clock;
  assign line_1580_reset = reset;
  assign line_1580_valid = 2'h2 == deq2_StartIndex ^ line_1580_valid_reg;
  assign line_1581_clock = clock;
  assign line_1581_reset = reset;
  assign line_1581_valid = 2'h3 == deq2_StartIndex ^ line_1581_valid_reg;
  assign line_1582_clock = clock;
  assign line_1582_reset = reset;
  assign line_1582_valid = 2'h0 == deq2_StartIndex ^ line_1582_valid_reg;
  assign line_1583_clock = clock;
  assign line_1583_reset = reset;
  assign line_1583_valid = 2'h1 == deq2_StartIndex ^ line_1583_valid_reg;
  assign line_1584_clock = clock;
  assign line_1584_reset = reset;
  assign line_1584_valid = 2'h2 == deq2_StartIndex ^ line_1584_valid_reg;
  assign line_1585_clock = clock;
  assign line_1585_reset = reset;
  assign line_1585_valid = 2'h3 == deq2_StartIndex ^ line_1585_valid_reg;
  assign line_1586_clock = clock;
  assign line_1586_reset = reset;
  assign line_1586_valid = 2'h0 == deq2_StartIndex ^ line_1586_valid_reg;
  assign line_1587_clock = clock;
  assign line_1587_reset = reset;
  assign line_1587_valid = 2'h1 == deq2_StartIndex ^ line_1587_valid_reg;
  assign line_1588_clock = clock;
  assign line_1588_reset = reset;
  assign line_1588_valid = 2'h2 == deq2_StartIndex ^ line_1588_valid_reg;
  assign line_1589_clock = clock;
  assign line_1589_reset = reset;
  assign line_1589_valid = 2'h3 == deq2_StartIndex ^ line_1589_valid_reg;
  assign line_1590_clock = clock;
  assign line_1590_reset = reset;
  assign line_1590_valid = 2'h0 == deq2_StartIndex ^ line_1590_valid_reg;
  assign line_1591_clock = clock;
  assign line_1591_reset = reset;
  assign line_1591_valid = 2'h1 == deq2_StartIndex ^ line_1591_valid_reg;
  assign line_1592_clock = clock;
  assign line_1592_reset = reset;
  assign line_1592_valid = 2'h2 == deq2_StartIndex ^ line_1592_valid_reg;
  assign line_1593_clock = clock;
  assign line_1593_reset = reset;
  assign line_1593_valid = 2'h3 == deq2_StartIndex ^ line_1593_valid_reg;
  assign line_1594_clock = clock;
  assign line_1594_reset = reset;
  assign line_1594_valid = 2'h0 == deq2_StartIndex ^ line_1594_valid_reg;
  assign line_1595_clock = clock;
  assign line_1595_reset = reset;
  assign line_1595_valid = 2'h1 == deq2_StartIndex ^ line_1595_valid_reg;
  assign line_1596_clock = clock;
  assign line_1596_reset = reset;
  assign line_1596_valid = 2'h2 == deq2_StartIndex ^ line_1596_valid_reg;
  assign line_1597_clock = clock;
  assign line_1597_reset = reset;
  assign line_1597_valid = 2'h3 == deq2_StartIndex ^ line_1597_valid_reg;
  assign line_1598_clock = clock;
  assign line_1598_reset = reset;
  assign line_1598_valid = 2'h0 == deq2_StartIndex ^ line_1598_valid_reg;
  assign line_1599_clock = clock;
  assign line_1599_reset = reset;
  assign line_1599_valid = 2'h1 == deq2_StartIndex ^ line_1599_valid_reg;
  assign line_1600_clock = clock;
  assign line_1600_reset = reset;
  assign line_1600_valid = 2'h2 == deq2_StartIndex ^ line_1600_valid_reg;
  assign line_1601_clock = clock;
  assign line_1601_reset = reset;
  assign line_1601_valid = 2'h3 == deq2_StartIndex ^ line_1601_valid_reg;
  assign line_1602_clock = clock;
  assign line_1602_reset = reset;
  assign line_1602_valid = 2'h0 == deq2_StartIndex ^ line_1602_valid_reg;
  assign line_1603_clock = clock;
  assign line_1603_reset = reset;
  assign line_1603_valid = 2'h1 == deq2_StartIndex ^ line_1603_valid_reg;
  assign line_1604_clock = clock;
  assign line_1604_reset = reset;
  assign line_1604_valid = 2'h2 == deq2_StartIndex ^ line_1604_valid_reg;
  assign line_1605_clock = clock;
  assign line_1605_reset = reset;
  assign line_1605_valid = 2'h3 == deq2_StartIndex ^ line_1605_valid_reg;
  assign line_1606_clock = clock;
  assign line_1606_reset = reset;
  assign line_1606_valid = 2'h0 == deq2_StartIndex ^ line_1606_valid_reg;
  assign line_1607_clock = clock;
  assign line_1607_reset = reset;
  assign line_1607_valid = 2'h1 == deq2_StartIndex ^ line_1607_valid_reg;
  assign line_1608_clock = clock;
  assign line_1608_reset = reset;
  assign line_1608_valid = 2'h2 == deq2_StartIndex ^ line_1608_valid_reg;
  assign line_1609_clock = clock;
  assign line_1609_reset = reset;
  assign line_1609_valid = 2'h3 == deq2_StartIndex ^ line_1609_valid_reg;
  assign line_1610_clock = clock;
  assign line_1610_reset = reset;
  assign line_1610_valid = 2'h0 == deq2_StartIndex ^ line_1610_valid_reg;
  assign line_1611_clock = clock;
  assign line_1611_reset = reset;
  assign line_1611_valid = 2'h1 == deq2_StartIndex ^ line_1611_valid_reg;
  assign line_1612_clock = clock;
  assign line_1612_reset = reset;
  assign line_1612_valid = 2'h2 == deq2_StartIndex ^ line_1612_valid_reg;
  assign line_1613_clock = clock;
  assign line_1613_reset = reset;
  assign line_1613_valid = 2'h3 == deq2_StartIndex ^ line_1613_valid_reg;
  assign line_1614_clock = clock;
  assign line_1614_reset = reset;
  assign line_1614_valid = 2'h0 == deq2_StartIndex ^ line_1614_valid_reg;
  assign line_1615_clock = clock;
  assign line_1615_reset = reset;
  assign line_1615_valid = 2'h1 == deq2_StartIndex ^ line_1615_valid_reg;
  assign line_1616_clock = clock;
  assign line_1616_reset = reset;
  assign line_1616_valid = 2'h2 == deq2_StartIndex ^ line_1616_valid_reg;
  assign line_1617_clock = clock;
  assign line_1617_reset = reset;
  assign line_1617_valid = 2'h3 == deq2_StartIndex ^ line_1617_valid_reg;
  assign line_1618_clock = clock;
  assign line_1618_reset = reset;
  assign line_1618_valid = 2'h0 == deq2_StartIndex ^ line_1618_valid_reg;
  assign line_1619_clock = clock;
  assign line_1619_reset = reset;
  assign line_1619_valid = 2'h1 == deq2_StartIndex ^ line_1619_valid_reg;
  assign line_1620_clock = clock;
  assign line_1620_reset = reset;
  assign line_1620_valid = 2'h2 == deq2_StartIndex ^ line_1620_valid_reg;
  assign line_1621_clock = clock;
  assign line_1621_reset = reset;
  assign line_1621_valid = 2'h3 == deq2_StartIndex ^ line_1621_valid_reg;
  assign line_1622_clock = clock;
  assign line_1622_reset = reset;
  assign line_1622_valid = 2'h0 == deq2_StartIndex ^ line_1622_valid_reg;
  assign line_1623_clock = clock;
  assign line_1623_reset = reset;
  assign line_1623_valid = 2'h1 == deq2_StartIndex ^ line_1623_valid_reg;
  assign line_1624_clock = clock;
  assign line_1624_reset = reset;
  assign line_1624_valid = 2'h2 == deq2_StartIndex ^ line_1624_valid_reg;
  assign line_1625_clock = clock;
  assign line_1625_reset = reset;
  assign line_1625_valid = 2'h3 == deq2_StartIndex ^ line_1625_valid_reg;
  assign line_1626_clock = clock;
  assign line_1626_reset = reset;
  assign line_1626_valid = dequeueFire ^ line_1626_valid_reg;
  assign line_1627_clock = clock;
  assign line_1627_reset = reset;
  assign line_1627_valid = frontend_io_flushVec[1] ^ line_1627_valid_reg;
  assign io_imem_mem_req_valid = io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_mem_req_bits_addr = io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_dmem_mem_req_valid = io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_addr = io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_size = io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_cmd = io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wmask = io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wdata = io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_frontend_req_ready = dmemXbar_io_in_3_req_ready; // @[src/main/scala/nutcore/NutCore.scala 222:23]
  assign isWFI = frontend_isWFI;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_out_0_ready = ringBufferAllowin | ~frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_iaf = itlb_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 189:21]
  assign frontend_io_sfence_vma_invalid = backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 215:36]
  assign frontend_io_wfi_invalid = backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 216:29]
  assign frontend_REG_valid = backend_REG_valid;
  assign frontend_REG_pc = backend_REG_pc;
  assign frontend_REG_isMissPredict = backend_REG_isMissPredict;
  assign frontend_REG_actualTarget = backend_REG_actualTarget;
  assign frontend_REG_actualTaken = backend_REG_actualTaken;
  assign frontend_REG_fuOpType = backend_REG_fuOpType;
  assign frontend_REG_btbType = backend_REG_btbType;
  assign frontend_REG_isRVC = backend_REG_isRVC;
  assign frontend_flushICache = backend_flushICache;
  assign frontend_flushTLB = backend_flushTLB;
  assign frontend_intrVecIDU = backend_intrVecIDU;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = ringBufferHead != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 2'h3 == ringBufferTail ? dataBuffer_3_cf_instr : _GEN_2244; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pc : _GEN_2240; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pnpc : _GEN_2236; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_1 : _GEN_2164; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_2 : _GEN_2168; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_12 : _GEN_2208; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_1 : _GEN_2116; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_3 : _GEN_2124; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_5 : _GEN_2132; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_7 : _GEN_2140; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_9 : _GEN_2148; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_11 : _GEN_2156; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 2'h3 == ringBufferTail ? dataBuffer_3_cf_brIdx : _GEN_2108; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_crossBoundaryFault = 2'h3 == ringBufferTail ? dataBuffer_3_cf_crossBoundaryFault :
    _GEN_2100; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src1Type : _GEN_2084; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src2Type : _GEN_2080; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuType : _GEN_2076; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuOpType : _GEN_2072; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc1 : _GEN_2068; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc2 : _GEN_2064; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfWen : _GEN_2060; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfDest : _GEN_2056; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_isNutCoreTrap = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_isNutCoreTrap : _GEN_2052; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 2'h3 == ringBufferTail ? dataBuffer_3_data_imm : _GEN_2024; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[src/main/scala/nutcore/NutCore.scala 219:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_memMMU_dmem_loadPF = dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_storePF = dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_laf = dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_saf = dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_extra_meip_0 = io_extra_meip_0;
  assign backend_paddr = dtlb_paddr;
  assign backend__T_12 = dtlb__T_12_0;
  assign backend_scIsSuccess = dtlb_scIsSuccess_0;
  assign backend_io_extra_mtip = io_extra_mtip;
  assign backend_vmEnable = dtlb_vmEnable_0;
  assign backend_tlbFinish = dtlb_tlbFinish_0;
  assign backend_ismmio = io_dmem_cache_ismmio_0;
  assign backend__T_13_0 = dtlb__T_13_1;
  assign backend_io_extra_msip = io_extra_msip;
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_0_req_bits_addr = io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_valid = io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_addr = io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_cmd = io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wmask = io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wdata = io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_1_req_valid = filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_addr = filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_cmd = filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_wdata = filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_valid = filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_addr = filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_cmd = filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_wdata = filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_out_req_ready = io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_valid = io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_cmd = io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_rdata = io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_out_req_ready = io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_valid = io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_rdata = io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_user = io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_mem_req_ready = filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_valid = filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_bits_rdata = filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_flush = frontend_io_flushVec[0]; // @[src/main/scala/nutcore/NutCore.scala 184:35]
  assign itlb_io_csrMMU_priviledgeMode = backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign itlb_CSRSATP = backend_satp;
  assign itlb_MOUFlushTLB = backend_flushTLB;
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_in_req_valid = itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_addr = itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_cmd = itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_wdata = itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_out_req_ready = dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_valid = dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_bits_rdata = dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_u = backend_io_memMMU_imem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_imem_cache_clock = clock;
  assign io_imem_cache_reset = reset;
  assign io_imem_cache_io_in_req_valid = itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/NutCore.scala 193:19]
  assign io_imem_cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign dtlb_clock = clock;
  assign dtlb_reset = reset;
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_mem_req_ready = filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_valid = filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_bits_rdata = filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_csrMMU_priviledgeMode = backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_sum = backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_mxr = backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_lr = backend_lr;
  assign dtlb_scInflight = backend_scInflight;
  assign dtlb_amoReq = backend_amoReq;
  assign dtlb_lrAddr = backend_lrAddr;
  assign dtlb_CSRSATP = backend_satp;
  assign dtlb_MOUFlushTLB = backend_flushTLB;
  assign filter_1_clock = clock;
  assign filter_1_reset = reset;
  assign filter_1_io_in_req_valid = dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_addr = dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_cmd = dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_wdata = dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_out_req_ready = dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_valid = dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_bits_rdata = dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_u = backend_io_memMMU_dmem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_dmem_cache_clock = clock;
  assign io_dmem_cache_reset = reset;
  assign io_dmem_cache_io_in_req_valid = dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_cmd = mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_instr <= _GEN_1125;
        end
      end else begin
        dataBuffer_0_cf_instr <= _GEN_1125;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pc <= _GEN_1129;
        end
      end else begin
        dataBuffer_0_cf_pc <= _GEN_1129;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pnpc <= _GEN_1133;
        end
      end else begin
        dataBuffer_0_cf_pnpc <= _GEN_1133;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_1 <= _GEN_1153;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_1 <= _GEN_1153;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_2 <= _GEN_1157;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_2 <= _GEN_1157;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_12 <= _GEN_1197;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_12 <= _GEN_1197;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_1 <= _GEN_1217;
        end
      end else begin
        dataBuffer_0_cf_intrVec_1 <= _GEN_1217;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_3 <= _GEN_1225;
        end
      end else begin
        dataBuffer_0_cf_intrVec_3 <= _GEN_1225;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_5 <= _GEN_1233;
        end
      end else begin
        dataBuffer_0_cf_intrVec_5 <= _GEN_1233;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_7 <= _GEN_1241;
        end
      end else begin
        dataBuffer_0_cf_intrVec_7 <= _GEN_1241;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_9 <= _GEN_1249;
        end
      end else begin
        dataBuffer_0_cf_intrVec_9 <= _GEN_1249;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_11 <= _GEN_1257;
        end
      end else begin
        dataBuffer_0_cf_intrVec_11 <= _GEN_1257;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_brIdx <= _GEN_1261;
        end
      end else begin
        dataBuffer_0_cf_brIdx <= _GEN_1261;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_crossBoundaryFault <= _GEN_1269;
        end
      end else begin
        dataBuffer_0_cf_crossBoundaryFault <= _GEN_1269;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src1Type <= _GEN_1285;
        end
      end else begin
        dataBuffer_0_ctrl_src1Type <= _GEN_1285;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src2Type <= _GEN_1289;
        end
      end else begin
        dataBuffer_0_ctrl_src2Type <= _GEN_1289;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuType <= _GEN_1293;
        end
      end else begin
        dataBuffer_0_ctrl_fuType <= _GEN_1293;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuOpType <= _GEN_1297;
        end
      end else begin
        dataBuffer_0_ctrl_fuOpType <= _GEN_1297;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc1 <= _GEN_1301;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc1 <= _GEN_1301;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc2 <= _GEN_1305;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc2 <= _GEN_1305;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfWen <= _GEN_1309;
        end
      end else begin
        dataBuffer_0_ctrl_rfWen <= _GEN_1309;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfDest <= _GEN_1313;
        end
      end else begin
        dataBuffer_0_ctrl_rfDest <= _GEN_1313;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_1317;
        end
      end else begin
        dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_1317;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_data_imm <= _GEN_1345;
        end
      end else begin
        dataBuffer_0_data_imm <= _GEN_1345;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_instr <= _GEN_1126;
        end
      end else begin
        dataBuffer_1_cf_instr <= _GEN_1126;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pc <= _GEN_1130;
        end
      end else begin
        dataBuffer_1_cf_pc <= _GEN_1130;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pnpc <= _GEN_1134;
        end
      end else begin
        dataBuffer_1_cf_pnpc <= _GEN_1134;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_1 <= _GEN_1154;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_1 <= _GEN_1154;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_2 <= _GEN_1158;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_2 <= _GEN_1158;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_12 <= _GEN_1198;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_12 <= _GEN_1198;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_1 <= _GEN_1218;
        end
      end else begin
        dataBuffer_1_cf_intrVec_1 <= _GEN_1218;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_3 <= _GEN_1226;
        end
      end else begin
        dataBuffer_1_cf_intrVec_3 <= _GEN_1226;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_5 <= _GEN_1234;
        end
      end else begin
        dataBuffer_1_cf_intrVec_5 <= _GEN_1234;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_7 <= _GEN_1242;
        end
      end else begin
        dataBuffer_1_cf_intrVec_7 <= _GEN_1242;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_9 <= _GEN_1250;
        end
      end else begin
        dataBuffer_1_cf_intrVec_9 <= _GEN_1250;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_11 <= _GEN_1258;
        end
      end else begin
        dataBuffer_1_cf_intrVec_11 <= _GEN_1258;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_brIdx <= _GEN_1262;
        end
      end else begin
        dataBuffer_1_cf_brIdx <= _GEN_1262;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_crossBoundaryFault <= _GEN_1270;
        end
      end else begin
        dataBuffer_1_cf_crossBoundaryFault <= _GEN_1270;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src1Type <= _GEN_1286;
        end
      end else begin
        dataBuffer_1_ctrl_src1Type <= _GEN_1286;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src2Type <= _GEN_1290;
        end
      end else begin
        dataBuffer_1_ctrl_src2Type <= _GEN_1290;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuType <= _GEN_1294;
        end
      end else begin
        dataBuffer_1_ctrl_fuType <= _GEN_1294;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuOpType <= _GEN_1298;
        end
      end else begin
        dataBuffer_1_ctrl_fuOpType <= _GEN_1298;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc1 <= _GEN_1302;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc1 <= _GEN_1302;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc2 <= _GEN_1306;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc2 <= _GEN_1306;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfWen <= _GEN_1310;
        end
      end else begin
        dataBuffer_1_ctrl_rfWen <= _GEN_1310;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfDest <= _GEN_1314;
        end
      end else begin
        dataBuffer_1_ctrl_rfDest <= _GEN_1314;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_1318;
        end
      end else begin
        dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_1318;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_data_imm <= _GEN_1346;
        end
      end else begin
        dataBuffer_1_data_imm <= _GEN_1346;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_instr <= _GEN_1127;
        end
      end else begin
        dataBuffer_2_cf_instr <= _GEN_1127;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pc <= _GEN_1131;
        end
      end else begin
        dataBuffer_2_cf_pc <= _GEN_1131;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pnpc <= _GEN_1135;
        end
      end else begin
        dataBuffer_2_cf_pnpc <= _GEN_1135;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_1 <= _GEN_1155;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_1 <= _GEN_1155;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_2 <= _GEN_1159;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_2 <= _GEN_1159;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_12 <= _GEN_1199;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_12 <= _GEN_1199;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_1 <= _GEN_1219;
        end
      end else begin
        dataBuffer_2_cf_intrVec_1 <= _GEN_1219;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_3 <= _GEN_1227;
        end
      end else begin
        dataBuffer_2_cf_intrVec_3 <= _GEN_1227;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_5 <= _GEN_1235;
        end
      end else begin
        dataBuffer_2_cf_intrVec_5 <= _GEN_1235;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_7 <= _GEN_1243;
        end
      end else begin
        dataBuffer_2_cf_intrVec_7 <= _GEN_1243;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_9 <= _GEN_1251;
        end
      end else begin
        dataBuffer_2_cf_intrVec_9 <= _GEN_1251;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_11 <= _GEN_1259;
        end
      end else begin
        dataBuffer_2_cf_intrVec_11 <= _GEN_1259;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_brIdx <= _GEN_1263;
        end
      end else begin
        dataBuffer_2_cf_brIdx <= _GEN_1263;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_crossBoundaryFault <= _GEN_1271;
        end
      end else begin
        dataBuffer_2_cf_crossBoundaryFault <= _GEN_1271;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src1Type <= _GEN_1287;
        end
      end else begin
        dataBuffer_2_ctrl_src1Type <= _GEN_1287;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src2Type <= _GEN_1291;
        end
      end else begin
        dataBuffer_2_ctrl_src2Type <= _GEN_1291;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuType <= _GEN_1295;
        end
      end else begin
        dataBuffer_2_ctrl_fuType <= _GEN_1295;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuOpType <= _GEN_1299;
        end
      end else begin
        dataBuffer_2_ctrl_fuOpType <= _GEN_1299;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc1 <= _GEN_1303;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc1 <= _GEN_1303;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc2 <= _GEN_1307;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc2 <= _GEN_1307;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfWen <= _GEN_1311;
        end
      end else begin
        dataBuffer_2_ctrl_rfWen <= _GEN_1311;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfDest <= _GEN_1315;
        end
      end else begin
        dataBuffer_2_ctrl_rfDest <= _GEN_1315;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_1319;
        end
      end else begin
        dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_1319;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_data_imm <= _GEN_1347;
        end
      end else begin
        dataBuffer_2_data_imm <= _GEN_1347;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_instr <= _GEN_1128;
        end
      end else begin
        dataBuffer_3_cf_instr <= _GEN_1128;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pc <= _GEN_1132;
        end
      end else begin
        dataBuffer_3_cf_pc <= _GEN_1132;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pnpc <= _GEN_1136;
        end
      end else begin
        dataBuffer_3_cf_pnpc <= _GEN_1136;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_1 <= _GEN_1156;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_1 <= _GEN_1156;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_2 <= _GEN_1160;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_2 <= _GEN_1160;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_12 <= _GEN_1200;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_12 <= _GEN_1200;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_1 <= _GEN_1220;
        end
      end else begin
        dataBuffer_3_cf_intrVec_1 <= _GEN_1220;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_3 <= _GEN_1228;
        end
      end else begin
        dataBuffer_3_cf_intrVec_3 <= _GEN_1228;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_5 <= _GEN_1236;
        end
      end else begin
        dataBuffer_3_cf_intrVec_5 <= _GEN_1236;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_7 <= _GEN_1244;
        end
      end else begin
        dataBuffer_3_cf_intrVec_7 <= _GEN_1244;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_9 <= _GEN_1252;
        end
      end else begin
        dataBuffer_3_cf_intrVec_9 <= _GEN_1252;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_11 <= _GEN_1260;
        end
      end else begin
        dataBuffer_3_cf_intrVec_11 <= _GEN_1260;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_brIdx <= _GEN_1264;
        end
      end else begin
        dataBuffer_3_cf_brIdx <= _GEN_1264;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_crossBoundaryFault <= _GEN_1272;
        end
      end else begin
        dataBuffer_3_cf_crossBoundaryFault <= _GEN_1272;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src1Type <= _GEN_1288;
        end
      end else begin
        dataBuffer_3_ctrl_src1Type <= _GEN_1288;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src2Type <= _GEN_1292;
        end
      end else begin
        dataBuffer_3_ctrl_src2Type <= _GEN_1292;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuType <= _GEN_1296;
        end
      end else begin
        dataBuffer_3_ctrl_fuType <= _GEN_1296;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuOpType <= _GEN_1300;
        end
      end else begin
        dataBuffer_3_ctrl_fuOpType <= _GEN_1300;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc1 <= _GEN_1304;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc1 <= _GEN_1304;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc2 <= _GEN_1308;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc2 <= _GEN_1308;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfWen <= _GEN_1312;
        end
      end else begin
        dataBuffer_3_ctrl_rfWen <= _GEN_1312;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfDest <= _GEN_1316;
        end
      end else begin
        dataBuffer_3_ctrl_rfDest <= _GEN_1316;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_1320;
        end
      end else begin
        dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_1320;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_data_imm <= _GEN_1348;
        end
      end else begin
        dataBuffer_3_data_imm <= _GEN_1348;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 30:33]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 72:24]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      ringBufferHead <= _ringBufferHead_T_1; // @[src/main/scala/utils/PipelineVector.scala 47:24]
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 31:33]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 73:24]
    end else if (dequeueFire) begin // @[src/main/scala/utils/PipelineVector.scala 66:22]
      ringBufferTail <= _ringBufferTail_T_1; // @[src/main/scala/utils/PipelineVector.scala 67:24]
    end
    line_727_valid_reg <= wen;
    line_728_valid_reg <= enqueueFire_0;
    line_729_valid_reg <= 2'h0 == _T_1[1:0];
    line_730_valid_reg <= 2'h1 == _T_1[1:0];
    line_731_valid_reg <= 2'h2 == _T_1[1:0];
    line_732_valid_reg <= 2'h3 == _T_1[1:0];
    line_733_valid_reg <= 2'h0 == _T_1[1:0];
    line_734_valid_reg <= 2'h1 == _T_1[1:0];
    line_735_valid_reg <= 2'h2 == _T_1[1:0];
    line_736_valid_reg <= 2'h3 == _T_1[1:0];
    line_737_valid_reg <= 2'h0 == _T_1[1:0];
    line_738_valid_reg <= 2'h1 == _T_1[1:0];
    line_739_valid_reg <= 2'h2 == _T_1[1:0];
    line_740_valid_reg <= 2'h3 == _T_1[1:0];
    line_741_valid_reg <= 2'h0 == _T_1[1:0];
    line_742_valid_reg <= 2'h1 == _T_1[1:0];
    line_743_valid_reg <= 2'h2 == _T_1[1:0];
    line_744_valid_reg <= 2'h3 == _T_1[1:0];
    line_745_valid_reg <= 2'h0 == _T_1[1:0];
    line_746_valid_reg <= 2'h1 == _T_1[1:0];
    line_747_valid_reg <= 2'h2 == _T_1[1:0];
    line_748_valid_reg <= 2'h3 == _T_1[1:0];
    line_749_valid_reg <= 2'h0 == _T_1[1:0];
    line_750_valid_reg <= 2'h1 == _T_1[1:0];
    line_751_valid_reg <= 2'h2 == _T_1[1:0];
    line_752_valid_reg <= 2'h3 == _T_1[1:0];
    line_753_valid_reg <= 2'h0 == _T_1[1:0];
    line_754_valid_reg <= 2'h1 == _T_1[1:0];
    line_755_valid_reg <= 2'h2 == _T_1[1:0];
    line_756_valid_reg <= 2'h3 == _T_1[1:0];
    line_757_valid_reg <= 2'h0 == _T_1[1:0];
    line_758_valid_reg <= 2'h1 == _T_1[1:0];
    line_759_valid_reg <= 2'h2 == _T_1[1:0];
    line_760_valid_reg <= 2'h3 == _T_1[1:0];
    line_761_valid_reg <= 2'h0 == _T_1[1:0];
    line_762_valid_reg <= 2'h1 == _T_1[1:0];
    line_763_valid_reg <= 2'h2 == _T_1[1:0];
    line_764_valid_reg <= 2'h3 == _T_1[1:0];
    line_765_valid_reg <= 2'h0 == _T_1[1:0];
    line_766_valid_reg <= 2'h1 == _T_1[1:0];
    line_767_valid_reg <= 2'h2 == _T_1[1:0];
    line_768_valid_reg <= 2'h3 == _T_1[1:0];
    line_769_valid_reg <= 2'h0 == _T_1[1:0];
    line_770_valid_reg <= 2'h1 == _T_1[1:0];
    line_771_valid_reg <= 2'h2 == _T_1[1:0];
    line_772_valid_reg <= 2'h3 == _T_1[1:0];
    line_773_valid_reg <= 2'h0 == _T_1[1:0];
    line_774_valid_reg <= 2'h1 == _T_1[1:0];
    line_775_valid_reg <= 2'h2 == _T_1[1:0];
    line_776_valid_reg <= 2'h3 == _T_1[1:0];
    line_777_valid_reg <= 2'h0 == _T_1[1:0];
    line_778_valid_reg <= 2'h1 == _T_1[1:0];
    line_779_valid_reg <= 2'h2 == _T_1[1:0];
    line_780_valid_reg <= 2'h3 == _T_1[1:0];
    line_781_valid_reg <= 2'h0 == _T_1[1:0];
    line_782_valid_reg <= 2'h1 == _T_1[1:0];
    line_783_valid_reg <= 2'h2 == _T_1[1:0];
    line_784_valid_reg <= 2'h3 == _T_1[1:0];
    line_785_valid_reg <= 2'h0 == _T_1[1:0];
    line_786_valid_reg <= 2'h1 == _T_1[1:0];
    line_787_valid_reg <= 2'h2 == _T_1[1:0];
    line_788_valid_reg <= 2'h3 == _T_1[1:0];
    line_789_valid_reg <= 2'h0 == _T_1[1:0];
    line_790_valid_reg <= 2'h1 == _T_1[1:0];
    line_791_valid_reg <= 2'h2 == _T_1[1:0];
    line_792_valid_reg <= 2'h3 == _T_1[1:0];
    line_793_valid_reg <= 2'h0 == _T_1[1:0];
    line_794_valid_reg <= 2'h1 == _T_1[1:0];
    line_795_valid_reg <= 2'h2 == _T_1[1:0];
    line_796_valid_reg <= 2'h3 == _T_1[1:0];
    line_797_valid_reg <= 2'h0 == _T_1[1:0];
    line_798_valid_reg <= 2'h1 == _T_1[1:0];
    line_799_valid_reg <= 2'h2 == _T_1[1:0];
    line_800_valid_reg <= 2'h3 == _T_1[1:0];
    line_801_valid_reg <= 2'h0 == _T_1[1:0];
    line_802_valid_reg <= 2'h1 == _T_1[1:0];
    line_803_valid_reg <= 2'h2 == _T_1[1:0];
    line_804_valid_reg <= 2'h3 == _T_1[1:0];
    line_805_valid_reg <= 2'h0 == _T_1[1:0];
    line_806_valid_reg <= 2'h1 == _T_1[1:0];
    line_807_valid_reg <= 2'h2 == _T_1[1:0];
    line_808_valid_reg <= 2'h3 == _T_1[1:0];
    line_809_valid_reg <= 2'h0 == _T_1[1:0];
    line_810_valid_reg <= 2'h1 == _T_1[1:0];
    line_811_valid_reg <= 2'h2 == _T_1[1:0];
    line_812_valid_reg <= 2'h3 == _T_1[1:0];
    line_813_valid_reg <= 2'h0 == _T_1[1:0];
    line_814_valid_reg <= 2'h1 == _T_1[1:0];
    line_815_valid_reg <= 2'h2 == _T_1[1:0];
    line_816_valid_reg <= 2'h3 == _T_1[1:0];
    line_817_valid_reg <= 2'h0 == _T_1[1:0];
    line_818_valid_reg <= 2'h1 == _T_1[1:0];
    line_819_valid_reg <= 2'h2 == _T_1[1:0];
    line_820_valid_reg <= 2'h3 == _T_1[1:0];
    line_821_valid_reg <= 2'h0 == _T_1[1:0];
    line_822_valid_reg <= 2'h1 == _T_1[1:0];
    line_823_valid_reg <= 2'h2 == _T_1[1:0];
    line_824_valid_reg <= 2'h3 == _T_1[1:0];
    line_825_valid_reg <= 2'h0 == _T_1[1:0];
    line_826_valid_reg <= 2'h1 == _T_1[1:0];
    line_827_valid_reg <= 2'h2 == _T_1[1:0];
    line_828_valid_reg <= 2'h3 == _T_1[1:0];
    line_829_valid_reg <= 2'h0 == _T_1[1:0];
    line_830_valid_reg <= 2'h1 == _T_1[1:0];
    line_831_valid_reg <= 2'h2 == _T_1[1:0];
    line_832_valid_reg <= 2'h3 == _T_1[1:0];
    line_833_valid_reg <= 2'h0 == _T_1[1:0];
    line_834_valid_reg <= 2'h1 == _T_1[1:0];
    line_835_valid_reg <= 2'h2 == _T_1[1:0];
    line_836_valid_reg <= 2'h3 == _T_1[1:0];
    line_837_valid_reg <= 2'h0 == _T_1[1:0];
    line_838_valid_reg <= 2'h1 == _T_1[1:0];
    line_839_valid_reg <= 2'h2 == _T_1[1:0];
    line_840_valid_reg <= 2'h3 == _T_1[1:0];
    line_841_valid_reg <= 2'h0 == _T_1[1:0];
    line_842_valid_reg <= 2'h1 == _T_1[1:0];
    line_843_valid_reg <= 2'h2 == _T_1[1:0];
    line_844_valid_reg <= 2'h3 == _T_1[1:0];
    line_845_valid_reg <= 2'h0 == _T_1[1:0];
    line_846_valid_reg <= 2'h1 == _T_1[1:0];
    line_847_valid_reg <= 2'h2 == _T_1[1:0];
    line_848_valid_reg <= 2'h3 == _T_1[1:0];
    line_849_valid_reg <= 2'h0 == _T_1[1:0];
    line_850_valid_reg <= 2'h1 == _T_1[1:0];
    line_851_valid_reg <= 2'h2 == _T_1[1:0];
    line_852_valid_reg <= 2'h3 == _T_1[1:0];
    line_853_valid_reg <= 2'h0 == _T_1[1:0];
    line_854_valid_reg <= 2'h1 == _T_1[1:0];
    line_855_valid_reg <= 2'h2 == _T_1[1:0];
    line_856_valid_reg <= 2'h3 == _T_1[1:0];
    line_857_valid_reg <= 2'h0 == _T_1[1:0];
    line_858_valid_reg <= 2'h1 == _T_1[1:0];
    line_859_valid_reg <= 2'h2 == _T_1[1:0];
    line_860_valid_reg <= 2'h3 == _T_1[1:0];
    line_861_valid_reg <= 2'h0 == _T_1[1:0];
    line_862_valid_reg <= 2'h1 == _T_1[1:0];
    line_863_valid_reg <= 2'h2 == _T_1[1:0];
    line_864_valid_reg <= 2'h3 == _T_1[1:0];
    line_865_valid_reg <= 2'h0 == _T_1[1:0];
    line_866_valid_reg <= 2'h1 == _T_1[1:0];
    line_867_valid_reg <= 2'h2 == _T_1[1:0];
    line_868_valid_reg <= 2'h3 == _T_1[1:0];
    line_869_valid_reg <= 2'h0 == _T_1[1:0];
    line_870_valid_reg <= 2'h1 == _T_1[1:0];
    line_871_valid_reg <= 2'h2 == _T_1[1:0];
    line_872_valid_reg <= 2'h3 == _T_1[1:0];
    line_873_valid_reg <= 2'h0 == _T_1[1:0];
    line_874_valid_reg <= 2'h1 == _T_1[1:0];
    line_875_valid_reg <= 2'h2 == _T_1[1:0];
    line_876_valid_reg <= 2'h3 == _T_1[1:0];
    line_877_valid_reg <= 2'h0 == _T_1[1:0];
    line_878_valid_reg <= 2'h1 == _T_1[1:0];
    line_879_valid_reg <= 2'h2 == _T_1[1:0];
    line_880_valid_reg <= 2'h3 == _T_1[1:0];
    line_881_valid_reg <= 2'h0 == _T_1[1:0];
    line_882_valid_reg <= 2'h1 == _T_1[1:0];
    line_883_valid_reg <= 2'h2 == _T_1[1:0];
    line_884_valid_reg <= 2'h3 == _T_1[1:0];
    line_885_valid_reg <= 2'h0 == _T_1[1:0];
    line_886_valid_reg <= 2'h1 == _T_1[1:0];
    line_887_valid_reg <= 2'h2 == _T_1[1:0];
    line_888_valid_reg <= 2'h3 == _T_1[1:0];
    line_889_valid_reg <= 2'h0 == _T_1[1:0];
    line_890_valid_reg <= 2'h1 == _T_1[1:0];
    line_891_valid_reg <= 2'h2 == _T_1[1:0];
    line_892_valid_reg <= 2'h3 == _T_1[1:0];
    line_893_valid_reg <= 2'h0 == _T_1[1:0];
    line_894_valid_reg <= 2'h1 == _T_1[1:0];
    line_895_valid_reg <= 2'h2 == _T_1[1:0];
    line_896_valid_reg <= 2'h3 == _T_1[1:0];
    line_897_valid_reg <= 2'h0 == _T_1[1:0];
    line_898_valid_reg <= 2'h1 == _T_1[1:0];
    line_899_valid_reg <= 2'h2 == _T_1[1:0];
    line_900_valid_reg <= 2'h3 == _T_1[1:0];
    line_901_valid_reg <= 2'h0 == _T_1[1:0];
    line_902_valid_reg <= 2'h1 == _T_1[1:0];
    line_903_valid_reg <= 2'h2 == _T_1[1:0];
    line_904_valid_reg <= 2'h3 == _T_1[1:0];
    line_905_valid_reg <= 2'h0 == _T_1[1:0];
    line_906_valid_reg <= 2'h1 == _T_1[1:0];
    line_907_valid_reg <= 2'h2 == _T_1[1:0];
    line_908_valid_reg <= 2'h3 == _T_1[1:0];
    line_909_valid_reg <= 2'h0 == _T_1[1:0];
    line_910_valid_reg <= 2'h1 == _T_1[1:0];
    line_911_valid_reg <= 2'h2 == _T_1[1:0];
    line_912_valid_reg <= 2'h3 == _T_1[1:0];
    line_913_valid_reg <= 2'h0 == _T_1[1:0];
    line_914_valid_reg <= 2'h1 == _T_1[1:0];
    line_915_valid_reg <= 2'h2 == _T_1[1:0];
    line_916_valid_reg <= 2'h3 == _T_1[1:0];
    line_917_valid_reg <= 2'h0 == _T_1[1:0];
    line_918_valid_reg <= 2'h1 == _T_1[1:0];
    line_919_valid_reg <= 2'h2 == _T_1[1:0];
    line_920_valid_reg <= 2'h3 == _T_1[1:0];
    line_921_valid_reg <= 2'h0 == _T_1[1:0];
    line_922_valid_reg <= 2'h1 == _T_1[1:0];
    line_923_valid_reg <= 2'h2 == _T_1[1:0];
    line_924_valid_reg <= 2'h3 == _T_1[1:0];
    line_925_valid_reg <= 2'h0 == _T_1[1:0];
    line_926_valid_reg <= 2'h1 == _T_1[1:0];
    line_927_valid_reg <= 2'h2 == _T_1[1:0];
    line_928_valid_reg <= 2'h3 == _T_1[1:0];
    line_929_valid_reg <= 2'h0 == _T_1[1:0];
    line_930_valid_reg <= 2'h1 == _T_1[1:0];
    line_931_valid_reg <= 2'h2 == _T_1[1:0];
    line_932_valid_reg <= 2'h3 == _T_1[1:0];
    line_933_valid_reg <= 2'h0 == _T_1[1:0];
    line_934_valid_reg <= 2'h1 == _T_1[1:0];
    line_935_valid_reg <= 2'h2 == _T_1[1:0];
    line_936_valid_reg <= 2'h3 == _T_1[1:0];
    line_937_valid_reg <= 2'h0 == _T_1[1:0];
    line_938_valid_reg <= 2'h1 == _T_1[1:0];
    line_939_valid_reg <= 2'h2 == _T_1[1:0];
    line_940_valid_reg <= 2'h3 == _T_1[1:0];
    line_941_valid_reg <= 2'h0 == _T_1[1:0];
    line_942_valid_reg <= 2'h1 == _T_1[1:0];
    line_943_valid_reg <= 2'h2 == _T_1[1:0];
    line_944_valid_reg <= 2'h3 == _T_1[1:0];
    line_945_valid_reg <= 2'h0 == _T_1[1:0];
    line_946_valid_reg <= 2'h1 == _T_1[1:0];
    line_947_valid_reg <= 2'h2 == _T_1[1:0];
    line_948_valid_reg <= 2'h3 == _T_1[1:0];
    line_949_valid_reg <= 2'h0 == _T_1[1:0];
    line_950_valid_reg <= 2'h1 == _T_1[1:0];
    line_951_valid_reg <= 2'h2 == _T_1[1:0];
    line_952_valid_reg <= 2'h3 == _T_1[1:0];
    line_953_valid_reg <= enqueueFire_1;
    line_954_valid_reg <= 2'h0 == _T_4;
    line_955_valid_reg <= 2'h1 == _T_4;
    line_956_valid_reg <= 2'h2 == _T_4;
    line_957_valid_reg <= 2'h3 == _T_4;
    line_958_valid_reg <= 2'h0 == _T_4;
    line_959_valid_reg <= 2'h1 == _T_4;
    line_960_valid_reg <= 2'h2 == _T_4;
    line_961_valid_reg <= 2'h3 == _T_4;
    line_962_valid_reg <= 2'h0 == _T_4;
    line_963_valid_reg <= 2'h1 == _T_4;
    line_964_valid_reg <= 2'h2 == _T_4;
    line_965_valid_reg <= 2'h3 == _T_4;
    line_966_valid_reg <= 2'h0 == _T_4;
    line_967_valid_reg <= 2'h1 == _T_4;
    line_968_valid_reg <= 2'h2 == _T_4;
    line_969_valid_reg <= 2'h3 == _T_4;
    line_970_valid_reg <= 2'h0 == _T_4;
    line_971_valid_reg <= 2'h1 == _T_4;
    line_972_valid_reg <= 2'h2 == _T_4;
    line_973_valid_reg <= 2'h3 == _T_4;
    line_974_valid_reg <= 2'h0 == _T_4;
    line_975_valid_reg <= 2'h1 == _T_4;
    line_976_valid_reg <= 2'h2 == _T_4;
    line_977_valid_reg <= 2'h3 == _T_4;
    line_978_valid_reg <= 2'h0 == _T_4;
    line_979_valid_reg <= 2'h1 == _T_4;
    line_980_valid_reg <= 2'h2 == _T_4;
    line_981_valid_reg <= 2'h3 == _T_4;
    line_982_valid_reg <= 2'h0 == _T_4;
    line_983_valid_reg <= 2'h1 == _T_4;
    line_984_valid_reg <= 2'h2 == _T_4;
    line_985_valid_reg <= 2'h3 == _T_4;
    line_986_valid_reg <= 2'h0 == _T_4;
    line_987_valid_reg <= 2'h1 == _T_4;
    line_988_valid_reg <= 2'h2 == _T_4;
    line_989_valid_reg <= 2'h3 == _T_4;
    line_990_valid_reg <= 2'h0 == _T_4;
    line_991_valid_reg <= 2'h1 == _T_4;
    line_992_valid_reg <= 2'h2 == _T_4;
    line_993_valid_reg <= 2'h3 == _T_4;
    line_994_valid_reg <= 2'h0 == _T_4;
    line_995_valid_reg <= 2'h1 == _T_4;
    line_996_valid_reg <= 2'h2 == _T_4;
    line_997_valid_reg <= 2'h3 == _T_4;
    line_998_valid_reg <= 2'h0 == _T_4;
    line_999_valid_reg <= 2'h1 == _T_4;
    line_1000_valid_reg <= 2'h2 == _T_4;
    line_1001_valid_reg <= 2'h3 == _T_4;
    line_1002_valid_reg <= 2'h0 == _T_4;
    line_1003_valid_reg <= 2'h1 == _T_4;
    line_1004_valid_reg <= 2'h2 == _T_4;
    line_1005_valid_reg <= 2'h3 == _T_4;
    line_1006_valid_reg <= 2'h0 == _T_4;
    line_1007_valid_reg <= 2'h1 == _T_4;
    line_1008_valid_reg <= 2'h2 == _T_4;
    line_1009_valid_reg <= 2'h3 == _T_4;
    line_1010_valid_reg <= 2'h0 == _T_4;
    line_1011_valid_reg <= 2'h1 == _T_4;
    line_1012_valid_reg <= 2'h2 == _T_4;
    line_1013_valid_reg <= 2'h3 == _T_4;
    line_1014_valid_reg <= 2'h0 == _T_4;
    line_1015_valid_reg <= 2'h1 == _T_4;
    line_1016_valid_reg <= 2'h2 == _T_4;
    line_1017_valid_reg <= 2'h3 == _T_4;
    line_1018_valid_reg <= 2'h0 == _T_4;
    line_1019_valid_reg <= 2'h1 == _T_4;
    line_1020_valid_reg <= 2'h2 == _T_4;
    line_1021_valid_reg <= 2'h3 == _T_4;
    line_1022_valid_reg <= 2'h0 == _T_4;
    line_1023_valid_reg <= 2'h1 == _T_4;
    line_1024_valid_reg <= 2'h2 == _T_4;
    line_1025_valid_reg <= 2'h3 == _T_4;
    line_1026_valid_reg <= 2'h0 == _T_4;
    line_1027_valid_reg <= 2'h1 == _T_4;
    line_1028_valid_reg <= 2'h2 == _T_4;
    line_1029_valid_reg <= 2'h3 == _T_4;
    line_1030_valid_reg <= 2'h0 == _T_4;
    line_1031_valid_reg <= 2'h1 == _T_4;
    line_1032_valid_reg <= 2'h2 == _T_4;
    line_1033_valid_reg <= 2'h3 == _T_4;
    line_1034_valid_reg <= 2'h0 == _T_4;
    line_1035_valid_reg <= 2'h1 == _T_4;
    line_1036_valid_reg <= 2'h2 == _T_4;
    line_1037_valid_reg <= 2'h3 == _T_4;
    line_1038_valid_reg <= 2'h0 == _T_4;
    line_1039_valid_reg <= 2'h1 == _T_4;
    line_1040_valid_reg <= 2'h2 == _T_4;
    line_1041_valid_reg <= 2'h3 == _T_4;
    line_1042_valid_reg <= 2'h0 == _T_4;
    line_1043_valid_reg <= 2'h1 == _T_4;
    line_1044_valid_reg <= 2'h2 == _T_4;
    line_1045_valid_reg <= 2'h3 == _T_4;
    line_1046_valid_reg <= 2'h0 == _T_4;
    line_1047_valid_reg <= 2'h1 == _T_4;
    line_1048_valid_reg <= 2'h2 == _T_4;
    line_1049_valid_reg <= 2'h3 == _T_4;
    line_1050_valid_reg <= 2'h0 == _T_4;
    line_1051_valid_reg <= 2'h1 == _T_4;
    line_1052_valid_reg <= 2'h2 == _T_4;
    line_1053_valid_reg <= 2'h3 == _T_4;
    line_1054_valid_reg <= 2'h0 == _T_4;
    line_1055_valid_reg <= 2'h1 == _T_4;
    line_1056_valid_reg <= 2'h2 == _T_4;
    line_1057_valid_reg <= 2'h3 == _T_4;
    line_1058_valid_reg <= 2'h0 == _T_4;
    line_1059_valid_reg <= 2'h1 == _T_4;
    line_1060_valid_reg <= 2'h2 == _T_4;
    line_1061_valid_reg <= 2'h3 == _T_4;
    line_1062_valid_reg <= 2'h0 == _T_4;
    line_1063_valid_reg <= 2'h1 == _T_4;
    line_1064_valid_reg <= 2'h2 == _T_4;
    line_1065_valid_reg <= 2'h3 == _T_4;
    line_1066_valid_reg <= 2'h0 == _T_4;
    line_1067_valid_reg <= 2'h1 == _T_4;
    line_1068_valid_reg <= 2'h2 == _T_4;
    line_1069_valid_reg <= 2'h3 == _T_4;
    line_1070_valid_reg <= 2'h0 == _T_4;
    line_1071_valid_reg <= 2'h1 == _T_4;
    line_1072_valid_reg <= 2'h2 == _T_4;
    line_1073_valid_reg <= 2'h3 == _T_4;
    line_1074_valid_reg <= 2'h0 == _T_4;
    line_1075_valid_reg <= 2'h1 == _T_4;
    line_1076_valid_reg <= 2'h2 == _T_4;
    line_1077_valid_reg <= 2'h3 == _T_4;
    line_1078_valid_reg <= 2'h0 == _T_4;
    line_1079_valid_reg <= 2'h1 == _T_4;
    line_1080_valid_reg <= 2'h2 == _T_4;
    line_1081_valid_reg <= 2'h3 == _T_4;
    line_1082_valid_reg <= 2'h0 == _T_4;
    line_1083_valid_reg <= 2'h1 == _T_4;
    line_1084_valid_reg <= 2'h2 == _T_4;
    line_1085_valid_reg <= 2'h3 == _T_4;
    line_1086_valid_reg <= 2'h0 == _T_4;
    line_1087_valid_reg <= 2'h1 == _T_4;
    line_1088_valid_reg <= 2'h2 == _T_4;
    line_1089_valid_reg <= 2'h3 == _T_4;
    line_1090_valid_reg <= 2'h0 == _T_4;
    line_1091_valid_reg <= 2'h1 == _T_4;
    line_1092_valid_reg <= 2'h2 == _T_4;
    line_1093_valid_reg <= 2'h3 == _T_4;
    line_1094_valid_reg <= 2'h0 == _T_4;
    line_1095_valid_reg <= 2'h1 == _T_4;
    line_1096_valid_reg <= 2'h2 == _T_4;
    line_1097_valid_reg <= 2'h3 == _T_4;
    line_1098_valid_reg <= 2'h0 == _T_4;
    line_1099_valid_reg <= 2'h1 == _T_4;
    line_1100_valid_reg <= 2'h2 == _T_4;
    line_1101_valid_reg <= 2'h3 == _T_4;
    line_1102_valid_reg <= 2'h0 == _T_4;
    line_1103_valid_reg <= 2'h1 == _T_4;
    line_1104_valid_reg <= 2'h2 == _T_4;
    line_1105_valid_reg <= 2'h3 == _T_4;
    line_1106_valid_reg <= 2'h0 == _T_4;
    line_1107_valid_reg <= 2'h1 == _T_4;
    line_1108_valid_reg <= 2'h2 == _T_4;
    line_1109_valid_reg <= 2'h3 == _T_4;
    line_1110_valid_reg <= 2'h0 == _T_4;
    line_1111_valid_reg <= 2'h1 == _T_4;
    line_1112_valid_reg <= 2'h2 == _T_4;
    line_1113_valid_reg <= 2'h3 == _T_4;
    line_1114_valid_reg <= 2'h0 == _T_4;
    line_1115_valid_reg <= 2'h1 == _T_4;
    line_1116_valid_reg <= 2'h2 == _T_4;
    line_1117_valid_reg <= 2'h3 == _T_4;
    line_1118_valid_reg <= 2'h0 == _T_4;
    line_1119_valid_reg <= 2'h1 == _T_4;
    line_1120_valid_reg <= 2'h2 == _T_4;
    line_1121_valid_reg <= 2'h3 == _T_4;
    line_1122_valid_reg <= 2'h0 == _T_4;
    line_1123_valid_reg <= 2'h1 == _T_4;
    line_1124_valid_reg <= 2'h2 == _T_4;
    line_1125_valid_reg <= 2'h3 == _T_4;
    line_1126_valid_reg <= 2'h0 == _T_4;
    line_1127_valid_reg <= 2'h1 == _T_4;
    line_1128_valid_reg <= 2'h2 == _T_4;
    line_1129_valid_reg <= 2'h3 == _T_4;
    line_1130_valid_reg <= 2'h0 == _T_4;
    line_1131_valid_reg <= 2'h1 == _T_4;
    line_1132_valid_reg <= 2'h2 == _T_4;
    line_1133_valid_reg <= 2'h3 == _T_4;
    line_1134_valid_reg <= 2'h0 == _T_4;
    line_1135_valid_reg <= 2'h1 == _T_4;
    line_1136_valid_reg <= 2'h2 == _T_4;
    line_1137_valid_reg <= 2'h3 == _T_4;
    line_1138_valid_reg <= 2'h0 == _T_4;
    line_1139_valid_reg <= 2'h1 == _T_4;
    line_1140_valid_reg <= 2'h2 == _T_4;
    line_1141_valid_reg <= 2'h3 == _T_4;
    line_1142_valid_reg <= 2'h0 == _T_4;
    line_1143_valid_reg <= 2'h1 == _T_4;
    line_1144_valid_reg <= 2'h2 == _T_4;
    line_1145_valid_reg <= 2'h3 == _T_4;
    line_1146_valid_reg <= 2'h0 == _T_4;
    line_1147_valid_reg <= 2'h1 == _T_4;
    line_1148_valid_reg <= 2'h2 == _T_4;
    line_1149_valid_reg <= 2'h3 == _T_4;
    line_1150_valid_reg <= 2'h0 == _T_4;
    line_1151_valid_reg <= 2'h1 == _T_4;
    line_1152_valid_reg <= 2'h2 == _T_4;
    line_1153_valid_reg <= 2'h3 == _T_4;
    line_1154_valid_reg <= 2'h0 == _T_4;
    line_1155_valid_reg <= 2'h1 == _T_4;
    line_1156_valid_reg <= 2'h2 == _T_4;
    line_1157_valid_reg <= 2'h3 == _T_4;
    line_1158_valid_reg <= 2'h0 == _T_4;
    line_1159_valid_reg <= 2'h1 == _T_4;
    line_1160_valid_reg <= 2'h2 == _T_4;
    line_1161_valid_reg <= 2'h3 == _T_4;
    line_1162_valid_reg <= 2'h0 == _T_4;
    line_1163_valid_reg <= 2'h1 == _T_4;
    line_1164_valid_reg <= 2'h2 == _T_4;
    line_1165_valid_reg <= 2'h3 == _T_4;
    line_1166_valid_reg <= 2'h0 == _T_4;
    line_1167_valid_reg <= 2'h1 == _T_4;
    line_1168_valid_reg <= 2'h2 == _T_4;
    line_1169_valid_reg <= 2'h3 == _T_4;
    line_1170_valid_reg <= 2'h0 == _T_4;
    line_1171_valid_reg <= 2'h1 == _T_4;
    line_1172_valid_reg <= 2'h2 == _T_4;
    line_1173_valid_reg <= 2'h3 == _T_4;
    line_1174_valid_reg <= 2'h0 == _T_4;
    line_1175_valid_reg <= 2'h1 == _T_4;
    line_1176_valid_reg <= 2'h2 == _T_4;
    line_1177_valid_reg <= 2'h3 == _T_4;
    line_1178_valid_reg <= 2'h0 == ringBufferTail;
    line_1179_valid_reg <= 2'h1 == ringBufferTail;
    line_1180_valid_reg <= 2'h2 == ringBufferTail;
    line_1181_valid_reg <= 2'h3 == ringBufferTail;
    line_1182_valid_reg <= 2'h0 == ringBufferTail;
    line_1183_valid_reg <= 2'h1 == ringBufferTail;
    line_1184_valid_reg <= 2'h2 == ringBufferTail;
    line_1185_valid_reg <= 2'h3 == ringBufferTail;
    line_1186_valid_reg <= 2'h0 == ringBufferTail;
    line_1187_valid_reg <= 2'h1 == ringBufferTail;
    line_1188_valid_reg <= 2'h2 == ringBufferTail;
    line_1189_valid_reg <= 2'h3 == ringBufferTail;
    line_1190_valid_reg <= 2'h0 == ringBufferTail;
    line_1191_valid_reg <= 2'h1 == ringBufferTail;
    line_1192_valid_reg <= 2'h2 == ringBufferTail;
    line_1193_valid_reg <= 2'h3 == ringBufferTail;
    line_1194_valid_reg <= 2'h0 == ringBufferTail;
    line_1195_valid_reg <= 2'h1 == ringBufferTail;
    line_1196_valid_reg <= 2'h2 == ringBufferTail;
    line_1197_valid_reg <= 2'h3 == ringBufferTail;
    line_1198_valid_reg <= 2'h0 == ringBufferTail;
    line_1199_valid_reg <= 2'h1 == ringBufferTail;
    line_1200_valid_reg <= 2'h2 == ringBufferTail;
    line_1201_valid_reg <= 2'h3 == ringBufferTail;
    line_1202_valid_reg <= 2'h0 == ringBufferTail;
    line_1203_valid_reg <= 2'h1 == ringBufferTail;
    line_1204_valid_reg <= 2'h2 == ringBufferTail;
    line_1205_valid_reg <= 2'h3 == ringBufferTail;
    line_1206_valid_reg <= 2'h0 == ringBufferTail;
    line_1207_valid_reg <= 2'h1 == ringBufferTail;
    line_1208_valid_reg <= 2'h2 == ringBufferTail;
    line_1209_valid_reg <= 2'h3 == ringBufferTail;
    line_1210_valid_reg <= 2'h0 == ringBufferTail;
    line_1211_valid_reg <= 2'h1 == ringBufferTail;
    line_1212_valid_reg <= 2'h2 == ringBufferTail;
    line_1213_valid_reg <= 2'h3 == ringBufferTail;
    line_1214_valid_reg <= 2'h0 == ringBufferTail;
    line_1215_valid_reg <= 2'h1 == ringBufferTail;
    line_1216_valid_reg <= 2'h2 == ringBufferTail;
    line_1217_valid_reg <= 2'h3 == ringBufferTail;
    line_1218_valid_reg <= 2'h0 == ringBufferTail;
    line_1219_valid_reg <= 2'h1 == ringBufferTail;
    line_1220_valid_reg <= 2'h2 == ringBufferTail;
    line_1221_valid_reg <= 2'h3 == ringBufferTail;
    line_1222_valid_reg <= 2'h0 == ringBufferTail;
    line_1223_valid_reg <= 2'h1 == ringBufferTail;
    line_1224_valid_reg <= 2'h2 == ringBufferTail;
    line_1225_valid_reg <= 2'h3 == ringBufferTail;
    line_1226_valid_reg <= 2'h0 == ringBufferTail;
    line_1227_valid_reg <= 2'h1 == ringBufferTail;
    line_1228_valid_reg <= 2'h2 == ringBufferTail;
    line_1229_valid_reg <= 2'h3 == ringBufferTail;
    line_1230_valid_reg <= 2'h0 == ringBufferTail;
    line_1231_valid_reg <= 2'h1 == ringBufferTail;
    line_1232_valid_reg <= 2'h2 == ringBufferTail;
    line_1233_valid_reg <= 2'h3 == ringBufferTail;
    line_1234_valid_reg <= 2'h0 == ringBufferTail;
    line_1235_valid_reg <= 2'h1 == ringBufferTail;
    line_1236_valid_reg <= 2'h2 == ringBufferTail;
    line_1237_valid_reg <= 2'h3 == ringBufferTail;
    line_1238_valid_reg <= 2'h0 == ringBufferTail;
    line_1239_valid_reg <= 2'h1 == ringBufferTail;
    line_1240_valid_reg <= 2'h2 == ringBufferTail;
    line_1241_valid_reg <= 2'h3 == ringBufferTail;
    line_1242_valid_reg <= 2'h0 == ringBufferTail;
    line_1243_valid_reg <= 2'h1 == ringBufferTail;
    line_1244_valid_reg <= 2'h2 == ringBufferTail;
    line_1245_valid_reg <= 2'h3 == ringBufferTail;
    line_1246_valid_reg <= 2'h0 == ringBufferTail;
    line_1247_valid_reg <= 2'h1 == ringBufferTail;
    line_1248_valid_reg <= 2'h2 == ringBufferTail;
    line_1249_valid_reg <= 2'h3 == ringBufferTail;
    line_1250_valid_reg <= 2'h0 == ringBufferTail;
    line_1251_valid_reg <= 2'h1 == ringBufferTail;
    line_1252_valid_reg <= 2'h2 == ringBufferTail;
    line_1253_valid_reg <= 2'h3 == ringBufferTail;
    line_1254_valid_reg <= 2'h0 == ringBufferTail;
    line_1255_valid_reg <= 2'h1 == ringBufferTail;
    line_1256_valid_reg <= 2'h2 == ringBufferTail;
    line_1257_valid_reg <= 2'h3 == ringBufferTail;
    line_1258_valid_reg <= 2'h0 == ringBufferTail;
    line_1259_valid_reg <= 2'h1 == ringBufferTail;
    line_1260_valid_reg <= 2'h2 == ringBufferTail;
    line_1261_valid_reg <= 2'h3 == ringBufferTail;
    line_1262_valid_reg <= 2'h0 == ringBufferTail;
    line_1263_valid_reg <= 2'h1 == ringBufferTail;
    line_1264_valid_reg <= 2'h2 == ringBufferTail;
    line_1265_valid_reg <= 2'h3 == ringBufferTail;
    line_1266_valid_reg <= 2'h0 == ringBufferTail;
    line_1267_valid_reg <= 2'h1 == ringBufferTail;
    line_1268_valid_reg <= 2'h2 == ringBufferTail;
    line_1269_valid_reg <= 2'h3 == ringBufferTail;
    line_1270_valid_reg <= 2'h0 == ringBufferTail;
    line_1271_valid_reg <= 2'h1 == ringBufferTail;
    line_1272_valid_reg <= 2'h2 == ringBufferTail;
    line_1273_valid_reg <= 2'h3 == ringBufferTail;
    line_1274_valid_reg <= 2'h0 == ringBufferTail;
    line_1275_valid_reg <= 2'h1 == ringBufferTail;
    line_1276_valid_reg <= 2'h2 == ringBufferTail;
    line_1277_valid_reg <= 2'h3 == ringBufferTail;
    line_1278_valid_reg <= 2'h0 == ringBufferTail;
    line_1279_valid_reg <= 2'h1 == ringBufferTail;
    line_1280_valid_reg <= 2'h2 == ringBufferTail;
    line_1281_valid_reg <= 2'h3 == ringBufferTail;
    line_1282_valid_reg <= 2'h0 == ringBufferTail;
    line_1283_valid_reg <= 2'h1 == ringBufferTail;
    line_1284_valid_reg <= 2'h2 == ringBufferTail;
    line_1285_valid_reg <= 2'h3 == ringBufferTail;
    line_1286_valid_reg <= 2'h0 == ringBufferTail;
    line_1287_valid_reg <= 2'h1 == ringBufferTail;
    line_1288_valid_reg <= 2'h2 == ringBufferTail;
    line_1289_valid_reg <= 2'h3 == ringBufferTail;
    line_1290_valid_reg <= 2'h0 == ringBufferTail;
    line_1291_valid_reg <= 2'h1 == ringBufferTail;
    line_1292_valid_reg <= 2'h2 == ringBufferTail;
    line_1293_valid_reg <= 2'h3 == ringBufferTail;
    line_1294_valid_reg <= 2'h0 == ringBufferTail;
    line_1295_valid_reg <= 2'h1 == ringBufferTail;
    line_1296_valid_reg <= 2'h2 == ringBufferTail;
    line_1297_valid_reg <= 2'h3 == ringBufferTail;
    line_1298_valid_reg <= 2'h0 == ringBufferTail;
    line_1299_valid_reg <= 2'h1 == ringBufferTail;
    line_1300_valid_reg <= 2'h2 == ringBufferTail;
    line_1301_valid_reg <= 2'h3 == ringBufferTail;
    line_1302_valid_reg <= 2'h0 == ringBufferTail;
    line_1303_valid_reg <= 2'h1 == ringBufferTail;
    line_1304_valid_reg <= 2'h2 == ringBufferTail;
    line_1305_valid_reg <= 2'h3 == ringBufferTail;
    line_1306_valid_reg <= 2'h0 == ringBufferTail;
    line_1307_valid_reg <= 2'h1 == ringBufferTail;
    line_1308_valid_reg <= 2'h2 == ringBufferTail;
    line_1309_valid_reg <= 2'h3 == ringBufferTail;
    line_1310_valid_reg <= 2'h0 == ringBufferTail;
    line_1311_valid_reg <= 2'h1 == ringBufferTail;
    line_1312_valid_reg <= 2'h2 == ringBufferTail;
    line_1313_valid_reg <= 2'h3 == ringBufferTail;
    line_1314_valid_reg <= 2'h0 == ringBufferTail;
    line_1315_valid_reg <= 2'h1 == ringBufferTail;
    line_1316_valid_reg <= 2'h2 == ringBufferTail;
    line_1317_valid_reg <= 2'h3 == ringBufferTail;
    line_1318_valid_reg <= 2'h0 == ringBufferTail;
    line_1319_valid_reg <= 2'h1 == ringBufferTail;
    line_1320_valid_reg <= 2'h2 == ringBufferTail;
    line_1321_valid_reg <= 2'h3 == ringBufferTail;
    line_1322_valid_reg <= 2'h0 == ringBufferTail;
    line_1323_valid_reg <= 2'h1 == ringBufferTail;
    line_1324_valid_reg <= 2'h2 == ringBufferTail;
    line_1325_valid_reg <= 2'h3 == ringBufferTail;
    line_1326_valid_reg <= 2'h0 == ringBufferTail;
    line_1327_valid_reg <= 2'h1 == ringBufferTail;
    line_1328_valid_reg <= 2'h2 == ringBufferTail;
    line_1329_valid_reg <= 2'h3 == ringBufferTail;
    line_1330_valid_reg <= 2'h0 == ringBufferTail;
    line_1331_valid_reg <= 2'h1 == ringBufferTail;
    line_1332_valid_reg <= 2'h2 == ringBufferTail;
    line_1333_valid_reg <= 2'h3 == ringBufferTail;
    line_1334_valid_reg <= 2'h0 == ringBufferTail;
    line_1335_valid_reg <= 2'h1 == ringBufferTail;
    line_1336_valid_reg <= 2'h2 == ringBufferTail;
    line_1337_valid_reg <= 2'h3 == ringBufferTail;
    line_1338_valid_reg <= 2'h0 == ringBufferTail;
    line_1339_valid_reg <= 2'h1 == ringBufferTail;
    line_1340_valid_reg <= 2'h2 == ringBufferTail;
    line_1341_valid_reg <= 2'h3 == ringBufferTail;
    line_1342_valid_reg <= 2'h0 == ringBufferTail;
    line_1343_valid_reg <= 2'h1 == ringBufferTail;
    line_1344_valid_reg <= 2'h2 == ringBufferTail;
    line_1345_valid_reg <= 2'h3 == ringBufferTail;
    line_1346_valid_reg <= 2'h0 == ringBufferTail;
    line_1347_valid_reg <= 2'h1 == ringBufferTail;
    line_1348_valid_reg <= 2'h2 == ringBufferTail;
    line_1349_valid_reg <= 2'h3 == ringBufferTail;
    line_1350_valid_reg <= 2'h0 == ringBufferTail;
    line_1351_valid_reg <= 2'h1 == ringBufferTail;
    line_1352_valid_reg <= 2'h2 == ringBufferTail;
    line_1353_valid_reg <= 2'h3 == ringBufferTail;
    line_1354_valid_reg <= 2'h0 == ringBufferTail;
    line_1355_valid_reg <= 2'h1 == ringBufferTail;
    line_1356_valid_reg <= 2'h2 == ringBufferTail;
    line_1357_valid_reg <= 2'h3 == ringBufferTail;
    line_1358_valid_reg <= 2'h0 == ringBufferTail;
    line_1359_valid_reg <= 2'h1 == ringBufferTail;
    line_1360_valid_reg <= 2'h2 == ringBufferTail;
    line_1361_valid_reg <= 2'h3 == ringBufferTail;
    line_1362_valid_reg <= 2'h0 == ringBufferTail;
    line_1363_valid_reg <= 2'h1 == ringBufferTail;
    line_1364_valid_reg <= 2'h2 == ringBufferTail;
    line_1365_valid_reg <= 2'h3 == ringBufferTail;
    line_1366_valid_reg <= 2'h0 == ringBufferTail;
    line_1367_valid_reg <= 2'h1 == ringBufferTail;
    line_1368_valid_reg <= 2'h2 == ringBufferTail;
    line_1369_valid_reg <= 2'h3 == ringBufferTail;
    line_1370_valid_reg <= 2'h0 == ringBufferTail;
    line_1371_valid_reg <= 2'h1 == ringBufferTail;
    line_1372_valid_reg <= 2'h2 == ringBufferTail;
    line_1373_valid_reg <= 2'h3 == ringBufferTail;
    line_1374_valid_reg <= 2'h0 == ringBufferTail;
    line_1375_valid_reg <= 2'h1 == ringBufferTail;
    line_1376_valid_reg <= 2'h2 == ringBufferTail;
    line_1377_valid_reg <= 2'h3 == ringBufferTail;
    line_1378_valid_reg <= 2'h0 == ringBufferTail;
    line_1379_valid_reg <= 2'h1 == ringBufferTail;
    line_1380_valid_reg <= 2'h2 == ringBufferTail;
    line_1381_valid_reg <= 2'h3 == ringBufferTail;
    line_1382_valid_reg <= 2'h0 == ringBufferTail;
    line_1383_valid_reg <= 2'h1 == ringBufferTail;
    line_1384_valid_reg <= 2'h2 == ringBufferTail;
    line_1385_valid_reg <= 2'h3 == ringBufferTail;
    line_1386_valid_reg <= 2'h0 == ringBufferTail;
    line_1387_valid_reg <= 2'h1 == ringBufferTail;
    line_1388_valid_reg <= 2'h2 == ringBufferTail;
    line_1389_valid_reg <= 2'h3 == ringBufferTail;
    line_1390_valid_reg <= 2'h0 == ringBufferTail;
    line_1391_valid_reg <= 2'h1 == ringBufferTail;
    line_1392_valid_reg <= 2'h2 == ringBufferTail;
    line_1393_valid_reg <= 2'h3 == ringBufferTail;
    line_1394_valid_reg <= 2'h0 == ringBufferTail;
    line_1395_valid_reg <= 2'h1 == ringBufferTail;
    line_1396_valid_reg <= 2'h2 == ringBufferTail;
    line_1397_valid_reg <= 2'h3 == ringBufferTail;
    line_1398_valid_reg <= 2'h0 == ringBufferTail;
    line_1399_valid_reg <= 2'h1 == ringBufferTail;
    line_1400_valid_reg <= 2'h2 == ringBufferTail;
    line_1401_valid_reg <= 2'h3 == ringBufferTail;
    line_1402_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1403_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1404_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1405_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1406_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1407_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1408_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1409_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1410_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1411_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1412_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1413_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1414_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1415_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1416_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1417_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1418_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1419_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1420_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1421_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1422_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1423_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1424_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1425_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1426_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1427_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1428_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1429_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1430_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1431_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1432_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1433_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1434_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1435_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1436_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1437_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1438_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1439_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1440_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1441_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1442_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1443_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1444_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1445_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1446_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1447_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1448_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1449_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1450_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1451_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1452_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1453_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1454_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1455_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1456_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1457_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1458_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1459_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1460_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1461_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1462_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1463_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1464_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1465_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1466_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1467_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1468_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1469_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1470_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1471_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1472_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1473_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1474_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1475_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1476_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1477_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1478_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1479_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1480_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1481_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1482_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1483_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1484_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1485_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1486_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1487_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1488_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1489_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1490_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1491_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1492_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1493_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1494_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1495_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1496_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1497_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1498_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1499_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1500_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1501_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1502_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1503_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1504_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1505_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1506_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1507_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1508_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1509_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1510_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1511_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1512_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1513_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1514_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1515_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1516_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1517_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1518_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1519_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1520_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1521_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1522_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1523_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1524_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1525_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1526_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1527_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1528_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1529_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1530_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1531_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1532_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1533_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1534_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1535_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1536_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1537_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1538_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1539_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1540_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1541_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1542_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1543_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1544_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1545_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1546_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1547_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1548_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1549_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1550_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1551_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1552_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1553_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1554_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1555_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1556_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1557_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1558_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1559_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1560_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1561_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1562_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1563_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1564_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1565_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1566_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1567_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1568_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1569_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1570_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1571_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1572_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1573_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1574_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1575_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1576_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1577_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1578_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1579_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1580_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1581_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1582_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1583_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1584_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1585_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1586_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1587_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1588_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1589_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1590_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1591_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1592_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1593_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1594_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1595_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1596_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1597_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1598_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1599_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1600_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1601_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1602_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1603_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1604_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1605_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1606_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1607_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1608_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1609_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1610_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1611_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1612_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1613_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1614_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1615_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1616_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1617_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1618_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1619_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1620_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1621_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1622_valid_reg <= 2'h0 == deq2_StartIndex;
    line_1623_valid_reg <= 2'h1 == deq2_StartIndex;
    line_1624_valid_reg <= 2'h2 == deq2_StartIndex;
    line_1625_valid_reg <= 2'h3 == deq2_StartIndex;
    line_1626_valid_reg <= dequeueFire;
    line_1627_valid_reg <= frontend_io_flushVec[1];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataBuffer_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dataBuffer_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  dataBuffer_0_cf_crossBoundaryFault = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  dataBuffer_0_ctrl_isNutCoreTrap = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  dataBuffer_0_data_imm = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  dataBuffer_1_cf_instr = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  dataBuffer_1_cf_pc = _RAND_25[38:0];
  _RAND_26 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_12 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  dataBuffer_1_cf_crossBoundaryFault = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  dataBuffer_1_ctrl_isNutCoreTrap = _RAND_46[0:0];
  _RAND_47 = {2{`RANDOM}};
  dataBuffer_1_data_imm = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  dataBuffer_2_cf_instr = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  dataBuffer_2_cf_pc = _RAND_49[38:0];
  _RAND_50 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc = _RAND_50[38:0];
  _RAND_51 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  dataBuffer_2_cf_crossBoundaryFault = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  dataBuffer_2_ctrl_isNutCoreTrap = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  dataBuffer_2_data_imm = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  dataBuffer_3_cf_instr = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  dataBuffer_3_cf_pc = _RAND_73[38:0];
  _RAND_74 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc = _RAND_74[38:0];
  _RAND_75 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  dataBuffer_3_cf_crossBoundaryFault = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1 = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  dataBuffer_3_ctrl_isNutCoreTrap = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  dataBuffer_3_data_imm = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  ringBufferHead = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  ringBufferTail = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  line_727_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_728_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_729_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_730_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_731_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_732_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_733_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_734_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_735_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_736_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_737_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_738_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_739_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_740_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_741_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_742_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_743_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_744_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_745_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_746_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_747_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_748_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_749_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_750_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_751_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_752_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_753_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_754_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_755_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_756_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_757_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_758_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_759_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_760_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_761_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_762_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_763_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_764_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_765_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_766_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_767_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_768_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_769_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_770_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_771_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_772_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_773_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_774_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_775_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_776_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_777_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_778_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_779_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_780_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_781_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_782_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_783_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_784_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_785_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_786_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_787_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_788_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_789_valid_reg = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  line_790_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  line_791_valid_reg = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  line_792_valid_reg = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  line_793_valid_reg = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  line_794_valid_reg = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  line_795_valid_reg = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  line_796_valid_reg = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  line_797_valid_reg = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  line_798_valid_reg = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  line_799_valid_reg = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  line_800_valid_reg = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  line_801_valid_reg = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  line_802_valid_reg = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  line_803_valid_reg = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  line_804_valid_reg = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  line_805_valid_reg = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  line_806_valid_reg = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  line_807_valid_reg = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  line_808_valid_reg = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  line_809_valid_reg = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  line_810_valid_reg = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  line_811_valid_reg = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  line_812_valid_reg = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  line_813_valid_reg = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  line_814_valid_reg = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  line_815_valid_reg = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  line_816_valid_reg = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  line_817_valid_reg = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  line_818_valid_reg = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  line_819_valid_reg = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  line_820_valid_reg = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  line_821_valid_reg = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  line_822_valid_reg = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  line_823_valid_reg = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  line_824_valid_reg = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  line_825_valid_reg = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  line_826_valid_reg = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  line_827_valid_reg = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  line_828_valid_reg = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  line_829_valid_reg = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  line_830_valid_reg = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  line_831_valid_reg = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  line_832_valid_reg = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  line_833_valid_reg = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  line_834_valid_reg = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  line_835_valid_reg = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  line_836_valid_reg = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  line_837_valid_reg = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  line_838_valid_reg = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  line_839_valid_reg = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  line_840_valid_reg = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  line_841_valid_reg = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  line_842_valid_reg = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  line_843_valid_reg = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  line_844_valid_reg = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  line_845_valid_reg = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  line_846_valid_reg = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  line_847_valid_reg = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  line_848_valid_reg = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  line_849_valid_reg = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  line_850_valid_reg = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  line_851_valid_reg = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  line_852_valid_reg = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  line_853_valid_reg = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  line_854_valid_reg = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  line_855_valid_reg = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  line_856_valid_reg = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  line_857_valid_reg = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  line_858_valid_reg = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  line_859_valid_reg = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  line_860_valid_reg = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  line_861_valid_reg = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  line_862_valid_reg = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  line_863_valid_reg = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  line_864_valid_reg = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  line_865_valid_reg = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  line_866_valid_reg = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  line_867_valid_reg = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  line_868_valid_reg = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  line_869_valid_reg = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  line_870_valid_reg = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  line_871_valid_reg = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  line_872_valid_reg = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  line_873_valid_reg = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  line_874_valid_reg = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  line_875_valid_reg = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  line_876_valid_reg = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  line_877_valid_reg = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  line_878_valid_reg = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  line_879_valid_reg = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  line_880_valid_reg = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  line_881_valid_reg = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  line_882_valid_reg = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  line_883_valid_reg = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  line_884_valid_reg = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  line_885_valid_reg = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  line_886_valid_reg = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  line_887_valid_reg = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  line_888_valid_reg = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  line_889_valid_reg = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  line_890_valid_reg = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  line_891_valid_reg = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  line_892_valid_reg = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  line_893_valid_reg = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  line_894_valid_reg = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  line_895_valid_reg = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  line_896_valid_reg = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  line_897_valid_reg = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  line_898_valid_reg = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  line_899_valid_reg = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  line_900_valid_reg = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  line_901_valid_reg = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  line_902_valid_reg = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  line_903_valid_reg = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  line_904_valid_reg = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  line_905_valid_reg = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  line_906_valid_reg = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  line_907_valid_reg = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  line_908_valid_reg = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  line_909_valid_reg = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  line_910_valid_reg = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  line_911_valid_reg = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  line_912_valid_reg = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  line_913_valid_reg = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  line_914_valid_reg = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  line_915_valid_reg = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  line_916_valid_reg = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  line_917_valid_reg = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  line_918_valid_reg = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  line_919_valid_reg = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  line_920_valid_reg = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  line_921_valid_reg = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  line_922_valid_reg = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  line_923_valid_reg = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  line_924_valid_reg = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  line_925_valid_reg = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  line_926_valid_reg = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  line_927_valid_reg = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  line_928_valid_reg = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  line_929_valid_reg = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  line_930_valid_reg = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  line_931_valid_reg = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  line_932_valid_reg = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  line_933_valid_reg = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  line_934_valid_reg = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  line_935_valid_reg = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  line_936_valid_reg = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  line_937_valid_reg = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  line_938_valid_reg = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  line_939_valid_reg = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  line_940_valid_reg = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  line_941_valid_reg = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  line_942_valid_reg = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  line_943_valid_reg = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  line_944_valid_reg = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  line_945_valid_reg = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  line_946_valid_reg = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  line_947_valid_reg = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  line_948_valid_reg = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  line_949_valid_reg = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  line_950_valid_reg = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  line_951_valid_reg = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  line_952_valid_reg = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  line_953_valid_reg = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  line_954_valid_reg = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  line_955_valid_reg = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  line_956_valid_reg = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  line_957_valid_reg = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  line_958_valid_reg = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  line_959_valid_reg = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  line_960_valid_reg = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  line_961_valid_reg = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  line_962_valid_reg = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  line_963_valid_reg = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  line_964_valid_reg = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  line_965_valid_reg = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  line_966_valid_reg = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  line_967_valid_reg = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  line_968_valid_reg = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  line_969_valid_reg = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  line_970_valid_reg = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  line_971_valid_reg = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  line_972_valid_reg = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  line_973_valid_reg = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  line_974_valid_reg = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  line_975_valid_reg = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  line_976_valid_reg = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  line_977_valid_reg = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  line_978_valid_reg = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  line_979_valid_reg = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  line_980_valid_reg = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  line_981_valid_reg = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  line_982_valid_reg = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  line_983_valid_reg = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  line_984_valid_reg = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  line_985_valid_reg = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  line_986_valid_reg = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  line_987_valid_reg = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  line_988_valid_reg = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  line_989_valid_reg = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  line_990_valid_reg = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  line_991_valid_reg = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  line_992_valid_reg = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  line_993_valid_reg = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  line_994_valid_reg = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  line_995_valid_reg = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  line_996_valid_reg = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  line_997_valid_reg = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  line_998_valid_reg = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  line_999_valid_reg = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  line_1000_valid_reg = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  line_1001_valid_reg = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  line_1002_valid_reg = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  line_1003_valid_reg = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  line_1004_valid_reg = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  line_1005_valid_reg = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  line_1006_valid_reg = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  line_1007_valid_reg = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  line_1008_valid_reg = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  line_1009_valid_reg = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  line_1010_valid_reg = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  line_1011_valid_reg = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  line_1012_valid_reg = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  line_1013_valid_reg = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  line_1014_valid_reg = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  line_1015_valid_reg = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  line_1016_valid_reg = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  line_1017_valid_reg = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  line_1018_valid_reg = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  line_1019_valid_reg = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  line_1020_valid_reg = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  line_1021_valid_reg = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  line_1022_valid_reg = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  line_1023_valid_reg = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  line_1024_valid_reg = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  line_1025_valid_reg = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  line_1026_valid_reg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  line_1027_valid_reg = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  line_1028_valid_reg = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  line_1029_valid_reg = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  line_1030_valid_reg = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  line_1031_valid_reg = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  line_1032_valid_reg = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  line_1033_valid_reg = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  line_1034_valid_reg = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  line_1035_valid_reg = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  line_1036_valid_reg = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  line_1037_valid_reg = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  line_1038_valid_reg = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  line_1039_valid_reg = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  line_1040_valid_reg = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  line_1041_valid_reg = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  line_1042_valid_reg = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  line_1043_valid_reg = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  line_1044_valid_reg = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  line_1045_valid_reg = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  line_1046_valid_reg = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  line_1047_valid_reg = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  line_1048_valid_reg = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  line_1049_valid_reg = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  line_1050_valid_reg = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  line_1051_valid_reg = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  line_1052_valid_reg = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  line_1053_valid_reg = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  line_1054_valid_reg = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  line_1055_valid_reg = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  line_1056_valid_reg = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  line_1057_valid_reg = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  line_1058_valid_reg = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  line_1059_valid_reg = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  line_1060_valid_reg = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  line_1061_valid_reg = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  line_1062_valid_reg = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  line_1063_valid_reg = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  line_1064_valid_reg = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  line_1065_valid_reg = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  line_1066_valid_reg = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  line_1067_valid_reg = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  line_1068_valid_reg = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  line_1069_valid_reg = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  line_1070_valid_reg = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  line_1071_valid_reg = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  line_1072_valid_reg = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  line_1073_valid_reg = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  line_1074_valid_reg = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  line_1075_valid_reg = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  line_1076_valid_reg = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  line_1077_valid_reg = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  line_1078_valid_reg = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  line_1079_valid_reg = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  line_1080_valid_reg = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  line_1081_valid_reg = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  line_1082_valid_reg = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  line_1083_valid_reg = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  line_1084_valid_reg = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  line_1085_valid_reg = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  line_1086_valid_reg = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  line_1087_valid_reg = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  line_1088_valid_reg = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  line_1089_valid_reg = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  line_1090_valid_reg = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  line_1091_valid_reg = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  line_1092_valid_reg = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  line_1093_valid_reg = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  line_1094_valid_reg = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  line_1095_valid_reg = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  line_1096_valid_reg = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  line_1097_valid_reg = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  line_1098_valid_reg = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  line_1099_valid_reg = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  line_1100_valid_reg = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  line_1101_valid_reg = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  line_1102_valid_reg = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  line_1103_valid_reg = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  line_1104_valid_reg = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  line_1105_valid_reg = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  line_1106_valid_reg = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  line_1107_valid_reg = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  line_1108_valid_reg = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  line_1109_valid_reg = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  line_1110_valid_reg = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  line_1111_valid_reg = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  line_1112_valid_reg = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  line_1113_valid_reg = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  line_1114_valid_reg = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  line_1115_valid_reg = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  line_1116_valid_reg = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  line_1117_valid_reg = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  line_1118_valid_reg = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  line_1119_valid_reg = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  line_1120_valid_reg = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  line_1121_valid_reg = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  line_1122_valid_reg = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  line_1123_valid_reg = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  line_1124_valid_reg = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  line_1125_valid_reg = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  line_1126_valid_reg = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  line_1127_valid_reg = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  line_1128_valid_reg = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  line_1129_valid_reg = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  line_1130_valid_reg = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  line_1131_valid_reg = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  line_1132_valid_reg = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  line_1133_valid_reg = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  line_1134_valid_reg = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  line_1135_valid_reg = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  line_1136_valid_reg = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  line_1137_valid_reg = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  line_1138_valid_reg = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  line_1139_valid_reg = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  line_1140_valid_reg = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  line_1141_valid_reg = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  line_1142_valid_reg = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  line_1143_valid_reg = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  line_1144_valid_reg = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  line_1145_valid_reg = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  line_1146_valid_reg = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  line_1147_valid_reg = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  line_1148_valid_reg = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  line_1149_valid_reg = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  line_1150_valid_reg = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  line_1151_valid_reg = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  line_1152_valid_reg = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  line_1153_valid_reg = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  line_1154_valid_reg = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  line_1155_valid_reg = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  line_1156_valid_reg = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  line_1157_valid_reg = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  line_1158_valid_reg = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  line_1159_valid_reg = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  line_1160_valid_reg = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  line_1161_valid_reg = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  line_1162_valid_reg = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  line_1163_valid_reg = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  line_1164_valid_reg = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  line_1165_valid_reg = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  line_1166_valid_reg = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  line_1167_valid_reg = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  line_1168_valid_reg = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  line_1169_valid_reg = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  line_1170_valid_reg = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  line_1171_valid_reg = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  line_1172_valid_reg = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  line_1173_valid_reg = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  line_1174_valid_reg = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  line_1175_valid_reg = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  line_1176_valid_reg = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  line_1177_valid_reg = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  line_1178_valid_reg = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  line_1179_valid_reg = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  line_1180_valid_reg = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  line_1181_valid_reg = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  line_1182_valid_reg = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  line_1183_valid_reg = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  line_1184_valid_reg = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  line_1185_valid_reg = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  line_1186_valid_reg = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  line_1187_valid_reg = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  line_1188_valid_reg = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  line_1189_valid_reg = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  line_1190_valid_reg = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  line_1191_valid_reg = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  line_1192_valid_reg = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  line_1193_valid_reg = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  line_1194_valid_reg = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  line_1195_valid_reg = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  line_1196_valid_reg = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  line_1197_valid_reg = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  line_1198_valid_reg = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  line_1199_valid_reg = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  line_1200_valid_reg = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  line_1201_valid_reg = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  line_1202_valid_reg = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  line_1203_valid_reg = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  line_1204_valid_reg = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  line_1205_valid_reg = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  line_1206_valid_reg = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  line_1207_valid_reg = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  line_1208_valid_reg = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  line_1209_valid_reg = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  line_1210_valid_reg = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  line_1211_valid_reg = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  line_1212_valid_reg = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  line_1213_valid_reg = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  line_1214_valid_reg = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  line_1215_valid_reg = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  line_1216_valid_reg = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  line_1217_valid_reg = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  line_1218_valid_reg = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  line_1219_valid_reg = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  line_1220_valid_reg = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  line_1221_valid_reg = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  line_1222_valid_reg = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  line_1223_valid_reg = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  line_1224_valid_reg = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  line_1225_valid_reg = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  line_1226_valid_reg = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  line_1227_valid_reg = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  line_1228_valid_reg = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  line_1229_valid_reg = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  line_1230_valid_reg = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  line_1231_valid_reg = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  line_1232_valid_reg = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  line_1233_valid_reg = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  line_1234_valid_reg = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  line_1235_valid_reg = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  line_1236_valid_reg = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  line_1237_valid_reg = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  line_1238_valid_reg = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  line_1239_valid_reg = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  line_1240_valid_reg = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  line_1241_valid_reg = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  line_1242_valid_reg = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  line_1243_valid_reg = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  line_1244_valid_reg = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  line_1245_valid_reg = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  line_1246_valid_reg = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  line_1247_valid_reg = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  line_1248_valid_reg = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  line_1249_valid_reg = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  line_1250_valid_reg = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  line_1251_valid_reg = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  line_1252_valid_reg = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  line_1253_valid_reg = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  line_1254_valid_reg = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  line_1255_valid_reg = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  line_1256_valid_reg = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  line_1257_valid_reg = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  line_1258_valid_reg = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  line_1259_valid_reg = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  line_1260_valid_reg = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  line_1261_valid_reg = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  line_1262_valid_reg = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  line_1263_valid_reg = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  line_1264_valid_reg = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  line_1265_valid_reg = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  line_1266_valid_reg = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  line_1267_valid_reg = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  line_1268_valid_reg = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  line_1269_valid_reg = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  line_1270_valid_reg = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  line_1271_valid_reg = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  line_1272_valid_reg = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  line_1273_valid_reg = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  line_1274_valid_reg = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  line_1275_valid_reg = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  line_1276_valid_reg = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  line_1277_valid_reg = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  line_1278_valid_reg = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  line_1279_valid_reg = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  line_1280_valid_reg = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  line_1281_valid_reg = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  line_1282_valid_reg = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  line_1283_valid_reg = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  line_1284_valid_reg = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  line_1285_valid_reg = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  line_1286_valid_reg = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  line_1287_valid_reg = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  line_1288_valid_reg = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  line_1289_valid_reg = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  line_1290_valid_reg = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  line_1291_valid_reg = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  line_1292_valid_reg = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  line_1293_valid_reg = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  line_1294_valid_reg = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  line_1295_valid_reg = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  line_1296_valid_reg = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  line_1297_valid_reg = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  line_1298_valid_reg = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  line_1299_valid_reg = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  line_1300_valid_reg = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  line_1301_valid_reg = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  line_1302_valid_reg = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  line_1303_valid_reg = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  line_1304_valid_reg = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  line_1305_valid_reg = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  line_1306_valid_reg = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  line_1307_valid_reg = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  line_1308_valid_reg = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  line_1309_valid_reg = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  line_1310_valid_reg = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  line_1311_valid_reg = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  line_1312_valid_reg = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  line_1313_valid_reg = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  line_1314_valid_reg = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  line_1315_valid_reg = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  line_1316_valid_reg = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  line_1317_valid_reg = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  line_1318_valid_reg = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  line_1319_valid_reg = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  line_1320_valid_reg = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  line_1321_valid_reg = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  line_1322_valid_reg = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  line_1323_valid_reg = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  line_1324_valid_reg = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  line_1325_valid_reg = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  line_1326_valid_reg = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  line_1327_valid_reg = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  line_1328_valid_reg = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  line_1329_valid_reg = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  line_1330_valid_reg = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  line_1331_valid_reg = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  line_1332_valid_reg = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  line_1333_valid_reg = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  line_1334_valid_reg = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  line_1335_valid_reg = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  line_1336_valid_reg = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  line_1337_valid_reg = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  line_1338_valid_reg = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  line_1339_valid_reg = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  line_1340_valid_reg = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  line_1341_valid_reg = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  line_1342_valid_reg = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  line_1343_valid_reg = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  line_1344_valid_reg = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  line_1345_valid_reg = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  line_1346_valid_reg = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  line_1347_valid_reg = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  line_1348_valid_reg = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  line_1349_valid_reg = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  line_1350_valid_reg = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  line_1351_valid_reg = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  line_1352_valid_reg = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  line_1353_valid_reg = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  line_1354_valid_reg = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  line_1355_valid_reg = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  line_1356_valid_reg = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  line_1357_valid_reg = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  line_1358_valid_reg = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  line_1359_valid_reg = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  line_1360_valid_reg = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  line_1361_valid_reg = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  line_1362_valid_reg = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  line_1363_valid_reg = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  line_1364_valid_reg = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  line_1365_valid_reg = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  line_1366_valid_reg = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  line_1367_valid_reg = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  line_1368_valid_reg = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  line_1369_valid_reg = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  line_1370_valid_reg = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  line_1371_valid_reg = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  line_1372_valid_reg = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  line_1373_valid_reg = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  line_1374_valid_reg = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  line_1375_valid_reg = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  line_1376_valid_reg = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  line_1377_valid_reg = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  line_1378_valid_reg = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  line_1379_valid_reg = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  line_1380_valid_reg = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  line_1381_valid_reg = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  line_1382_valid_reg = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  line_1383_valid_reg = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  line_1384_valid_reg = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  line_1385_valid_reg = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  line_1386_valid_reg = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  line_1387_valid_reg = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  line_1388_valid_reg = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  line_1389_valid_reg = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  line_1390_valid_reg = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  line_1391_valid_reg = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  line_1392_valid_reg = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  line_1393_valid_reg = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  line_1394_valid_reg = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  line_1395_valid_reg = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  line_1396_valid_reg = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  line_1397_valid_reg = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  line_1398_valid_reg = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  line_1399_valid_reg = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  line_1400_valid_reg = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  line_1401_valid_reg = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  line_1402_valid_reg = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  line_1403_valid_reg = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  line_1404_valid_reg = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  line_1405_valid_reg = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  line_1406_valid_reg = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  line_1407_valid_reg = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  line_1408_valid_reg = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  line_1409_valid_reg = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  line_1410_valid_reg = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  line_1411_valid_reg = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  line_1412_valid_reg = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  line_1413_valid_reg = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  line_1414_valid_reg = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  line_1415_valid_reg = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  line_1416_valid_reg = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  line_1417_valid_reg = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  line_1418_valid_reg = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  line_1419_valid_reg = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  line_1420_valid_reg = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  line_1421_valid_reg = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  line_1422_valid_reg = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  line_1423_valid_reg = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  line_1424_valid_reg = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  line_1425_valid_reg = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  line_1426_valid_reg = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  line_1427_valid_reg = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  line_1428_valid_reg = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  line_1429_valid_reg = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  line_1430_valid_reg = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  line_1431_valid_reg = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  line_1432_valid_reg = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  line_1433_valid_reg = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  line_1434_valid_reg = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  line_1435_valid_reg = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  line_1436_valid_reg = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  line_1437_valid_reg = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  line_1438_valid_reg = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  line_1439_valid_reg = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  line_1440_valid_reg = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  line_1441_valid_reg = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  line_1442_valid_reg = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  line_1443_valid_reg = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  line_1444_valid_reg = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  line_1445_valid_reg = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  line_1446_valid_reg = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  line_1447_valid_reg = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  line_1448_valid_reg = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  line_1449_valid_reg = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  line_1450_valid_reg = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  line_1451_valid_reg = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  line_1452_valid_reg = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  line_1453_valid_reg = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  line_1454_valid_reg = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  line_1455_valid_reg = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  line_1456_valid_reg = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  line_1457_valid_reg = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  line_1458_valid_reg = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  line_1459_valid_reg = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  line_1460_valid_reg = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  line_1461_valid_reg = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  line_1462_valid_reg = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  line_1463_valid_reg = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  line_1464_valid_reg = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  line_1465_valid_reg = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  line_1466_valid_reg = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  line_1467_valid_reg = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  line_1468_valid_reg = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  line_1469_valid_reg = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  line_1470_valid_reg = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  line_1471_valid_reg = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  line_1472_valid_reg = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  line_1473_valid_reg = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  line_1474_valid_reg = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  line_1475_valid_reg = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  line_1476_valid_reg = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  line_1477_valid_reg = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  line_1478_valid_reg = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  line_1479_valid_reg = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  line_1480_valid_reg = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  line_1481_valid_reg = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  line_1482_valid_reg = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  line_1483_valid_reg = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  line_1484_valid_reg = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  line_1485_valid_reg = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  line_1486_valid_reg = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  line_1487_valid_reg = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  line_1488_valid_reg = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  line_1489_valid_reg = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  line_1490_valid_reg = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  line_1491_valid_reg = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  line_1492_valid_reg = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  line_1493_valid_reg = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  line_1494_valid_reg = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  line_1495_valid_reg = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  line_1496_valid_reg = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  line_1497_valid_reg = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  line_1498_valid_reg = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  line_1499_valid_reg = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  line_1500_valid_reg = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  line_1501_valid_reg = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  line_1502_valid_reg = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  line_1503_valid_reg = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  line_1504_valid_reg = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  line_1505_valid_reg = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  line_1506_valid_reg = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  line_1507_valid_reg = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  line_1508_valid_reg = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  line_1509_valid_reg = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  line_1510_valid_reg = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  line_1511_valid_reg = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  line_1512_valid_reg = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  line_1513_valid_reg = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  line_1514_valid_reg = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  line_1515_valid_reg = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  line_1516_valid_reg = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  line_1517_valid_reg = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  line_1518_valid_reg = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  line_1519_valid_reg = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  line_1520_valid_reg = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  line_1521_valid_reg = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  line_1522_valid_reg = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  line_1523_valid_reg = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  line_1524_valid_reg = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  line_1525_valid_reg = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  line_1526_valid_reg = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  line_1527_valid_reg = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  line_1528_valid_reg = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  line_1529_valid_reg = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  line_1530_valid_reg = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  line_1531_valid_reg = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  line_1532_valid_reg = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  line_1533_valid_reg = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  line_1534_valid_reg = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  line_1535_valid_reg = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  line_1536_valid_reg = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  line_1537_valid_reg = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  line_1538_valid_reg = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  line_1539_valid_reg = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  line_1540_valid_reg = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  line_1541_valid_reg = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  line_1542_valid_reg = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  line_1543_valid_reg = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  line_1544_valid_reg = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  line_1545_valid_reg = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  line_1546_valid_reg = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  line_1547_valid_reg = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  line_1548_valid_reg = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  line_1549_valid_reg = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  line_1550_valid_reg = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  line_1551_valid_reg = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  line_1552_valid_reg = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  line_1553_valid_reg = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  line_1554_valid_reg = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  line_1555_valid_reg = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  line_1556_valid_reg = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  line_1557_valid_reg = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  line_1558_valid_reg = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  line_1559_valid_reg = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  line_1560_valid_reg = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  line_1561_valid_reg = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  line_1562_valid_reg = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  line_1563_valid_reg = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  line_1564_valid_reg = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  line_1565_valid_reg = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  line_1566_valid_reg = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  line_1567_valid_reg = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  line_1568_valid_reg = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  line_1569_valid_reg = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  line_1570_valid_reg = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  line_1571_valid_reg = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  line_1572_valid_reg = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  line_1573_valid_reg = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  line_1574_valid_reg = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  line_1575_valid_reg = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  line_1576_valid_reg = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  line_1577_valid_reg = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  line_1578_valid_reg = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  line_1579_valid_reg = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  line_1580_valid_reg = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  line_1581_valid_reg = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  line_1582_valid_reg = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  line_1583_valid_reg = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  line_1584_valid_reg = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  line_1585_valid_reg = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  line_1586_valid_reg = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  line_1587_valid_reg = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  line_1588_valid_reg = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  line_1589_valid_reg = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  line_1590_valid_reg = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  line_1591_valid_reg = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  line_1592_valid_reg = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  line_1593_valid_reg = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  line_1594_valid_reg = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  line_1595_valid_reg = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  line_1596_valid_reg = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  line_1597_valid_reg = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  line_1598_valid_reg = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  line_1599_valid_reg = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  line_1600_valid_reg = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  line_1601_valid_reg = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  line_1602_valid_reg = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  line_1603_valid_reg = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  line_1604_valid_reg = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  line_1605_valid_reg = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  line_1606_valid_reg = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  line_1607_valid_reg = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  line_1608_valid_reg = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  line_1609_valid_reg = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  line_1610_valid_reg = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  line_1611_valid_reg = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  line_1612_valid_reg = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  line_1613_valid_reg = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  line_1614_valid_reg = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  line_1615_valid_reg = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  line_1616_valid_reg = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  line_1617_valid_reg = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  line_1618_valid_reg = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  line_1619_valid_reg = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  line_1620_valid_reg = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  line_1621_valid_reg = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  line_1622_valid_reg = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  line_1623_valid_reg = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  line_1624_valid_reg = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  line_1625_valid_reg = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  line_1626_valid_reg = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  line_1627_valid_reg = _RAND_998[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_0) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_2) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_0 & _GEN_3) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_225) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_226) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_227) begin
      cover(1'h1);
    end
    //
    if (wen & enqueueFire_1 & _GEN_228) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h1 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h2 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h3 == ringBufferTail) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h0 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h1 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h2 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (2'h3 == deq2_StartIndex) begin
      cover(1'h1);
    end
    //
    if (dequeueFire) begin
      cover(1'h1);
    end
    //
    if (frontend_io_flushVec[1]) begin
      cover(1'h1);
    end
  end
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_in_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_in_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_out_mem_resp_bits_rdata // @[src/main/scala/system/Coherence.scala 31:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/system/Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[src/main/scala/system/Coherence.scala 46:24]
  wire  _T_12 = ~reset; // @[src/main/scala/system/Coherence.scala 49:9]
  wire  line_1628_clock;
  wire  line_1628_reset;
  wire  line_1628_valid;
  reg  line_1628_valid_reg;
  wire  _reqLatch_T = ~inflight; // @[src/main/scala/system/Coherence.scala 52:42]
  reg [31:0] reqLatch_addr; // @[src/main/scala/system/Coherence.scala 52:27]
  wire  line_1629_clock;
  wire  line_1629_reset;
  wire  line_1629_valid;
  reg  line_1629_valid_reg;
  wire  _io_out_mem_req_valid_T_1 = io_in_req_valid & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 65:43]
  wire  _T_19 = 3'h0 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1630_clock;
  wire  line_1630_reset;
  wire  line_1630_valid;
  reg  line_1630_valid_reg;
  wire  _T_20 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1631_clock;
  wire  line_1631_reset;
  wire  line_1631_valid;
  reg  line_1631_valid_reg;
  wire  line_1632_clock;
  wire  line_1632_reset;
  wire  line_1632_valid;
  reg  line_1632_valid_reg;
  wire  _T_27 = 3'h1 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1633_clock;
  wire  line_1633_reset;
  wire  line_1633_valid;
  reg  line_1633_valid_reg;
  wire  line_1634_clock;
  wire  line_1634_reset;
  wire  line_1634_valid;
  reg  line_1634_valid_reg;
  wire  _T_29 = 3'h2 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1635_clock;
  wire  line_1635_reset;
  wire  line_1635_valid;
  reg  line_1635_valid_reg;
  wire  _T_31 = io_in_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire  _T_32 = io_in_resp_valid & _T_31; // @[src/main/scala/system/Coherence.scala 89:29]
  wire  line_1636_clock;
  wire  line_1636_reset;
  wire  line_1636_valid;
  reg  line_1636_valid_reg;
  wire [2:0] _GEN_40 = io_in_resp_valid & _T_31 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 89:{60,68}]
  wire  line_1637_clock;
  wire  line_1637_reset;
  wire  line_1637_valid;
  reg  line_1637_valid_reg;
  wire  _T_33 = 3'h3 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1638_clock;
  wire  line_1638_reset;
  wire  line_1638_valid;
  reg  line_1638_valid_reg;
  wire  _T_34 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1639_clock;
  wire  line_1639_reset;
  wire  line_1639_valid;
  reg  line_1639_valid_reg;
  wire [2:0] _GEN_41 = _T_34 ? 3'h4 : state; // @[src/main/scala/system/Coherence.scala 45:22 94:{36,44}]
  wire  line_1640_clock;
  wire  line_1640_reset;
  wire  line_1640_valid;
  reg  line_1640_valid_reg;
  wire  _T_35 = 3'h4 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1641_clock;
  wire  line_1641_reset;
  wire  line_1641_valid;
  reg  line_1641_valid_reg;
  wire  _T_36 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_37 = io_out_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire  _T_38 = _T_36 & _T_37; // @[src/main/scala/system/Coherence.scala 96:55]
  wire  line_1642_clock;
  wire  line_1642_reset;
  wire  line_1642_valid;
  reg  line_1642_valid_reg;
  wire [2:0] _GEN_42 = _T_36 & _T_37 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 96:101 45:22 96:93]
  wire  line_1643_clock;
  wire  line_1643_reset;
  wire  line_1643_valid;
  reg  line_1643_valid_reg;
  wire  _T_39 = 3'h5 == state; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  line_1644_clock;
  wire  line_1644_reset;
  wire  line_1644_valid;
  reg  line_1644_valid_reg;
  wire  line_1645_clock;
  wire  line_1645_reset;
  wire  line_1645_valid;
  reg  line_1645_valid_reg;
  wire [2:0] _GEN_43 = _T_36 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 97:{57,65}]
  wire [2:0] _GEN_44 = 3'h5 == state ? _GEN_43 : state; // @[src/main/scala/system/Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_45 = 3'h4 == state ? _GEN_42 : _GEN_44; // @[src/main/scala/system/Coherence.scala 74:18]
  wire [31:0] _GEN_46 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_51 = 3'h3 == state | _io_out_mem_req_valid_T_1; // @[src/main/scala/system/Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_52 = 3'h3 == state ? _GEN_41 : _GEN_45; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_54 = 3'h2 == state ? 1'h0 : io_out_mem_resp_valid; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_55 = 3'h2 == state ? 4'h0 : io_out_mem_resp_bits_cmd; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_56 = 3'h2 == state ? 64'h0 : io_out_mem_resp_bits_rdata; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [31:0] _GEN_58 = 3'h2 == state ? io_in_req_bits_addr : _GEN_46; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_63 = 3'h2 == state ? _io_out_mem_req_valid_T_1 : _GEN_51; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_66 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_54; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_67 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_55; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_68 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_56; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [31:0] _GEN_69 = 3'h1 == state ? io_in_req_bits_addr : _GEN_58; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_74 = 3'h1 == state ? _io_out_mem_req_valid_T_1 : _GEN_63; // @[src/main/scala/system/Coherence.scala 74:18]
  GEN_w1_line #(.COVER_INDEX(1628)) line_1628 (
    .clock(line_1628_clock),
    .reset(line_1628_reset),
    .valid(line_1628_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1629)) line_1629 (
    .clock(line_1629_clock),
    .reset(line_1629_reset),
    .valid(line_1629_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1630)) line_1630 (
    .clock(line_1630_clock),
    .reset(line_1630_reset),
    .valid(line_1630_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1631)) line_1631 (
    .clock(line_1631_clock),
    .reset(line_1631_reset),
    .valid(line_1631_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1632)) line_1632 (
    .clock(line_1632_clock),
    .reset(line_1632_reset),
    .valid(line_1632_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1633)) line_1633 (
    .clock(line_1633_clock),
    .reset(line_1633_reset),
    .valid(line_1633_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1634)) line_1634 (
    .clock(line_1634_clock),
    .reset(line_1634_reset),
    .valid(line_1634_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1635)) line_1635 (
    .clock(line_1635_clock),
    .reset(line_1635_reset),
    .valid(line_1635_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1636)) line_1636 (
    .clock(line_1636_clock),
    .reset(line_1636_reset),
    .valid(line_1636_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1637)) line_1637 (
    .clock(line_1637_clock),
    .reset(line_1637_reset),
    .valid(line_1637_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1638)) line_1638 (
    .clock(line_1638_clock),
    .reset(line_1638_reset),
    .valid(line_1638_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1639)) line_1639 (
    .clock(line_1639_clock),
    .reset(line_1639_reset),
    .valid(line_1639_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1640)) line_1640 (
    .clock(line_1640_clock),
    .reset(line_1640_reset),
    .valid(line_1640_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1641)) line_1641 (
    .clock(line_1641_clock),
    .reset(line_1641_reset),
    .valid(line_1641_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1642)) line_1642 (
    .clock(line_1642_clock),
    .reset(line_1642_reset),
    .valid(line_1642_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1643)) line_1643 (
    .clock(line_1643_clock),
    .reset(line_1643_reset),
    .valid(line_1643_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1644)) line_1644 (
    .clock(line_1644_clock),
    .reset(line_1644_reset),
    .valid(line_1644_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1645)) line_1645 (
    .clock(line_1645_clock),
    .reset(line_1645_reset),
    .valid(line_1645_valid)
  );
  assign line_1628_clock = clock;
  assign line_1628_reset = reset;
  assign line_1628_valid = _T_12 ^ line_1628_valid_reg;
  assign line_1629_clock = clock;
  assign line_1629_reset = reset;
  assign line_1629_valid = _reqLatch_T ^ line_1629_valid_reg;
  assign line_1630_clock = clock;
  assign line_1630_reset = reset;
  assign line_1630_valid = _T_19 ^ line_1630_valid_reg;
  assign line_1631_clock = clock;
  assign line_1631_reset = reset;
  assign line_1631_valid = _T_20 ^ line_1631_valid_reg;
  assign line_1632_clock = clock;
  assign line_1632_reset = reset;
  assign line_1632_valid = _T_19 ^ line_1632_valid_reg;
  assign line_1633_clock = clock;
  assign line_1633_reset = reset;
  assign line_1633_valid = _T_27 ^ line_1633_valid_reg;
  assign line_1634_clock = clock;
  assign line_1634_reset = reset;
  assign line_1634_valid = _T_27 ^ line_1634_valid_reg;
  assign line_1635_clock = clock;
  assign line_1635_reset = reset;
  assign line_1635_valid = _T_29 ^ line_1635_valid_reg;
  assign line_1636_clock = clock;
  assign line_1636_reset = reset;
  assign line_1636_valid = _T_32 ^ line_1636_valid_reg;
  assign line_1637_clock = clock;
  assign line_1637_reset = reset;
  assign line_1637_valid = _T_29 ^ line_1637_valid_reg;
  assign line_1638_clock = clock;
  assign line_1638_reset = reset;
  assign line_1638_valid = _T_33 ^ line_1638_valid_reg;
  assign line_1639_clock = clock;
  assign line_1639_reset = reset;
  assign line_1639_valid = _T_34 ^ line_1639_valid_reg;
  assign line_1640_clock = clock;
  assign line_1640_reset = reset;
  assign line_1640_valid = _T_33 ^ line_1640_valid_reg;
  assign line_1641_clock = clock;
  assign line_1641_reset = reset;
  assign line_1641_valid = _T_35 ^ line_1641_valid_reg;
  assign line_1642_clock = clock;
  assign line_1642_reset = reset;
  assign line_1642_valid = _T_38 ^ line_1642_valid_reg;
  assign line_1643_clock = clock;
  assign line_1643_reset = reset;
  assign line_1643_valid = _T_35 ^ line_1643_valid_reg;
  assign line_1644_clock = clock;
  assign line_1644_reset = reset;
  assign line_1644_valid = _T_39 ^ line_1644_valid_reg;
  assign line_1645_clock = clock;
  assign line_1645_reset = reset;
  assign line_1645_valid = _T_36 ^ line_1645_valid_reg;
  assign io_in_req_ready = io_out_mem_req_ready & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 66:43]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_66; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_67; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_68; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _io_out_mem_req_valid_T_1 : _GEN_74; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_69; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/system/Coherence.scala 72:14]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/system/Coherence.scala 45:22]
      state <= 3'h0; // @[src/main/scala/system/Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (_T_20) begin // @[src/main/scala/system/Coherence.scala 76:29]
        state <= 3'h4;
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (3'h2 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
        state <= _GEN_40;
      end else begin
        state <= _GEN_52;
      end
    end
    line_1628_valid_reg <= _T_12;
    if (~inflight) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_addr <= io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 52:27]
    end
    line_1629_valid_reg <= _reqLatch_T;
    line_1630_valid_reg <= _T_19;
    line_1631_valid_reg <= _T_20;
    line_1632_valid_reg <= _T_19;
    line_1633_valid_reg <= _T_27;
    line_1634_valid_reg <= _T_27;
    line_1635_valid_reg <= _T_29;
    line_1636_valid_reg <= _T_32;
    line_1637_valid_reg <= _T_29;
    line_1638_valid_reg <= _T_33;
    line_1639_valid_reg <= _T_34;
    line_1640_valid_reg <= _T_33;
    line_1641_valid_reg <= _T_35;
    line_1642_valid_reg <= _T_38;
    line_1643_valid_reg <= _T_35;
    line_1644_valid_reg <= _T_39;
    line_1645_valid_reg <= _T_36;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  line_1628_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  line_1629_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1630_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1631_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1632_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1633_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1634_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1635_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1636_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1637_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1638_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1639_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1640_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1641_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1642_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1643_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1644_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1645_valid_reg = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_12) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/system/Coherence.scala 49:9]
    end
    //
    if (_reqLatch_T) begin
      cover(1'h1);
    end
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_19) begin
      cover(1'h1);
    end
    //
    if (_T_19 & _T_20) begin
      cover(1'h1);
    end
    //
    if (_T_19 & _T_20) begin
      cover(1'h1);
    end
    //
    if (~_T_19) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & _T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & _T_29) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & _T_29 & _T_32) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & _T_33) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & _T_33 & _T_34) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33 & _T_35) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33 & _T_35 & _T_38) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33 & ~_T_35) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33 & ~_T_35 & _T_39) begin
      cover(1'h1);
    end
    //
    if (~_T_19 & ~_T_27 & ~_T_29 & ~_T_33 & ~_T_35 & _T_39 & _T_36) begin
      cover(1'h1);
    end
  end
endmodule
module LockingArbiter_2(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  line_1646_clock;
  wire  line_1646_reset;
  wire  line_1646_valid;
  reg  line_1646_valid_reg;
  wire  line_1647_clock;
  wire  line_1647_reset;
  wire  line_1647_valid;
  reg  line_1647_valid_reg;
  wire  line_1648_clock;
  wire  line_1648_reset;
  wire  line_1648_valid;
  reg  line_1648_valid_reg;
  wire  line_1649_clock;
  wire  line_1649_reset;
  wire  line_1649_valid;
  reg  line_1649_valid_reg;
  wire  line_1650_clock;
  wire  line_1650_reset;
  wire  line_1650_valid;
  reg  line_1650_valid_reg;
  wire  line_1651_clock;
  wire  line_1651_reset;
  wire  line_1651_valid;
  reg  line_1651_valid_reg;
  wire  line_1652_clock;
  wire  line_1652_reset;
  wire  line_1652_valid;
  reg  line_1652_valid_reg;
  wire  line_1653_clock;
  wire  line_1653_reset;
  wire  line_1653_valid;
  reg  line_1653_valid_reg;
  wire  line_1654_clock;
  wire  line_1654_reset;
  wire  line_1654_valid;
  reg  line_1654_valid_reg;
  wire  line_1655_clock;
  wire  line_1655_reset;
  wire  line_1655_valid;
  reg  line_1655_valid_reg;
  wire  line_1656_clock;
  wire  line_1656_reset;
  wire  line_1656_valid;
  reg  line_1656_valid_reg;
  wire  line_1657_clock;
  wire  line_1657_reset;
  wire  line_1657_valid;
  reg  line_1657_valid_reg;
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & wantsLock; // @[src/main/scala/chisel3/util/Arbiter.scala 64:22]
  wire  line_1658_clock;
  wire  line_1658_reset;
  wire  line_1658_valid;
  reg  line_1658_valid_reg;
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1659_clock;
  wire  line_1659_reset;
  wire  line_1659_valid;
  reg  line_1659_valid_reg;
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  line_1660_clock;
  wire  line_1660_reset;
  wire  line_1660_valid;
  reg  line_1660_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1646)) line_1646 (
    .clock(line_1646_clock),
    .reset(line_1646_reset),
    .valid(line_1646_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1647)) line_1647 (
    .clock(line_1647_clock),
    .reset(line_1647_reset),
    .valid(line_1647_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1648)) line_1648 (
    .clock(line_1648_clock),
    .reset(line_1648_reset),
    .valid(line_1648_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1649)) line_1649 (
    .clock(line_1649_clock),
    .reset(line_1649_reset),
    .valid(line_1649_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1650)) line_1650 (
    .clock(line_1650_clock),
    .reset(line_1650_reset),
    .valid(line_1650_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1651)) line_1651 (
    .clock(line_1651_clock),
    .reset(line_1651_reset),
    .valid(line_1651_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1652)) line_1652 (
    .clock(line_1652_clock),
    .reset(line_1652_reset),
    .valid(line_1652_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1653)) line_1653 (
    .clock(line_1653_clock),
    .reset(line_1653_reset),
    .valid(line_1653_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1654)) line_1654 (
    .clock(line_1654_clock),
    .reset(line_1654_reset),
    .valid(line_1654_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1655)) line_1655 (
    .clock(line_1655_clock),
    .reset(line_1655_reset),
    .valid(line_1655_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1656)) line_1656 (
    .clock(line_1656_clock),
    .reset(line_1656_reset),
    .valid(line_1656_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1657)) line_1657 (
    .clock(line_1657_clock),
    .reset(line_1657_reset),
    .valid(line_1657_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1658)) line_1658 (
    .clock(line_1658_clock),
    .reset(line_1658_reset),
    .valid(line_1658_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1659)) line_1659 (
    .clock(line_1659_clock),
    .reset(line_1659_reset),
    .valid(line_1659_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1660)) line_1660 (
    .clock(line_1660_clock),
    .reset(line_1660_reset),
    .valid(line_1660_valid)
  );
  assign line_1646_clock = clock;
  assign line_1646_reset = reset;
  assign line_1646_valid = ~io_chosen ^ line_1646_valid_reg;
  assign line_1647_clock = clock;
  assign line_1647_reset = reset;
  assign line_1647_valid = io_chosen ^ line_1647_valid_reg;
  assign line_1648_clock = clock;
  assign line_1648_reset = reset;
  assign line_1648_valid = ~io_chosen ^ line_1648_valid_reg;
  assign line_1649_clock = clock;
  assign line_1649_reset = reset;
  assign line_1649_valid = io_chosen ^ line_1649_valid_reg;
  assign line_1650_clock = clock;
  assign line_1650_reset = reset;
  assign line_1650_valid = ~io_chosen ^ line_1650_valid_reg;
  assign line_1651_clock = clock;
  assign line_1651_reset = reset;
  assign line_1651_valid = io_chosen ^ line_1651_valid_reg;
  assign line_1652_clock = clock;
  assign line_1652_reset = reset;
  assign line_1652_valid = ~io_chosen ^ line_1652_valid_reg;
  assign line_1653_clock = clock;
  assign line_1653_reset = reset;
  assign line_1653_valid = io_chosen ^ line_1653_valid_reg;
  assign line_1654_clock = clock;
  assign line_1654_reset = reset;
  assign line_1654_valid = ~io_chosen ^ line_1654_valid_reg;
  assign line_1655_clock = clock;
  assign line_1655_reset = reset;
  assign line_1655_valid = io_chosen ^ line_1655_valid_reg;
  assign line_1656_clock = clock;
  assign line_1656_reset = reset;
  assign line_1656_valid = ~io_chosen ^ line_1656_valid_reg;
  assign line_1657_clock = clock;
  assign line_1657_reset = reset;
  assign line_1657_valid = io_chosen ^ line_1657_valid_reg;
  assign line_1658_clock = clock;
  assign line_1658_reset = reset;
  assign line_1658_valid = _T_1 ^ line_1658_valid_reg;
  assign line_1659_clock = clock;
  assign line_1659_reset = reset;
  assign line_1659_valid = locked ^ line_1659_valid_reg;
  assign line_1660_clock = clock;
  assign line_1660_reset = reset;
  assign line_1660_valid = io_in_0_valid ^ line_1660_valid_reg;
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    line_1646_valid_reg <= ~io_chosen;
    line_1647_valid_reg <= io_chosen;
    line_1648_valid_reg <= ~io_chosen;
    line_1649_valid_reg <= io_chosen;
    line_1650_valid_reg <= ~io_chosen;
    line_1651_valid_reg <= io_chosen;
    line_1652_valid_reg <= ~io_chosen;
    line_1653_valid_reg <= io_chosen;
    line_1654_valid_reg <= ~io_chosen;
    line_1655_valid_reg <= io_chosen;
    line_1656_valid_reg <= ~io_chosen;
    line_1657_valid_reg <= io_chosen;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    line_1658_valid_reg <= _T_1;
    line_1659_valid_reg <= locked;
    line_1660_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1646_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1647_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1648_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1649_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1650_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1651_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1652_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1653_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1654_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1655_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1656_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1657_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lockCount_value = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  lockIdx = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1658_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1659_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1660_valid_reg = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (~io_chosen) begin
      cover(1'h1);
    end
    //
    if (io_chosen) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (locked) begin
      cover(1'h1);
    end
    //
    if (io_in_0_valid) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusCrossbarNto1_2(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_0_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_1_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:29]
  wire  _T_12 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_1661_clock;
  wire  line_1661_reset;
  wire  line_1661_valid;
  reg  line_1661_valid_reg;
  wire  _T_13 = ~(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
  wire  line_1662_clock;
  wire  line_1662_reset;
  wire  line_1662_valid;
  reg  line_1662_valid_reg;
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  line_1663_clock;
  wire  line_1663_reset;
  wire  line_1663_valid;
  reg  line_1663_valid_reg;
  wire  line_1664_clock;
  wire  line_1664_reset;
  wire  line_1664_valid;
  reg  line_1664_valid_reg;
  wire  line_1665_clock;
  wire  line_1665_reset;
  wire  line_1665_valid;
  reg  line_1665_valid_reg;
  wire  line_1666_clock;
  wire  line_1666_reset;
  wire  line_1666_valid;
  reg  line_1666_valid_reg;
  wire  _T_14 = 2'h0 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_1667_clock;
  wire  line_1667_reset;
  wire  line_1667_valid;
  reg  line_1667_valid_reg;
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1668_clock;
  wire  line_1668_reset;
  wire  line_1668_valid;
  reg  line_1668_valid_reg;
  wire  line_1669_clock;
  wire  line_1669_reset;
  wire  line_1669_valid;
  reg  line_1669_valid_reg;
  wire  line_1670_clock;
  wire  line_1670_reset;
  wire  line_1670_valid;
  reg  line_1670_valid_reg;
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire  _T_23 = _T_21 | _T_22; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:47]
  wire  line_1671_clock;
  wire  line_1671_reset;
  wire  line_1671_valid;
  reg  line_1671_valid_reg;
  wire [1:0] _GEN_21 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  line_1672_clock;
  wire  line_1672_reset;
  wire  line_1672_valid;
  reg  line_1672_valid_reg;
  wire  _T_24 = 2'h1 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_1673_clock;
  wire  line_1673_reset;
  wire  line_1673_valid;
  reg  line_1673_valid_reg;
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire  _T_27 = _T_25 & _T_26; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:48]
  wire  line_1674_clock;
  wire  line_1674_reset;
  wire  line_1674_valid;
  reg  line_1674_valid_reg;
  wire  line_1675_clock;
  wire  line_1675_reset;
  wire  line_1675_valid;
  reg  line_1675_valid_reg;
  wire  _T_28 = 2'h2 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
  wire  line_1676_clock;
  wire  line_1676_reset;
  wire  line_1676_valid;
  reg  line_1676_valid_reg;
  wire  line_1677_clock;
  wire  line_1677_reset;
  wire  line_1677_valid;
  reg  line_1677_valid_reg;
  wire [1:0] _GEN_26 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter_2 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w1_line #(.COVER_INDEX(1661)) line_1661 (
    .clock(line_1661_clock),
    .reset(line_1661_reset),
    .valid(line_1661_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1662)) line_1662 (
    .clock(line_1662_clock),
    .reset(line_1662_reset),
    .valid(line_1662_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1663)) line_1663 (
    .clock(line_1663_clock),
    .reset(line_1663_reset),
    .valid(line_1663_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1664)) line_1664 (
    .clock(line_1664_clock),
    .reset(line_1664_reset),
    .valid(line_1664_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1665)) line_1665 (
    .clock(line_1665_clock),
    .reset(line_1665_reset),
    .valid(line_1665_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1666)) line_1666 (
    .clock(line_1666_clock),
    .reset(line_1666_reset),
    .valid(line_1666_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1667)) line_1667 (
    .clock(line_1667_clock),
    .reset(line_1667_reset),
    .valid(line_1667_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1668)) line_1668 (
    .clock(line_1668_clock),
    .reset(line_1668_reset),
    .valid(line_1668_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1669)) line_1669 (
    .clock(line_1669_clock),
    .reset(line_1669_reset),
    .valid(line_1669_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1670)) line_1670 (
    .clock(line_1670_clock),
    .reset(line_1670_reset),
    .valid(line_1670_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1671)) line_1671 (
    .clock(line_1671_clock),
    .reset(line_1671_reset),
    .valid(line_1671_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1672)) line_1672 (
    .clock(line_1672_clock),
    .reset(line_1672_reset),
    .valid(line_1672_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1673)) line_1673 (
    .clock(line_1673_clock),
    .reset(line_1673_reset),
    .valid(line_1673_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1674)) line_1674 (
    .clock(line_1674_clock),
    .reset(line_1674_reset),
    .valid(line_1674_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1675)) line_1675 (
    .clock(line_1675_clock),
    .reset(line_1675_reset),
    .valid(line_1675_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1676)) line_1676 (
    .clock(line_1676_clock),
    .reset(line_1676_reset),
    .valid(line_1676_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1677)) line_1677 (
    .clock(line_1677_clock),
    .reset(line_1677_reset),
    .valid(line_1677_valid)
  );
  assign line_1661_clock = clock;
  assign line_1661_reset = reset;
  assign line_1661_valid = _T_12 ^ line_1661_valid_reg;
  assign line_1662_clock = clock;
  assign line_1662_reset = reset;
  assign line_1662_valid = _T_13 ^ line_1662_valid_reg;
  assign line_1663_clock = clock;
  assign line_1663_reset = reset;
  assign line_1663_valid = ~inflightSrc ^ line_1663_valid_reg;
  assign line_1664_clock = clock;
  assign line_1664_reset = reset;
  assign line_1664_valid = inflightSrc ^ line_1664_valid_reg;
  assign line_1665_clock = clock;
  assign line_1665_reset = reset;
  assign line_1665_valid = ~inflightSrc ^ line_1665_valid_reg;
  assign line_1666_clock = clock;
  assign line_1666_reset = reset;
  assign line_1666_valid = inflightSrc ^ line_1666_valid_reg;
  assign line_1667_clock = clock;
  assign line_1667_reset = reset;
  assign line_1667_valid = _T_14 ^ line_1667_valid_reg;
  assign line_1668_clock = clock;
  assign line_1668_reset = reset;
  assign line_1668_valid = _T_15 ^ line_1668_valid_reg;
  assign line_1669_clock = clock;
  assign line_1669_reset = reset;
  assign line_1669_valid = _T_4 ^ line_1669_valid_reg;
  assign line_1670_clock = clock;
  assign line_1670_reset = reset;
  assign line_1670_valid = _T_4 ^ line_1670_valid_reg;
  assign line_1671_clock = clock;
  assign line_1671_reset = reset;
  assign line_1671_valid = _T_23 ^ line_1671_valid_reg;
  assign line_1672_clock = clock;
  assign line_1672_reset = reset;
  assign line_1672_valid = _T_14 ^ line_1672_valid_reg;
  assign line_1673_clock = clock;
  assign line_1673_reset = reset;
  assign line_1673_valid = _T_24 ^ line_1673_valid_reg;
  assign line_1674_clock = clock;
  assign line_1674_reset = reset;
  assign line_1674_valid = _T_27 ^ line_1674_valid_reg;
  assign line_1675_clock = clock;
  assign line_1675_reset = reset;
  assign line_1675_valid = _T_24 ^ line_1675_valid_reg;
  assign line_1676_clock = clock;
  assign line_1676_reset = reset;
  assign line_1676_valid = _T_28 ^ line_1676_valid_reg;
  assign line_1677_clock = clock;
  assign line_1677_reset = reset;
  assign line_1677_valid = _T_25 ^ line_1677_valid_reg;
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_21;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_26;
    end
    line_1661_valid_reg <= _T_12;
    line_1662_valid_reg <= _T_13;
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    line_1663_valid_reg <= ~inflightSrc;
    line_1664_valid_reg <= inflightSrc;
    line_1665_valid_reg <= ~inflightSrc;
    line_1666_valid_reg <= inflightSrc;
    line_1667_valid_reg <= _T_14;
    line_1668_valid_reg <= _T_15;
    line_1669_valid_reg <= _T_4;
    line_1670_valid_reg <= _T_4;
    line_1671_valid_reg <= _T_23;
    line_1672_valid_reg <= _T_14;
    line_1673_valid_reg <= _T_24;
    line_1674_valid_reg <= _T_27;
    line_1675_valid_reg <= _T_24;
    line_1676_valid_reg <= _T_28;
    line_1677_valid_reg <= _T_25;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_1661_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1662_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  inflightSrc = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1663_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1664_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1665_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1666_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1667_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1668_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1669_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1670_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1671_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1672_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1673_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1674_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1675_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1676_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1677_valid_reg = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_12) begin
      cover(1'h1);
    end
    //
    if (_T_12 & _T_13) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (~inflightSrc) begin
      cover(1'h1);
    end
    //
    if (inflightSrc) begin
      cover(1'h1);
    end
    //
    if (~inflightSrc) begin
      cover(1'h1);
    end
    //
    if (inflightSrc) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_4) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _T_15 & _T_5 & _T_23) begin
      cover(1'h1);
    end
    //
    if (~_T_14) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & _T_24 & _T_27) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28) begin
      cover(1'h1);
    end
    //
    if (~_T_14 & ~_T_24 & _T_28 & _T_25) begin
      cover(1'h1);
    end
  end
endmodule
module AXI42SimpleBusConverter(
  input   clock,
  input   reset,
  input   io_out_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
  output  io_out_req_valid // @[src/main/scala/bus/simplebus/ToAXI4.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  _T_4 = io_out_req_ready & io_out_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1678_clock;
  wire  line_1678_reset;
  wire  line_1678_valid;
  reg  line_1678_valid_reg;
  wire  _T_28 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 137:32]
  wire  line_1679_clock;
  wire  line_1679_reset;
  wire  line_1679_valid;
  reg  line_1679_valid_reg;
  wire  _T_29 = ~_T_4; // @[src/main/scala/bus/simplebus/ToAXI4.scala 137:32]
  wire  line_1680_clock;
  wire  line_1680_reset;
  wire  line_1680_valid;
  reg  line_1680_valid_reg;
  wire  line_1681_clock;
  wire  line_1681_reset;
  wire  line_1681_valid;
  reg  line_1681_valid_reg;
  wire  line_1682_clock;
  wire  line_1682_reset;
  wire  line_1682_valid;
  reg  line_1682_valid_reg;
  wire  line_1683_clock;
  wire  line_1683_reset;
  wire  line_1683_valid;
  reg  line_1683_valid_reg;
  wire  line_1684_clock;
  wire  line_1684_reset;
  wire  line_1684_valid;
  reg  line_1684_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1678)) line_1678 (
    .clock(line_1678_clock),
    .reset(line_1678_reset),
    .valid(line_1678_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1679)) line_1679 (
    .clock(line_1679_clock),
    .reset(line_1679_reset),
    .valid(line_1679_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1680)) line_1680 (
    .clock(line_1680_clock),
    .reset(line_1680_reset),
    .valid(line_1680_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1681)) line_1681 (
    .clock(line_1681_clock),
    .reset(line_1681_reset),
    .valid(line_1681_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1682)) line_1682 (
    .clock(line_1682_clock),
    .reset(line_1682_reset),
    .valid(line_1682_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1683)) line_1683 (
    .clock(line_1683_clock),
    .reset(line_1683_reset),
    .valid(line_1683_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1684)) line_1684 (
    .clock(line_1684_clock),
    .reset(line_1684_reset),
    .valid(line_1684_valid)
  );
  assign line_1678_clock = clock;
  assign line_1678_reset = reset;
  assign line_1678_valid = _T_4 ^ line_1678_valid_reg;
  assign line_1679_clock = clock;
  assign line_1679_reset = reset;
  assign line_1679_valid = _T_28 ^ line_1679_valid_reg;
  assign line_1680_clock = clock;
  assign line_1680_reset = reset;
  assign line_1680_valid = _T_29 ^ line_1680_valid_reg;
  assign line_1681_clock = clock;
  assign line_1681_reset = reset;
  assign line_1681_valid = _T_28 ^ line_1681_valid_reg;
  assign line_1682_clock = clock;
  assign line_1682_reset = reset;
  assign line_1682_valid = _T_28 ^ line_1682_valid_reg;
  assign line_1683_clock = clock;
  assign line_1683_reset = reset;
  assign line_1683_valid = _T_28 ^ line_1683_valid_reg;
  assign line_1684_clock = clock;
  assign line_1684_reset = reset;
  assign line_1684_valid = _T_28 ^ line_1684_valid_reg;
  assign io_out_req_valid = 1'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 127:52]
  always @(posedge clock) begin
    line_1678_valid_reg <= _T_4;
    line_1679_valid_reg <= _T_28;
    line_1680_valid_reg <= _T_29;
    line_1681_valid_reg <= _T_28;
    line_1682_valid_reg <= _T_28;
    line_1683_valid_reg <= _T_28;
    line_1684_valid_reg <= _T_28;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1678_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1679_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1680_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1681_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1682_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1683_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1684_valid_reg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2MemPortConverter(
  input   clock,
  input   reset
);
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusAddressMapper(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1685_clock;
  wire  line_1685_reset;
  wire  line_1685_valid;
  reg  line_1685_valid_reg;
  wire [2:0] _io_out_ar_bits_len_T_1 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:30]
  wire  _io_out_w_bits_last_T = io_in_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _io_out_w_bits_last_T_1 = io_in_req_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [2:0] _io_in_resp_bits_cmd_T = io_out_r_bits_last ? 3'h6 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:28]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1686_clock;
  wire  line_1686_reset;
  wire  line_1686_valid;
  reg  line_1686_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 & io_out_w_bits_last | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1687_clock;
  wire  line_1687_reset;
  wire  line_1687_valid;
  reg  line_1687_valid_reg;
  wire  _wAck_T_1 = _wSend_T_1 & io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 188:41]
  wire  line_1688_clock;
  wire  line_1688_reset;
  wire  line_1688_valid;
  reg  line_1688_valid_reg;
  wire  _GEN_9 = _wAck_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1689_clock;
  wire  line_1689_reset;
  wire  line_1689_valid;
  reg  line_1689_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1690_clock;
  wire  line_1690_reset;
  wire  line_1690_valid;
  reg  line_1690_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1685)) line_1685 (
    .clock(line_1685_clock),
    .reset(line_1685_reset),
    .valid(line_1685_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1686)) line_1686 (
    .clock(line_1686_clock),
    .reset(line_1686_reset),
    .valid(line_1686_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1687)) line_1687 (
    .clock(line_1687_clock),
    .reset(line_1687_reset),
    .valid(line_1687_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1688)) line_1688 (
    .clock(line_1688_clock),
    .reset(line_1688_reset),
    .valid(line_1688_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1689)) line_1689 (
    .clock(line_1689_clock),
    .reset(line_1689_reset),
    .valid(line_1689_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1690)) line_1690 (
    .clock(line_1690_clock),
    .reset(line_1690_reset),
    .valid(line_1690_valid)
  );
  assign line_1685_clock = clock;
  assign line_1685_reset = reset;
  assign line_1685_valid = _T_2 ^ line_1685_valid_reg;
  assign line_1686_clock = clock;
  assign line_1686_reset = reset;
  assign line_1686_valid = _awAck_T ^ line_1686_valid_reg;
  assign line_1687_clock = clock;
  assign line_1687_reset = reset;
  assign line_1687_valid = wSend ^ line_1687_valid_reg;
  assign line_1688_clock = clock;
  assign line_1688_reset = reset;
  assign line_1688_valid = _wAck_T_1 ^ line_1688_valid_reg;
  assign line_1689_clock = clock;
  assign line_1689_reset = reset;
  assign line_1689_valid = wSend ^ line_1689_valid_reg;
  assign line_1690_clock = clock;
  assign line_1690_reset = reset;
  assign line_1690_valid = _wen_T_1 ^ line_1690_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : 1'h1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _io_in_resp_bits_cmd_T}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_w_bits_last = _io_out_w_bits_last_T | _io_out_w_bits_last_T_1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 177:54]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_ar_bits_len = {{5'd0}, _io_out_ar_bits_len_T_1}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:24]
  assign io_out_ar_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 170:24]
  always @(posedge clock) begin
    line_1685_valid_reg <= _T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1686_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1687_valid_reg <= wSend;
    line_1688_valid_reg <= _wAck_T_1;
    line_1689_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1690_valid_reg <= _wen_T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1685_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  awAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1686_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wAck = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1687_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1688_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1689_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1690_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wAck_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_out_2_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h80000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [2:0] _outSelVec_enc_T = outMatchVec_2 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _outSelVec_enc_T_1 = outMatchVec_1 ? 3'h2 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] outSelVec_enc = outMatchVec_0 ? 3'h1 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  line_1691_clock;
  wire  line_1691_reset;
  wire  line_1691_valid;
  reg  line_1691_valid_reg;
  wire [2:0] _reqInvalidAddr_T = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
  wire  line_1692_clock;
  wire  line_1692_reset;
  wire  line_1692_valid;
  reg  line_1692_valid_reg;
  wire  _T_3 = ~(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
  wire  line_1693_clock;
  wire  line_1693_reset;
  wire  line_1693_valid;
  reg  line_1693_valid_reg;
  wire  _T_4 = 2'h0 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1694_clock;
  wire  line_1694_reset;
  wire  line_1694_valid;
  reg  line_1694_valid_reg;
  wire  line_1695_clock;
  wire  line_1695_reset;
  wire  line_1695_valid;
  reg  line_1695_valid_reg;
  wire  line_1696_clock;
  wire  line_1696_reset;
  wire  line_1696_valid;
  reg  line_1696_valid_reg;
  wire  line_1697_clock;
  wire  line_1697_reset;
  wire  line_1697_valid;
  reg  line_1697_valid_reg;
  wire  _T_6 = 2'h1 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1698_clock;
  wire  line_1698_reset;
  wire  line_1698_valid;
  reg  line_1698_valid_reg;
  wire  line_1699_clock;
  wire  line_1699_reset;
  wire  line_1699_valid;
  reg  line_1699_valid_reg;
  wire [1:0] _GEN_17 = io_in_resp_valid ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  line_1700_clock;
  wire  line_1700_reset;
  wire  line_1700_valid;
  reg  line_1700_valid_reg;
  wire  _T_8 = 2'h2 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1701_clock;
  wire  line_1701_reset;
  wire  line_1701_valid;
  reg  line_1701_valid_reg;
  wire  line_1702_clock;
  wire  line_1702_reset;
  wire  line_1702_valid;
  reg  line_1702_valid_reg;
  wire  _io_in_req_ready_T_4 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_4 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_5 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_6 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_7 = outSelRespVec_2 ? io_out_2_resp_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_8 = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  GEN_w1_line #(.COVER_INDEX(1691)) line_1691 (
    .clock(line_1691_clock),
    .reset(line_1691_reset),
    .valid(line_1691_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1692)) line_1692 (
    .clock(line_1692_clock),
    .reset(line_1692_reset),
    .valid(line_1692_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1693)) line_1693 (
    .clock(line_1693_clock),
    .reset(line_1693_reset),
    .valid(line_1693_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1694)) line_1694 (
    .clock(line_1694_clock),
    .reset(line_1694_reset),
    .valid(line_1694_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1695)) line_1695 (
    .clock(line_1695_clock),
    .reset(line_1695_reset),
    .valid(line_1695_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1696)) line_1696 (
    .clock(line_1696_clock),
    .reset(line_1696_reset),
    .valid(line_1696_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1697)) line_1697 (
    .clock(line_1697_clock),
    .reset(line_1697_reset),
    .valid(line_1697_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1698)) line_1698 (
    .clock(line_1698_clock),
    .reset(line_1698_reset),
    .valid(line_1698_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1699)) line_1699 (
    .clock(line_1699_clock),
    .reset(line_1699_reset),
    .valid(line_1699_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1700)) line_1700 (
    .clock(line_1700_clock),
    .reset(line_1700_reset),
    .valid(line_1700_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1701)) line_1701 (
    .clock(line_1701_clock),
    .reset(line_1701_reset),
    .valid(line_1701_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1702)) line_1702 (
    .clock(line_1702_clock),
    .reset(line_1702_reset),
    .valid(line_1702_valid)
  );
  assign line_1691_clock = clock;
  assign line_1691_reset = reset;
  assign line_1691_valid = _outSelRespVec_T_2 ^ line_1691_valid_reg;
  assign line_1692_clock = clock;
  assign line_1692_reset = reset;
  assign line_1692_valid = _T_2 ^ line_1692_valid_reg;
  assign line_1693_clock = clock;
  assign line_1693_reset = reset;
  assign line_1693_valid = _T_3 ^ line_1693_valid_reg;
  assign line_1694_clock = clock;
  assign line_1694_reset = reset;
  assign line_1694_valid = _T_4 ^ line_1694_valid_reg;
  assign line_1695_clock = clock;
  assign line_1695_reset = reset;
  assign line_1695_valid = _outSelRespVec_T ^ line_1695_valid_reg;
  assign line_1696_clock = clock;
  assign line_1696_reset = reset;
  assign line_1696_valid = reqInvalidAddr ^ line_1696_valid_reg;
  assign line_1697_clock = clock;
  assign line_1697_reset = reset;
  assign line_1697_valid = _T_4 ^ line_1697_valid_reg;
  assign line_1698_clock = clock;
  assign line_1698_reset = reset;
  assign line_1698_valid = _T_6 ^ line_1698_valid_reg;
  assign line_1699_clock = clock;
  assign line_1699_reset = reset;
  assign line_1699_valid = io_in_resp_valid ^ line_1699_valid_reg;
  assign line_1700_clock = clock;
  assign line_1700_reset = reset;
  assign line_1700_valid = _T_6 ^ line_1700_valid_reg;
  assign line_1701_clock = clock;
  assign line_1701_reset = reset;
  assign line_1701_valid = _T_8 ^ line_1701_valid_reg;
  assign line_1702_clock = clock;
  assign line_1702_reset = reset;
  assign line_1702_valid = io_in_resp_valid ^ line_1702_valid_reg;
  assign io_in_req_ready = _io_in_req_ready_T_4 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_4 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_8 | _io_in_resp_bits_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_3 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_17;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_17;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    line_1691_valid_reg <= _outSelRespVec_T_2;
    line_1692_valid_reg <= _T_2;
    line_1693_valid_reg <= _T_3;
    line_1694_valid_reg <= _T_4;
    line_1695_valid_reg <= _outSelRespVec_T;
    line_1696_valid_reg <= reqInvalidAddr;
    line_1697_valid_reg <= _T_4;
    line_1698_valid_reg <= _T_6;
    line_1699_valid_reg <= io_in_resp_valid;
    line_1700_valid_reg <= _T_6;
    line_1701_valid_reg <= _T_8;
    line_1702_valid_reg <= io_in_resp_valid;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1691_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1692_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1693_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1694_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1695_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1696_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1697_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1698_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1699_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1700_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1701_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1702_valid_reg = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_outSelRespVec_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _outSelRespVec_T) begin
      cover(1'h1);
    end
    //
    if (_T_4 & reqInvalidAddr) begin
      cover(1'h1);
    end
    //
    if (~_T_4) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_6 & io_in_resp_valid) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6 & _T_8) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6 & _T_8 & io_in_resp_valid) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_mtip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_msip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         isWFI_0,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _fullMask_T_8 = io__in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_9 = io__in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_10 = io__in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_11 = io__in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_12 = io__in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_13 = io__in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_14 = io__in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_15 = io__in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] fullMask = {_fullMask_T_15,_fullMask_T_14,_fullMask_T_13,_fullMask_T_12,_fullMask_T_11,_fullMask_T_10,
    _fullMask_T_9,_fullMask_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1703_clock;
  wire  line_1703_reset;
  wire  line_1703_valid;
  reg  line_1703_valid_reg;
  wire  _GEN_15 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1704_clock;
  wire  line_1704_reset;
  wire  line_1704_valid;
  reg  line_1704_valid_reg;
  wire  _GEN_16 = _r_busy_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1705_clock;
  wire  line_1705_reset;
  wire  line_1705_valid;
  reg  line_1705_valid_reg;
  wire  _GEN_17 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1706_clock;
  wire  line_1706_reset;
  wire  line_1706_valid;
  reg  line_1706_valid_reg;
  wire  _GEN_18 = _io_in_r_valid_T_2 | _GEN_17; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1707_clock;
  wire  line_1707_reset;
  wire  line_1707_valid;
  reg  line_1707_valid_reg;
  wire  _GEN_19 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1708_clock;
  wire  line_1708_reset;
  wire  line_1708_valid;
  reg  line_1708_valid_reg;
  wire  _GEN_20 = _w_busy_T | _GEN_19; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1709_clock;
  wire  line_1709_reset;
  wire  line_1709_valid;
  reg  line_1709_valid_reg;
  wire  _GEN_21 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1710_clock;
  wire  line_1710_reset;
  wire  line_1710_valid;
  reg  line_1710_valid_reg;
  wire  _GEN_22 = _io_in_b_valid_T | _GEN_21; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  reg [63:0] freq_reg; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire [15:0] freq = freq_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 38:22]
  reg [63:0] inc_reg; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire [15:0] inc = inc_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 40:20]
  reg [15:0] cnt; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[src/main/scala/device/AXI4CLINT.scala 43:21]
  wire  tick = nextCnt == freq; // @[src/main/scala/device/AXI4CLINT.scala 45:23]
  wire  line_1711_clock;
  wire  line_1711_reset;
  wire  line_1711_valid;
  reg  line_1711_valid_reg;
  wire [63:0] _GEN_30 = {{48'd0}, inc}; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_1 = mtime + _GEN_30; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire  line_1712_clock;
  wire  line_1712_reset;
  wire  line_1712_valid;
  reg  line_1712_valid_reg;
  wire [63:0] _mtime_T_3 = mtime + 64'h186a0; // @[src/main/scala/device/AXI4CLINT.scala 51:35]
  wire  _io_in_r_bits_data_T = 16'h0 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 16'h8000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 16'hbff8 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 16'h8008 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_4 = 16'h4000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T ? msip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_1 ? freq_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_2 ? mtime : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_8 = _io_in_r_bits_data_T_3 ? inc_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_4 ? mtimecmp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_5 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_11 = _io_in_r_bits_data_T_10 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_12 = _io_in_r_bits_data_T_11 | _io_in_r_bits_data_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_21 = _io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h0; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1713_clock;
  wire  line_1713_reset;
  wire  line_1713_valid;
  reg  line_1713_valid_reg;
  wire [63:0] _msip_T = io__in_w_bits_data & fullMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _msip_T_1 = ~fullMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _msip_T_2 = msip & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _msip_T_3 = _msip_T | _msip_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_23 = _io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8000; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1714_clock;
  wire  line_1714_reset;
  wire  line_1714_valid;
  reg  line_1714_valid_reg;
  wire [63:0] _freq_reg_T_2 = freq_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _freq_reg_T_3 = _msip_T | _freq_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_25 = _io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'hbff8; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1715_clock;
  wire  line_1715_reset;
  wire  line_1715_valid;
  reg  line_1715_valid_reg;
  wire [63:0] _mtime_T_6 = mtime & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtime_T_7 = _msip_T | _mtime_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_27 = _io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8008; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1716_clock;
  wire  line_1716_reset;
  wire  line_1716_valid;
  reg  line_1716_valid_reg;
  wire [63:0] _inc_reg_T_2 = inc_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _inc_reg_T_3 = _msip_T | _inc_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_29 = _io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h4000; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1717_clock;
  wire  line_1717_reset;
  wire  line_1717_valid;
  reg  line_1717_valid_reg;
  wire [63:0] _mtimecmp_T_2 = mtimecmp & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtimecmp_T_3 = _msip_T | _mtimecmp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  reg  io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  GEN_w1_line #(.COVER_INDEX(1703)) line_1703 (
    .clock(line_1703_clock),
    .reset(line_1703_reset),
    .valid(line_1703_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1704)) line_1704 (
    .clock(line_1704_clock),
    .reset(line_1704_reset),
    .valid(line_1704_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1705)) line_1705 (
    .clock(line_1705_clock),
    .reset(line_1705_reset),
    .valid(line_1705_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1706)) line_1706 (
    .clock(line_1706_clock),
    .reset(line_1706_reset),
    .valid(line_1706_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1707)) line_1707 (
    .clock(line_1707_clock),
    .reset(line_1707_reset),
    .valid(line_1707_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1708)) line_1708 (
    .clock(line_1708_clock),
    .reset(line_1708_reset),
    .valid(line_1708_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1709)) line_1709 (
    .clock(line_1709_clock),
    .reset(line_1709_reset),
    .valid(line_1709_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1710)) line_1710 (
    .clock(line_1710_clock),
    .reset(line_1710_reset),
    .valid(line_1710_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1711)) line_1711 (
    .clock(line_1711_clock),
    .reset(line_1711_reset),
    .valid(line_1711_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1712)) line_1712 (
    .clock(line_1712_clock),
    .reset(line_1712_reset),
    .valid(line_1712_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1713)) line_1713 (
    .clock(line_1713_clock),
    .reset(line_1713_reset),
    .valid(line_1713_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1714)) line_1714 (
    .clock(line_1714_clock),
    .reset(line_1714_reset),
    .valid(line_1714_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1715)) line_1715 (
    .clock(line_1715_clock),
    .reset(line_1715_reset),
    .valid(line_1715_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1716)) line_1716 (
    .clock(line_1716_clock),
    .reset(line_1716_reset),
    .valid(line_1716_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1717)) line_1717 (
    .clock(line_1717_clock),
    .reset(line_1717_reset),
    .valid(line_1717_valid)
  );
  assign line_1703_clock = clock;
  assign line_1703_reset = reset;
  assign line_1703_valid = _r_busy_T_1 ^ line_1703_valid_reg;
  assign line_1704_clock = clock;
  assign line_1704_reset = reset;
  assign line_1704_valid = _r_busy_T ^ line_1704_valid_reg;
  assign line_1705_clock = clock;
  assign line_1705_reset = reset;
  assign line_1705_valid = _r_busy_T_1 ^ line_1705_valid_reg;
  assign line_1706_clock = clock;
  assign line_1706_reset = reset;
  assign line_1706_valid = _io_in_r_valid_T_2 ^ line_1706_valid_reg;
  assign line_1707_clock = clock;
  assign line_1707_reset = reset;
  assign line_1707_valid = _w_busy_T_1 ^ line_1707_valid_reg;
  assign line_1708_clock = clock;
  assign line_1708_reset = reset;
  assign line_1708_valid = _w_busy_T ^ line_1708_valid_reg;
  assign line_1709_clock = clock;
  assign line_1709_reset = reset;
  assign line_1709_valid = _w_busy_T_1 ^ line_1709_valid_reg;
  assign line_1710_clock = clock;
  assign line_1710_reset = reset;
  assign line_1710_valid = _io_in_b_valid_T ^ line_1710_valid_reg;
  assign line_1711_clock = clock;
  assign line_1711_reset = reset;
  assign line_1711_valid = tick ^ line_1711_valid_reg;
  assign line_1712_clock = clock;
  assign line_1712_reset = reset;
  assign line_1712_valid = isWFI_0 ^ line_1712_valid_reg;
  assign line_1713_clock = clock;
  assign line_1713_reset = reset;
  assign line_1713_valid = _T_21 ^ line_1713_valid_reg;
  assign line_1714_clock = clock;
  assign line_1714_reset = reset;
  assign line_1714_valid = _T_23 ^ line_1714_valid_reg;
  assign line_1715_clock = clock;
  assign line_1715_reset = reset;
  assign line_1715_valid = _T_25 ^ line_1715_valid_reg;
  assign line_1716_clock = clock;
  assign line_1716_reset = reset;
  assign line_1716_valid = _T_27 ^ line_1716_valid_reg;
  assign line_1717_clock = clock;
  assign line_1717_reset = reset;
  assign line_1717_valid = _T_29 ^ line_1717_valid_reg;
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = _io_in_r_bits_data_T_12 | _io_in_r_bits_data_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__extra_mtip = io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:21]
  assign io__extra_msip = io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_16;
    end
    line_1703_valid_reg <= _r_busy_T_1;
    line_1704_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_18;
    end
    line_1705_valid_reg <= _r_busy_T_1;
    line_1706_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_20;
    end
    line_1707_valid_reg <= _w_busy_T_1;
    line_1708_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_22;
    end
    line_1709_valid_reg <= _w_busy_T_1;
    line_1710_valid_reg <= _io_in_b_valid_T;
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'hbff8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtime <= _mtime_T_7; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (isWFI_0) begin // @[src/main/scala/device/AXI4CLINT.scala 51:18]
      mtime <= _mtime_T_3; // @[src/main/scala/device/AXI4CLINT.scala 51:26]
    end else if (tick) begin // @[src/main/scala/device/AXI4CLINT.scala 46:15]
      mtime <= _mtime_T_1; // @[src/main/scala/device/AXI4CLINT.scala 46:23]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h4000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtimecmp <= _mtimecmp_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      msip <= _msip_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 37:25]
      freq_reg <= 64'h2710; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      freq_reg <= _freq_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 39:24]
      inc_reg <= 64'h1; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8008) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      inc_reg <= _inc_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 42:20]
      cnt <= 16'h0; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end else if (nextCnt < freq) begin // @[src/main/scala/device/AXI4CLINT.scala 44:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    line_1711_valid_reg <= tick;
    line_1712_valid_reg <= isWFI_0;
    line_1713_valid_reg <= _T_21;
    line_1714_valid_reg <= _T_23;
    line_1715_valid_reg <= _T_25;
    line_1716_valid_reg <= _T_27;
    line_1717_valid_reg <= _T_29;
    io_extra_mtip_REG <= mtime >= mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 66:38]
    io_extra_msip_REG <= msip != 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 67:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1703_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1704_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1705_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1706_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1707_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1708_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1709_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1710_valid_reg = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  mtime = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  mtimecmp = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  msip = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  freq_reg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  inc_reg = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  cnt = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  line_1711_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_1712_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_1713_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_1714_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_1715_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_1716_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_1717_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_extra_mtip_REG = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  io_extra_msip_REG = _RAND_27[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (tick) begin
      cover(1'h1);
    end
    //
    if (isWFI_0) begin
      cover(1'h1);
    end
    //
    if (_T_21) begin
      cover(1'h1);
    end
    //
    if (_T_23) begin
      cover(1'h1);
    end
    //
    if (_T_25) begin
      cover(1'h1);
    end
    //
    if (_T_27) begin
      cover(1'h1);
    end
    //
    if (_T_29) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1718_clock;
  wire  line_1718_reset;
  wire  line_1718_valid;
  reg  line_1718_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1719_clock;
  wire  line_1719_reset;
  wire  line_1719_valid;
  reg  line_1719_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1720_clock;
  wire  line_1720_reset;
  wire  line_1720_valid;
  reg  line_1720_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1721_clock;
  wire  line_1721_reset;
  wire  line_1721_valid;
  reg  line_1721_valid_reg;
  wire  line_1722_clock;
  wire  line_1722_reset;
  wire  line_1722_valid;
  reg  line_1722_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1723_clock;
  wire  line_1723_reset;
  wire  line_1723_valid;
  reg  line_1723_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1724_clock;
  wire  line_1724_reset;
  wire  line_1724_valid;
  reg  line_1724_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1718)) line_1718 (
    .clock(line_1718_clock),
    .reset(line_1718_reset),
    .valid(line_1718_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1719)) line_1719 (
    .clock(line_1719_clock),
    .reset(line_1719_reset),
    .valid(line_1719_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1720)) line_1720 (
    .clock(line_1720_clock),
    .reset(line_1720_reset),
    .valid(line_1720_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1721)) line_1721 (
    .clock(line_1721_clock),
    .reset(line_1721_reset),
    .valid(line_1721_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1722)) line_1722 (
    .clock(line_1722_clock),
    .reset(line_1722_reset),
    .valid(line_1722_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1723)) line_1723 (
    .clock(line_1723_clock),
    .reset(line_1723_reset),
    .valid(line_1723_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1724)) line_1724 (
    .clock(line_1724_clock),
    .reset(line_1724_reset),
    .valid(line_1724_valid)
  );
  assign line_1718_clock = clock;
  assign line_1718_reset = reset;
  assign line_1718_valid = _T_2 ^ line_1718_valid_reg;
  assign line_1719_clock = clock;
  assign line_1719_reset = reset;
  assign line_1719_valid = _T_3 ^ line_1719_valid_reg;
  assign line_1720_clock = clock;
  assign line_1720_reset = reset;
  assign line_1720_valid = _awAck_T ^ line_1720_valid_reg;
  assign line_1721_clock = clock;
  assign line_1721_reset = reset;
  assign line_1721_valid = wSend ^ line_1721_valid_reg;
  assign line_1722_clock = clock;
  assign line_1722_reset = reset;
  assign line_1722_valid = _wSend_T_1 ^ line_1722_valid_reg;
  assign line_1723_clock = clock;
  assign line_1723_reset = reset;
  assign line_1723_valid = wSend ^ line_1723_valid_reg;
  assign line_1724_clock = clock;
  assign line_1724_reset = reset;
  assign line_1724_valid = _wen_T_1 ^ line_1724_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1718_valid_reg <= _T_2;
    line_1719_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1720_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1721_valid_reg <= wSend;
    line_1722_valid_reg <= _wSend_T_1;
    line_1723_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1724_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1718_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1719_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1720_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1721_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1722_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1723_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1724_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_meip_0, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1725_clock;
  wire  line_1725_reset;
  wire  line_1725_valid;
  reg  line_1725_valid_reg;
  wire  _GEN_19 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1726_clock;
  wire  line_1726_reset;
  wire  line_1726_valid;
  reg  line_1726_valid_reg;
  wire  _GEN_20 = _r_busy_T | _GEN_19; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1727_clock;
  wire  line_1727_reset;
  wire  line_1727_valid;
  reg  line_1727_valid_reg;
  wire  _GEN_21 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1728_clock;
  wire  line_1728_reset;
  wire  line_1728_valid;
  reg  line_1728_valid_reg;
  wire  _GEN_22 = _io_in_r_valid_T_2 | _GEN_21; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1729_clock;
  wire  line_1729_reset;
  wire  line_1729_valid;
  reg  line_1729_valid_reg;
  wire  _GEN_23 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1730_clock;
  wire  line_1730_reset;
  wire  line_1730_valid;
  reg  line_1730_valid_reg;
  wire  _GEN_24 = _w_busy_T | _GEN_23; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1731_clock;
  wire  line_1731_reset;
  wire  line_1731_valid;
  reg  line_1731_valid_reg;
  wire  _GEN_25 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1732_clock;
  wire  line_1732_reset;
  wire  line_1732_valid;
  reg  line_1732_valid_reg;
  wire  _GEN_26 = _io_in_b_valid_T | _GEN_25; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  reg [31:0] enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  wire  _T_4 = _r_busy_T_1 & io__in_ar_bits_addr[25:0] == 26'h200004; // @[src/main/scala/device/AXI4PLIC.scala 68:25]
  wire  line_1733_clock;
  wire  line_1733_reset;
  wire  line_1733_valid;
  reg  line_1733_valid_reg;
  wire [7:0] _T_12 = io__in_w_bits_strb >> io__in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4PLIC.scala 89:85]
  wire [7:0] _T_21 = _T_12[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_22 = _T_12[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_23 = _T_12[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_24 = _T_12[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_25 = _T_12[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_26 = _T_12[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_27 = _T_12[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_28 = _T_12[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_29 = {_T_28,_T_27,_T_26,_T_25,_T_24,_T_23,_T_22,_T_21}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T_1 = 26'h2000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 26'h4 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 26'h200000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_6 = _rdata_T_1 ? enable_0_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_8 = _rdata_T_3 ? priority_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_9 = _rdata_T_4 ? threshold_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_6 | _rdata_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] rdata = _rdata_T_12 | _rdata_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_32 = _io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h2000; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1734_clock;
  wire  line_1734_reset;
  wire  line_1734_valid;
  reg  line_1734_valid_reg;
  wire [31:0] _enable_0_0_T = io__in_w_bits_data[31:0] & _T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _enable_0_0_T_1 = ~_T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _enable_0_0_T_2 = enable_0_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _enable_0_0_T_3 = _enable_0_0_T | _enable_0_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_34 = _io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200004; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1735_clock;
  wire  line_1735_reset;
  wire  line_1735_valid;
  reg  line_1735_valid_reg;
  wire  _GEN_14 = ~_enable_0_0_T[0]; // @[src/main/scala/device/AXI4PLIC.scala 60:27]
  wire  line_1736_clock;
  wire  line_1736_reset;
  wire  line_1736_valid;
  reg  line_1736_valid_reg;
  wire  line_1737_clock;
  wire  line_1737_reset;
  wire  line_1737_valid;
  reg  line_1737_valid_reg;
  wire  _T_36 = _io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h4; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1738_clock;
  wire  line_1738_reset;
  wire  line_1738_valid;
  reg  line_1738_valid_reg;
  wire [31:0] _priority_0_T_2 = priority_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _priority_0_T_3 = _enable_0_0_T | _priority_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_38 = _io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200000; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1739_clock;
  wire  line_1739_reset;
  wire  line_1739_valid;
  reg  line_1739_valid_reg;
  wire [31:0] _threshold_0_T_2 = threshold_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _threshold_0_T_3 = _enable_0_0_T | _threshold_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  GEN_w1_line #(.COVER_INDEX(1725)) line_1725 (
    .clock(line_1725_clock),
    .reset(line_1725_reset),
    .valid(line_1725_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1726)) line_1726 (
    .clock(line_1726_clock),
    .reset(line_1726_reset),
    .valid(line_1726_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1727)) line_1727 (
    .clock(line_1727_clock),
    .reset(line_1727_reset),
    .valid(line_1727_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1728)) line_1728 (
    .clock(line_1728_clock),
    .reset(line_1728_reset),
    .valid(line_1728_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1729)) line_1729 (
    .clock(line_1729_clock),
    .reset(line_1729_reset),
    .valid(line_1729_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1730)) line_1730 (
    .clock(line_1730_clock),
    .reset(line_1730_reset),
    .valid(line_1730_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1731)) line_1731 (
    .clock(line_1731_clock),
    .reset(line_1731_reset),
    .valid(line_1731_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1732)) line_1732 (
    .clock(line_1732_clock),
    .reset(line_1732_reset),
    .valid(line_1732_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1733)) line_1733 (
    .clock(line_1733_clock),
    .reset(line_1733_reset),
    .valid(line_1733_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1734)) line_1734 (
    .clock(line_1734_clock),
    .reset(line_1734_reset),
    .valid(line_1734_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1735)) line_1735 (
    .clock(line_1735_clock),
    .reset(line_1735_reset),
    .valid(line_1735_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1736)) line_1736 (
    .clock(line_1736_clock),
    .reset(line_1736_reset),
    .valid(line_1736_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1737)) line_1737 (
    .clock(line_1737_clock),
    .reset(line_1737_reset),
    .valid(line_1737_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1738)) line_1738 (
    .clock(line_1738_clock),
    .reset(line_1738_reset),
    .valid(line_1738_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1739)) line_1739 (
    .clock(line_1739_clock),
    .reset(line_1739_reset),
    .valid(line_1739_valid)
  );
  assign line_1725_clock = clock;
  assign line_1725_reset = reset;
  assign line_1725_valid = _r_busy_T_1 ^ line_1725_valid_reg;
  assign line_1726_clock = clock;
  assign line_1726_reset = reset;
  assign line_1726_valid = _r_busy_T ^ line_1726_valid_reg;
  assign line_1727_clock = clock;
  assign line_1727_reset = reset;
  assign line_1727_valid = _r_busy_T_1 ^ line_1727_valid_reg;
  assign line_1728_clock = clock;
  assign line_1728_reset = reset;
  assign line_1728_valid = _io_in_r_valid_T_2 ^ line_1728_valid_reg;
  assign line_1729_clock = clock;
  assign line_1729_reset = reset;
  assign line_1729_valid = _w_busy_T_1 ^ line_1729_valid_reg;
  assign line_1730_clock = clock;
  assign line_1730_reset = reset;
  assign line_1730_valid = _w_busy_T ^ line_1730_valid_reg;
  assign line_1731_clock = clock;
  assign line_1731_reset = reset;
  assign line_1731_valid = _w_busy_T_1 ^ line_1731_valid_reg;
  assign line_1732_clock = clock;
  assign line_1732_reset = reset;
  assign line_1732_valid = _io_in_b_valid_T ^ line_1732_valid_reg;
  assign line_1733_clock = clock;
  assign line_1733_reset = reset;
  assign line_1733_valid = _T_4 ^ line_1733_valid_reg;
  assign line_1734_clock = clock;
  assign line_1734_reset = reset;
  assign line_1734_valid = _T_32 ^ line_1734_valid_reg;
  assign line_1735_clock = clock;
  assign line_1735_reset = reset;
  assign line_1735_valid = _T_34 ^ line_1735_valid_reg;
  assign line_1736_clock = clock;
  assign line_1736_reset = reset;
  assign line_1736_valid = ~_enable_0_0_T[0] ^ line_1736_valid_reg;
  assign line_1737_clock = clock;
  assign line_1737_reset = reset;
  assign line_1737_valid = _enable_0_0_T[0] ^ line_1737_valid_reg;
  assign line_1738_clock = clock;
  assign line_1738_reset = reset;
  assign line_1738_valid = _T_36 ^ line_1738_valid_reg;
  assign line_1739_clock = clock;
  assign line_1739_reset = reset;
  assign line_1739_valid = _T_38 ^ line_1739_valid_reg;
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = {rdata,rdata}; // @[src/main/scala/device/AXI4PLIC.scala 91:25]
  assign io__extra_meip_0 = 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_20;
    end
    line_1725_valid_reg <= _r_busy_T_1;
    line_1726_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_22;
    end
    line_1727_valid_reg <= _r_busy_T_1;
    line_1728_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_24;
    end
    line_1729_valid_reg <= _w_busy_T_1;
    line_1730_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_26;
    end
    line_1731_valid_reg <= _w_busy_T_1;
    line_1732_valid_reg <= _io_in_b_valid_T;
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      priority_0 <= _priority_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h2000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      enable_0_0 <= _enable_0_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      threshold_0 <= _threshold_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    line_1733_valid_reg <= _T_4;
    line_1734_valid_reg <= _T_32;
    line_1735_valid_reg <= _T_34;
    line_1736_valid_reg <= ~_enable_0_0_T[0];
    line_1737_valid_reg <= _enable_0_0_T[0];
    line_1738_valid_reg <= _T_36;
    line_1739_valid_reg <= _T_38;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1725_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1726_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1727_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1728_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1729_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1730_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1731_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1732_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  priority_0 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  enable_0_0 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  threshold_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  line_1733_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1734_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1735_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1736_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_1737_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_1738_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_1739_valid_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_32) begin
      cover(1'h1);
    end
    //
    if (_T_34) begin
      cover(1'h1);
    end
    //
    if (_T_34 & _GEN_14) begin
      cover(1'h1);
    end
    //
    if (_T_34 & _enable_0_0_T[0]) begin
      cover(1'h1);
    end
    //
    if (_T_36) begin
      cover(1'h1);
    end
    //
    if (_T_38) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_2(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1740_clock;
  wire  line_1740_reset;
  wire  line_1740_valid;
  reg  line_1740_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1741_clock;
  wire  line_1741_reset;
  wire  line_1741_valid;
  reg  line_1741_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1742_clock;
  wire  line_1742_reset;
  wire  line_1742_valid;
  reg  line_1742_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1743_clock;
  wire  line_1743_reset;
  wire  line_1743_valid;
  reg  line_1743_valid_reg;
  wire  line_1744_clock;
  wire  line_1744_reset;
  wire  line_1744_valid;
  reg  line_1744_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1745_clock;
  wire  line_1745_reset;
  wire  line_1745_valid;
  reg  line_1745_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1746_clock;
  wire  line_1746_reset;
  wire  line_1746_valid;
  reg  line_1746_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1740)) line_1740 (
    .clock(line_1740_clock),
    .reset(line_1740_reset),
    .valid(line_1740_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1741)) line_1741 (
    .clock(line_1741_clock),
    .reset(line_1741_reset),
    .valid(line_1741_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1742)) line_1742 (
    .clock(line_1742_clock),
    .reset(line_1742_reset),
    .valid(line_1742_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1743)) line_1743 (
    .clock(line_1743_clock),
    .reset(line_1743_reset),
    .valid(line_1743_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1744)) line_1744 (
    .clock(line_1744_clock),
    .reset(line_1744_reset),
    .valid(line_1744_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1745)) line_1745 (
    .clock(line_1745_clock),
    .reset(line_1745_reset),
    .valid(line_1745_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1746)) line_1746 (
    .clock(line_1746_clock),
    .reset(line_1746_reset),
    .valid(line_1746_valid)
  );
  assign line_1740_clock = clock;
  assign line_1740_reset = reset;
  assign line_1740_valid = _T_2 ^ line_1740_valid_reg;
  assign line_1741_clock = clock;
  assign line_1741_reset = reset;
  assign line_1741_valid = _T_3 ^ line_1741_valid_reg;
  assign line_1742_clock = clock;
  assign line_1742_reset = reset;
  assign line_1742_valid = _awAck_T ^ line_1742_valid_reg;
  assign line_1743_clock = clock;
  assign line_1743_reset = reset;
  assign line_1743_valid = wSend ^ line_1743_valid_reg;
  assign line_1744_clock = clock;
  assign line_1744_reset = reset;
  assign line_1744_valid = _wSend_T_1 ^ line_1744_valid_reg;
  assign line_1745_clock = clock;
  assign line_1745_reset = reset;
  assign line_1745_valid = wSend ^ line_1745_valid_reg;
  assign line_1746_clock = clock;
  assign line_1746_reset = reset;
  assign line_1746_valid = _wen_T_1 ^ line_1746_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1740_valid_reg <= _T_2;
    line_1741_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1742_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1743_valid_reg <= wSend;
    line_1744_valid_reg <= _wSend_T_1;
    line_1745_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1746_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1740_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1741_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1742_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1743_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1744_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1745_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1746_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_aw_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_aw_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_aw_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_w_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mem_w_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_w_bits_strb, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_b_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_ar_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_ar_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_ar_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mem_ar_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mem_r_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_req_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_req_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_resp_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_resp_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/system/NutShell.scala 45:14]
);
  wire  nutcore_clock; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_reset; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [2:0] nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_isWFI; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  cohMg_clock; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_reset; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  xbar_clock; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_reset; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  axi2sb_clock; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_reset; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  memport_bridge_clock; // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
  wire  memport_bridge_reset; // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
  wire  memAddrMap_clock; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_reset; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_in_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  io_mem_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  clint_clock; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_reset; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [7:0] clint_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_isWFI_0; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] clint_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_clock; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_reset; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [7:0] plic_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] plic_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  NutCore nutcore ( // @[src/main/scala/system/NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_size(nutcore_io_dmem_mem_req_bits_size),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wmask(nutcore_io_dmem_mem_req_bits_wmask),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .isWFI(nutcore_isWFI),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_msip(nutcore_io_extra_msip)
  );
  CoherenceManager cohMg ( // @[src/main/scala/system/NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_2 xbar ( // @[src/main/scala/system/NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[src/main/scala/system/NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid)
  );
  SimpleBus2MemPortConverter memport_bridge ( // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
    .clock(memport_bridge_clock),
    .reset(memport_bridge_reset)
  );
  SimpleBusAddressMapper memAddrMap ( // @[src/main/scala/system/NutShell.scala 93:26]
    .clock(memAddrMap_clock),
    .reset(memAddrMap_reset),
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_size(memAddrMap_io_in_req_bits_size),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(memAddrMap_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_size(memAddrMap_io_out_req_bits_size),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(memAddrMap_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter io_mem_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(io_mem_bridge_clock),
    .reset(io_mem_bridge_reset),
    .io_in_req_ready(io_mem_bridge_io_in_req_ready),
    .io_in_req_valid(io_mem_bridge_io_in_req_valid),
    .io_in_req_bits_addr(io_mem_bridge_io_in_req_bits_addr),
    .io_in_req_bits_size(io_mem_bridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_mem_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_mem_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_mem_bridge_io_in_req_bits_wdata),
    .io_in_resp_valid(io_mem_bridge_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_mem_bridge_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_mem_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(io_mem_bridge_io_out_aw_ready),
    .io_out_aw_valid(io_mem_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(io_mem_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(io_mem_bridge_io_out_w_ready),
    .io_out_w_valid(io_mem_bridge_io_out_w_valid),
    .io_out_w_bits_data(io_mem_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(io_mem_bridge_io_out_w_bits_strb),
    .io_out_w_bits_last(io_mem_bridge_io_out_w_bits_last),
    .io_out_b_valid(io_mem_bridge_io_out_b_valid),
    .io_out_ar_valid(io_mem_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(io_mem_bridge_io_out_ar_bits_addr),
    .io_out_ar_bits_len(io_mem_bridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(io_mem_bridge_io_out_ar_bits_size),
    .io_out_r_valid(io_mem_bridge_io_out_r_valid),
    .io_out_r_bits_data(io_mem_bridge_io_out_r_bits_data),
    .io_out_r_bits_last(io_mem_bridge_io_out_r_bits_last)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[src/main/scala/system/NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_cmd(mmioXbar_io_out_2_resp_bits_cmd),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  AXI4CLINT clint ( // @[src/main/scala/system/NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_aw_ready(clint_io__in_aw_ready),
    .io__in_aw_valid(clint_io__in_aw_valid),
    .io__in_aw_bits_addr(clint_io__in_aw_bits_addr),
    .io__in_w_ready(clint_io__in_w_ready),
    .io__in_w_valid(clint_io__in_w_valid),
    .io__in_w_bits_data(clint_io__in_w_bits_data),
    .io__in_w_bits_strb(clint_io__in_w_bits_strb),
    .io__in_b_ready(clint_io__in_b_ready),
    .io__in_b_valid(clint_io__in_b_valid),
    .io__in_ar_ready(clint_io__in_ar_ready),
    .io__in_ar_valid(clint_io__in_ar_valid),
    .io__in_ar_bits_addr(clint_io__in_ar_bits_addr),
    .io__in_r_ready(clint_io__in_r_ready),
    .io__in_r_valid(clint_io__in_r_valid),
    .io__in_r_bits_data(clint_io__in_r_bits_data),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .isWFI_0(clint_isWFI_0),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_1 clint_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(clint_io_in_bridge_clock),
    .reset(clint_io_in_bridge_reset),
    .io_in_req_ready(clint_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(clint_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(clint_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(clint_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(clint_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(clint_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(clint_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(clint_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(clint_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(clint_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(clint_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(clint_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(clint_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(clint_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(clint_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(clint_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(clint_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(clint_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(clint_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(clint_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(clint_io_in_bridge_io_out_r_bits_data)
  );
  AXI4PLIC plic ( // @[src/main/scala/system/NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_aw_ready(plic_io__in_aw_ready),
    .io__in_aw_valid(plic_io__in_aw_valid),
    .io__in_aw_bits_addr(plic_io__in_aw_bits_addr),
    .io__in_w_ready(plic_io__in_w_ready),
    .io__in_w_valid(plic_io__in_w_valid),
    .io__in_w_bits_data(plic_io__in_w_bits_data),
    .io__in_w_bits_strb(plic_io__in_w_bits_strb),
    .io__in_b_ready(plic_io__in_b_ready),
    .io__in_b_valid(plic_io__in_b_valid),
    .io__in_ar_ready(plic_io__in_ar_ready),
    .io__in_ar_valid(plic_io__in_ar_valid),
    .io__in_ar_bits_addr(plic_io__in_ar_bits_addr),
    .io__in_r_ready(plic_io__in_r_ready),
    .io__in_r_valid(plic_io__in_r_valid),
    .io__in_r_bits_data(plic_io__in_r_bits_data),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_2 plic_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(plic_io_in_bridge_clock),
    .reset(plic_io_in_bridge_reset),
    .io_in_req_ready(plic_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(plic_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(plic_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(plic_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(plic_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(plic_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(plic_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(plic_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(plic_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(plic_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(plic_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(plic_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(plic_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(plic_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(plic_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(plic_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(plic_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(plic_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(plic_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(plic_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(plic_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(plic_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(plic_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(plic_io_in_bridge_io_out_r_bits_data)
  );
  assign io_mem_aw_valid = io_mem_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_addr = io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_valid = io_mem_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_data = io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_strb = io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_last = io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_valid = io_mem_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_addr = io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_len = io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_size = io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mmio_req_valid = mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_resp_ready = mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_out_req_ready = memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_valid = memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[src/main/scala/system/NutShell.scala 63:23]
  assign memport_bridge_clock = clock;
  assign memport_bridge_reset = reset;
  assign memAddrMap_clock = clock;
  assign memAddrMap_reset = reset;
  assign memAddrMap_io_in_req_valid = xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_addr = xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_size = xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_cmd = xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wmask = xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wdata = xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_out_req_ready = io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_clock = clock;
  assign io_mem_bridge_reset = reset;
  assign io_mem_bridge_io_in_req_valid = memAddrMap_io_out_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_size = memAddrMap_io_out_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wmask = memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_out_aw_ready = io_mem_aw_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_w_ready = io_mem_w_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_b_valid = io_mem_b_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_valid = io_mem_r_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_data = io_mem_r_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_last = io_mem_r_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_valid = io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_aw_valid = clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_aw_bits_addr = clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_valid = clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_data = clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_strb = clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_b_ready = clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_valid = clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_bits_addr = clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_r_ready = clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_isWFI_0 = nutcore_isWFI;
  assign clint_io_in_bridge_clock = clock;
  assign clint_io_in_bridge_reset = reset;
  assign clint_io_in_bridge_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_out_aw_ready = clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_w_ready = clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_b_valid = clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_ar_ready = clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_valid = clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_bits_data = clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_aw_valid = plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_aw_bits_addr = plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_valid = plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_data = plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_strb = plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_b_ready = plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_valid = plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_bits_addr = plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_r_ready = plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_clock = clock;
  assign plic_io_in_bridge_reset = reset;
  assign plic_io_in_bridge_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_out_aw_ready = plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_w_ready = plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_b_valid = plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_ar_ready = plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_valid = plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_bits_data = plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module DifftestMem1P(
  input         clock,
  input         reset,
  input         read_valid, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input  [63:0] read_index, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  output [63:0] read_data_0, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input         write_valid, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_index, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_data_0, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_mask_0 // @[difftest/src/main/scala/common/Mem.scala 204:17]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  helper_0_r_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_w_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_mask; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_clock; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  _T_1 = ~reset; // @[difftest/src/main/scala/common/Mem.scala 214:16]
  wire [64:0] _T_3 = read_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 215:26]
  wire [65:0] _T_4 = {{1'd0}, _T_3}; // @[difftest/src/main/scala/common/Mem.scala 215:39]
  wire [64:0] _T_9 = write_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 223:27]
  wire [65:0] _T_10 = {{1'd0}, _T_9}; // @[difftest/src/main/scala/common/Mem.scala 223:40]
  wire  line_1747_clock;
  wire  line_1747_reset;
  wire  line_1747_valid;
  reg  line_1747_valid_reg;
  wire  _T_17 = ~(~read_valid | ~write_valid); // @[difftest/src/main/scala/common/Mem.scala 263:9]
  wire  line_1748_clock;
  wire  line_1748_reset;
  wire  line_1748_valid;
  reg  line_1748_valid_reg;
  MemRWHelper helper_0 ( // @[difftest/src/main/scala/common/Mem.scala 197:49]
    .r_enable(helper_0_r_enable),
    .r_index(helper_0_r_index),
    .r_data(helper_0_r_data),
    .w_enable(helper_0_w_enable),
    .w_index(helper_0_w_index),
    .w_data(helper_0_w_data),
    .w_mask(helper_0_w_mask),
    .clock(helper_0_clock)
  );
  GEN_w1_line #(.COVER_INDEX(1747)) line_1747 (
    .clock(line_1747_clock),
    .reset(line_1747_reset),
    .valid(line_1747_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1748)) line_1748 (
    .clock(line_1748_clock),
    .reset(line_1748_reset),
    .valid(line_1748_valid)
  );
  assign line_1747_clock = clock;
  assign line_1747_reset = reset;
  assign line_1747_valid = _T_1 ^ line_1747_valid_reg;
  assign line_1748_clock = clock;
  assign line_1748_reset = reset;
  assign line_1748_valid = _T_17 ^ line_1748_valid_reg;
  assign read_data_0 = helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 211:13]
  assign helper_0_r_enable = ~reset & read_valid; // @[difftest/src/main/scala/common/Mem.scala 214:30]
  assign helper_0_r_index = _T_4[63:0]; // @[difftest/src/main/scala/common/Mem.scala 102:13]
  assign helper_0_w_enable = _T_1 & write_valid; // @[difftest/src/main/scala/common/Mem.scala 222:30]
  assign helper_0_w_index = _T_10[63:0]; // @[difftest/src/main/scala/common/Mem.scala 150:13]
  assign helper_0_w_data = write_data_0; // @[difftest/src/main/scala/common/Mem.scala 151:12]
  assign helper_0_w_mask = write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 152:12]
  assign helper_0_clock = clock; // @[difftest/src/main/scala/common/Mem.scala 220:13]
  always @(posedge clock) begin
    line_1747_valid_reg <= _T_1;
    line_1748_valid_reg <= _T_17;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~(~read_valid | ~write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed: read and write come at the same cycle\n    at Mem.scala:263 assert(!read.valid || !write.valid, \"read and write come at the same cycle\")\n"
            ); // @[difftest/src/main/scala/common/Mem.scala 263:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1747_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1748_valid_reg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_1 & _T_17) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      assert(~read_valid | ~write_valid); // @[difftest/src/main/scala/common/Mem.scala 263:9]
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_bits_last, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_bits_last // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
`endif // RANDOMIZE_REG_INIT
  wire  rdata_mem_clock; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_reset; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_read_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_write_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [7:0] _fullMask_T_8 = io_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_9 = io_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_10 = io_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_11 = io_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_12 = io_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_13 = io_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_14 = io_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_15 = io_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [31:0] fullMask_lo = {_fullMask_T_11,_fullMask_T_10,_fullMask_T_9,_fullMask_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire [31:0] fullMask_hi = {_fullMask_T_15,_fullMask_T_14,_fullMask_T_13,_fullMask_T_12}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  reg [7:0] c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [7:0] readBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _len_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [7:0] len_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_1749_clock;
  wire  line_1749_reset;
  wire  line_1749_valid;
  reg  line_1749_valid_reg;
  wire [7:0] _GEN_28 = _len_T ? io_in_ar_bits_len : len_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg [1:0] burst_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_1750_clock;
  wire  line_1750_reset;
  wire  line_1750_valid;
  reg  line_1750_valid_reg;
  wire [1:0] _GEN_29 = _len_T ? 2'h2 : burst_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [31:0] _wrapAddr_WIRE = {{24'd0}, io_in_ar_bits_len}; // @[src/main/scala/device/AXI4Slave.scala 45:{69,69}]
  wire [38:0] _GEN_47 = {{7'd0}, _wrapAddr_WIRE}; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T = _GEN_47 << io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T_1 = ~_wrapAddr_T; // @[src/main/scala/device/AXI4Slave.scala 45:42]
  wire [38:0] _GEN_56 = {{7'd0}, io_in_ar_bits_addr}; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  wire [38:0] wrapAddr = _GEN_56 & _wrapAddr_T_1; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  reg [38:0] raddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_1751_clock;
  wire  line_1751_reset;
  wire  line_1751_valid;
  reg  line_1751_valid_reg;
  wire [38:0] _GEN_30 = _len_T ? wrapAddr : raddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  wire  line_1752_clock;
  wire  line_1752_reset;
  wire  line_1752_valid;
  reg  line_1752_valid_reg;
  wire [7:0] _value_T_1 = readBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T_2 = _GEN_29 == 2'h2 & readBeatCnt == _GEN_28; // @[src/main/scala/device/AXI4Slave.scala 50:51]
  wire  line_1753_clock;
  wire  line_1753_reset;
  wire  line_1753_valid;
  reg  line_1753_valid_reg;
  wire [7:0] _GEN_31 = _GEN_29 == 2'h2 & readBeatCnt == _GEN_28 ? 8'h0 : _value_T_1; // @[src/main/scala/device/AXI4Slave.scala 50:{77,93} src/main/scala/chisel3/util/Counter.scala 77:15]
  wire [7:0] _GEN_32 = ren ? _GEN_31 : readBeatCnt; // @[src/main/scala/device/AXI4Slave.scala 48:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_1754_clock;
  wire  line_1754_reset;
  wire  line_1754_valid;
  reg  line_1754_valid_reg;
  wire [7:0] _value_T_3 = c_value + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1755_clock;
  wire  line_1755_reset;
  wire  line_1755_valid;
  reg  line_1755_valid_reg;
  wire  line_1756_clock;
  wire  line_1756_reset;
  wire  line_1756_valid;
  reg  line_1756_valid_reg;
  wire [31:0] _value_T_4 = io_in_ar_bits_addr >> io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 57:45]
  wire [31:0] _value_T_5 = _value_T_4 & _wrapAddr_WIRE; // @[src/main/scala/device/AXI4Slave.scala 57:67]
  wire  _T_5 = io_in_ar_bits_len != 8'h0; // @[src/main/scala/device/AXI4Slave.scala 58:32]
  wire  line_1757_clock;
  wire  line_1757_reset;
  wire  line_1757_valid;
  reg  line_1757_valid_reg;
  wire  _T_11 = io_in_ar_bits_len == 8'h7; // @[src/main/scala/device/AXI4Slave.scala 60:30]
  wire  _T_12 = io_in_ar_bits_len == 8'h1 | io_in_ar_bits_len == 8'h3 | _T_11; // @[src/main/scala/device/AXI4Slave.scala 59:71]
  wire  _T_14 = _T_12 | io_in_ar_bits_len == 8'hf; // @[src/main/scala/device/AXI4Slave.scala 60:38]
  wire  _T_16 = ~reset; // @[src/main/scala/device/AXI4Slave.scala 59:17]
  wire  line_1758_clock;
  wire  line_1758_reset;
  wire  line_1758_valid;
  reg  line_1758_valid_reg;
  wire  _T_17 = ~_T_14; // @[src/main/scala/device/AXI4Slave.scala 59:17]
  wire  line_1759_clock;
  wire  line_1759_reset;
  wire  line_1759_valid;
  reg  line_1759_valid_reg;
  wire [31:0] _GEN_35 = _len_T ? _value_T_5 : {{24'd0}, _GEN_32}; // @[src/main/scala/device/AXI4Slave.scala 56:29 57:23]
  wire  _r_busy_T_2 = io_in_r_valid & io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 70:56]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1760_clock;
  wire  line_1760_reset;
  wire  line_1760_valid;
  reg  line_1760_valid_reg;
  wire  _GEN_36 = _r_busy_T_2 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1761_clock;
  wire  line_1761_reset;
  wire  line_1761_valid;
  reg  line_1761_valid_reg;
  wire  _GEN_37 = _len_T | _GEN_36; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_valid_T_2 = ren & (_len_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1762_clock;
  wire  line_1762_reset;
  wire  line_1762_valid;
  reg  line_1762_valid_reg;
  wire  _GEN_38 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1763_clock;
  wire  line_1763_reset;
  wire  line_1763_valid;
  reg  line_1763_valid_reg;
  wire  _GEN_39 = _io_in_r_valid_T_2 | _GEN_38; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [7:0] writeBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _waddr_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [31:0] waddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_1764_clock;
  wire  line_1764_reset;
  wire  line_1764_valid;
  reg  line_1764_valid_reg;
  wire [31:0] _GEN_40 = _waddr_T ? io_in_aw_bits_addr : waddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  _T_18 = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1765_clock;
  wire  line_1765_reset;
  wire  line_1765_valid;
  reg  line_1765_valid_reg;
  wire [7:0] _value_T_7 = writeBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1766_clock;
  wire  line_1766_reset;
  wire  line_1766_valid;
  reg  line_1766_valid_reg;
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1767_clock;
  wire  line_1767_reset;
  wire  line_1767_valid;
  reg  line_1767_valid_reg;
  wire  _GEN_43 = io_in_b_valid ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1768_clock;
  wire  line_1768_reset;
  wire  line_1768_valid;
  reg  line_1768_valid_reg;
  wire  _GEN_44 = _waddr_T | _GEN_43; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T_1 = _T_18 & io_in_w_bits_last; // @[src/main/scala/device/AXI4Slave.scala 97:43]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1769_clock;
  wire  line_1769_reset;
  wire  line_1769_valid;
  reg  line_1769_valid_reg;
  wire  _GEN_45 = io_in_b_valid ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1770_clock;
  wire  line_1770_reset;
  wire  line_1770_valid;
  reg  line_1770_valid_reg;
  wire  _GEN_46 = _io_in_b_valid_T_1 | _GEN_45; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  line_1771_clock;
  wire  line_1771_reset;
  wire  line_1771_valid;
  reg  line_1771_valid_reg;
  wire  line_1772_clock;
  wire  line_1772_reset;
  wire  line_1772_valid;
  reg  line_1772_valid_reg;
  wire  line_1773_clock;
  wire  line_1773_reset;
  wire  line_1773_valid;
  reg  line_1773_valid_reg;
  wire  line_1774_clock;
  wire  line_1774_reset;
  wire  line_1774_valid;
  reg  line_1774_valid_reg;
  wire [31:0] _wIdx_T = _GEN_40 & 32'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [28:0] _GEN_58 = {{21'd0}, writeBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T[31:3] + _GEN_58; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [38:0] _rIdx_T = _GEN_30 & 39'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [35:0] _GEN_59 = {{28'd0}, readBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [35:0] rIdx = _rIdx_T[38:3] + _GEN_59; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'h10000000; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire  wen = _T_18 & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 37:25]
  wire  line_1775_clock;
  wire  line_1775_reset;
  wire  line_1775_valid;
  reg  line_1775_valid_reg;
  wire [31:0] rdata_lo = {io_in_w_bits_data[31:24],io_in_w_bits_data[23:16],io_in_w_bits_data[15:8],io_in_w_bits_data[7:
    0]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [31:0] rdata_hi = {io_in_w_bits_data[63:56],io_in_w_bits_data[55:48],io_in_w_bits_data[47:40],io_in_w_bits_data[
    39:32]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  reg  rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  reg  rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  reg [63:0] rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire  line_1776_clock;
  wire  line_1776_reset;
  wire  line_1776_valid;
  reg  line_1776_valid_reg;
  wire [63:0] _rdata_T_28_0 = rdata_REG ? rdata_mem_read_data_0 : rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:8]
  wire [31:0] rdata_lo_2 = {_rdata_T_28_0[31:24],_rdata_T_28_0[23:16],_rdata_T_28_0[15:8],_rdata_T_28_0[7:0]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] rdata_hi_2 = {_rdata_T_28_0[63:56],_rdata_T_28_0[55:48],_rdata_T_28_0[47:40],_rdata_T_28_0[39:32]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] _GEN_60 = reset ? 32'h0 : _GEN_35; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  DifftestMem1P rdata_mem ( // @[difftest/src/main/scala/common/Mem.scala 322:36]
    .clock(rdata_mem_clock),
    .reset(rdata_mem_reset),
    .read_valid(rdata_mem_read_valid),
    .read_index(rdata_mem_read_index),
    .read_data_0(rdata_mem_read_data_0),
    .write_valid(rdata_mem_write_valid),
    .write_index(rdata_mem_write_index),
    .write_data_0(rdata_mem_write_data_0),
    .write_mask_0(rdata_mem_write_mask_0)
  );
  GEN_w1_line #(.COVER_INDEX(1749)) line_1749 (
    .clock(line_1749_clock),
    .reset(line_1749_reset),
    .valid(line_1749_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1750)) line_1750 (
    .clock(line_1750_clock),
    .reset(line_1750_reset),
    .valid(line_1750_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1751)) line_1751 (
    .clock(line_1751_clock),
    .reset(line_1751_reset),
    .valid(line_1751_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1752)) line_1752 (
    .clock(line_1752_clock),
    .reset(line_1752_reset),
    .valid(line_1752_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1753)) line_1753 (
    .clock(line_1753_clock),
    .reset(line_1753_reset),
    .valid(line_1753_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1754)) line_1754 (
    .clock(line_1754_clock),
    .reset(line_1754_reset),
    .valid(line_1754_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1755)) line_1755 (
    .clock(line_1755_clock),
    .reset(line_1755_reset),
    .valid(line_1755_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1756)) line_1756 (
    .clock(line_1756_clock),
    .reset(line_1756_reset),
    .valid(line_1756_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1757)) line_1757 (
    .clock(line_1757_clock),
    .reset(line_1757_reset),
    .valid(line_1757_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1758)) line_1758 (
    .clock(line_1758_clock),
    .reset(line_1758_reset),
    .valid(line_1758_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1759)) line_1759 (
    .clock(line_1759_clock),
    .reset(line_1759_reset),
    .valid(line_1759_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1760)) line_1760 (
    .clock(line_1760_clock),
    .reset(line_1760_reset),
    .valid(line_1760_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1761)) line_1761 (
    .clock(line_1761_clock),
    .reset(line_1761_reset),
    .valid(line_1761_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1762)) line_1762 (
    .clock(line_1762_clock),
    .reset(line_1762_reset),
    .valid(line_1762_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1763)) line_1763 (
    .clock(line_1763_clock),
    .reset(line_1763_reset),
    .valid(line_1763_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1764)) line_1764 (
    .clock(line_1764_clock),
    .reset(line_1764_reset),
    .valid(line_1764_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1765)) line_1765 (
    .clock(line_1765_clock),
    .reset(line_1765_reset),
    .valid(line_1765_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1766)) line_1766 (
    .clock(line_1766_clock),
    .reset(line_1766_reset),
    .valid(line_1766_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1767)) line_1767 (
    .clock(line_1767_clock),
    .reset(line_1767_reset),
    .valid(line_1767_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1768)) line_1768 (
    .clock(line_1768_clock),
    .reset(line_1768_reset),
    .valid(line_1768_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1769)) line_1769 (
    .clock(line_1769_clock),
    .reset(line_1769_reset),
    .valid(line_1769_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1770)) line_1770 (
    .clock(line_1770_clock),
    .reset(line_1770_reset),
    .valid(line_1770_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1771)) line_1771 (
    .clock(line_1771_clock),
    .reset(line_1771_reset),
    .valid(line_1771_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1772)) line_1772 (
    .clock(line_1772_clock),
    .reset(line_1772_reset),
    .valid(line_1772_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1773)) line_1773 (
    .clock(line_1773_clock),
    .reset(line_1773_reset),
    .valid(line_1773_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1774)) line_1774 (
    .clock(line_1774_clock),
    .reset(line_1774_reset),
    .valid(line_1774_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1775)) line_1775 (
    .clock(line_1775_clock),
    .reset(line_1775_reset),
    .valid(line_1775_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1776)) line_1776 (
    .clock(line_1776_clock),
    .reset(line_1776_reset),
    .valid(line_1776_valid)
  );
  assign line_1749_clock = clock;
  assign line_1749_reset = reset;
  assign line_1749_valid = _len_T ^ line_1749_valid_reg;
  assign line_1750_clock = clock;
  assign line_1750_reset = reset;
  assign line_1750_valid = _len_T ^ line_1750_valid_reg;
  assign line_1751_clock = clock;
  assign line_1751_reset = reset;
  assign line_1751_valid = _len_T ^ line_1751_valid_reg;
  assign line_1752_clock = clock;
  assign line_1752_reset = reset;
  assign line_1752_valid = ren ^ line_1752_valid_reg;
  assign line_1753_clock = clock;
  assign line_1753_reset = reset;
  assign line_1753_valid = _T_2 ^ line_1753_valid_reg;
  assign line_1754_clock = clock;
  assign line_1754_reset = reset;
  assign line_1754_valid = io_in_r_valid ^ line_1754_valid_reg;
  assign line_1755_clock = clock;
  assign line_1755_reset = reset;
  assign line_1755_valid = io_in_r_bits_last ^ line_1755_valid_reg;
  assign line_1756_clock = clock;
  assign line_1756_reset = reset;
  assign line_1756_valid = _len_T ^ line_1756_valid_reg;
  assign line_1757_clock = clock;
  assign line_1757_reset = reset;
  assign line_1757_valid = _T_5 ^ line_1757_valid_reg;
  assign line_1758_clock = clock;
  assign line_1758_reset = reset;
  assign line_1758_valid = _T_16 ^ line_1758_valid_reg;
  assign line_1759_clock = clock;
  assign line_1759_reset = reset;
  assign line_1759_valid = _T_17 ^ line_1759_valid_reg;
  assign line_1760_clock = clock;
  assign line_1760_reset = reset;
  assign line_1760_valid = _r_busy_T_2 ^ line_1760_valid_reg;
  assign line_1761_clock = clock;
  assign line_1761_reset = reset;
  assign line_1761_valid = _len_T ^ line_1761_valid_reg;
  assign line_1762_clock = clock;
  assign line_1762_reset = reset;
  assign line_1762_valid = io_in_r_valid ^ line_1762_valid_reg;
  assign line_1763_clock = clock;
  assign line_1763_reset = reset;
  assign line_1763_valid = _io_in_r_valid_T_2 ^ line_1763_valid_reg;
  assign line_1764_clock = clock;
  assign line_1764_reset = reset;
  assign line_1764_valid = _waddr_T ^ line_1764_valid_reg;
  assign line_1765_clock = clock;
  assign line_1765_reset = reset;
  assign line_1765_valid = _T_18 ^ line_1765_valid_reg;
  assign line_1766_clock = clock;
  assign line_1766_reset = reset;
  assign line_1766_valid = io_in_w_bits_last ^ line_1766_valid_reg;
  assign line_1767_clock = clock;
  assign line_1767_reset = reset;
  assign line_1767_valid = io_in_b_valid ^ line_1767_valid_reg;
  assign line_1768_clock = clock;
  assign line_1768_reset = reset;
  assign line_1768_valid = _waddr_T ^ line_1768_valid_reg;
  assign line_1769_clock = clock;
  assign line_1769_reset = reset;
  assign line_1769_valid = io_in_b_valid ^ line_1769_valid_reg;
  assign line_1770_clock = clock;
  assign line_1770_reset = reset;
  assign line_1770_valid = _io_in_b_valid_T_1 ^ line_1770_valid_reg;
  assign line_1771_clock = clock;
  assign line_1771_reset = reset;
  assign line_1771_valid = _waddr_T ^ line_1771_valid_reg;
  assign line_1772_clock = clock;
  assign line_1772_reset = reset;
  assign line_1772_valid = _waddr_T ^ line_1772_valid_reg;
  assign line_1773_clock = clock;
  assign line_1773_reset = reset;
  assign line_1773_valid = _len_T ^ line_1773_valid_reg;
  assign line_1774_clock = clock;
  assign line_1774_reset = reset;
  assign line_1774_valid = _len_T ^ line_1774_valid_reg;
  assign line_1775_clock = clock;
  assign line_1775_reset = reset;
  assign line_1775_valid = wen ^ line_1775_valid_reg;
  assign line_1776_clock = clock;
  assign line_1776_reset = reset;
  assign line_1776_valid = rdata_REG_1 ^ line_1776_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {rdata_hi_2,rdata_lo_2}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  assign io_in_r_bits_last = c_value == _GEN_28; // @[src/main/scala/device/AXI4Slave.scala 47:36]
  assign rdata_mem_clock = clock;
  assign rdata_mem_reset = reset;
  assign rdata_mem_read_valid = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  assign rdata_mem_read_index = {{28'd0}, rIdx}; // @[difftest/src/main/scala/common/Mem.scala 237:16]
  assign rdata_mem_write_valid = _T_18 & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 37:25]
  assign rdata_mem_write_index = {{35'd0}, wIdx};
  assign rdata_mem_write_data_0 = {rdata_hi,rdata_lo}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  assign rdata_mem_write_mask_0 = {fullMask_hi,fullMask_lo}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      c_value <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_in_r_valid) begin // @[src/main/scala/device/AXI4Slave.scala 52:28]
      if (io_in_r_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 54:33]
        c_value <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 54:43]
      end else begin
        c_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    readBeatCnt <= _GEN_60[7:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= 8'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= io_in_ar_bits_len; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_1749_valid_reg <= _len_T;
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h2; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_1750_valid_reg <= _len_T;
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= 39'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= wrapAddr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_1751_valid_reg <= _len_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _len_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    line_1752_valid_reg <= ren;
    line_1753_valid_reg <= _T_2;
    line_1754_valid_reg <= io_in_r_valid;
    line_1755_valid_reg <= io_in_r_bits_last;
    line_1756_valid_reg <= _len_T;
    line_1757_valid_reg <= _T_5;
    line_1758_valid_reg <= _T_16;
    line_1759_valid_reg <= _T_17;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_37;
    end
    line_1760_valid_reg <= _r_busy_T_2;
    line_1761_valid_reg <= _len_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_39;
    end
    line_1762_valid_reg <= io_in_r_valid;
    line_1763_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T_18) begin // @[src/main/scala/device/AXI4Slave.scala 82:28]
      if (io_in_w_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 84:33]
        writeBeatCnt <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 84:43]
      end else begin
        writeBeatCnt <= _value_T_7; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= 32'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_waddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= io_in_aw_bits_addr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_1764_valid_reg <= _waddr_T;
    line_1765_valid_reg <= _T_18;
    line_1766_valid_reg <= io_in_w_bits_last;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_44;
    end
    line_1767_valid_reg <= io_in_b_valid;
    line_1768_valid_reg <= _waddr_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_46;
    end
    line_1769_valid_reg <= io_in_b_valid;
    line_1770_valid_reg <= _io_in_b_valid_T_1;
    line_1771_valid_reg <= _waddr_T;
    line_1772_valid_reg <= _waddr_T;
    line_1773_valid_reg <= _len_T;
    line_1774_valid_reg <= _len_T;
    line_1775_valid_reg <= wen;
    rdata_REG <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    rdata_REG_1 <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    if (rdata_REG_1) begin // @[difftest/src/main/scala/common/Mem.scala 238:42]
      rdata_r_0 <= rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    line_1776_valid_reg <= rdata_REG_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_len_T & _T_5 & _T_16 & ~_T_14) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at AXI4Slave.scala:59 assert(axi4.ar.bits.len === 1.U || axi4.ar.bits.len === 3.U ||\n"
            ); // @[src/main/scala/device/AXI4Slave.scala 59:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_value = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  readBeatCnt = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  len_r = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  line_1749_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  burst_r = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  line_1750_valid_reg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  raddr_r = _RAND_6[38:0];
  _RAND_7 = {1{`RANDOM}};
  line_1751_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ren_REG = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1752_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1753_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1754_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1755_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1756_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1757_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1758_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1759_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_busy = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1760_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1761_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_1762_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_1763_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  writeBeatCnt = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  waddr_r = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  line_1764_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_1765_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_1766_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  w_busy = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_1767_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_1768_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_1769_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_1770_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_1771_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_1772_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_1773_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_1774_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_1775_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  rdata_REG = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  rdata_REG_1 = _RAND_40[0:0];
  _RAND_41 = {2{`RANDOM}};
  rdata_r_0 = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  line_1776_valid_reg = _RAND_42[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (ren) begin
      cover(1'h1);
    end
    //
    if (ren & _T_2) begin
      cover(1'h1);
    end
    //
    if (io_in_r_valid) begin
      cover(1'h1);
    end
    //
    if (io_in_r_valid & io_in_r_bits_last) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (_len_T & _T_5) begin
      cover(1'h1);
    end
    //
    if (_len_T & _T_5 & _T_16) begin
      cover(1'h1);
    end
    //
    if (_len_T & _T_5 & _T_16 & _T_17) begin
      cover(1'h1);
    end
    //
    if (_len_T & _T_5 & ~reset) begin
      assert(_T_14); // @[src/main/scala/device/AXI4Slave.scala 59:17]
    end
    //
    if (_r_busy_T_2) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (io_in_r_valid) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_waddr_T) begin
      cover(1'h1);
    end
    //
    if (_T_18) begin
      cover(1'h1);
    end
    //
    if (_T_18 & io_in_w_bits_last) begin
      cover(1'h1);
    end
    //
    if (io_in_b_valid) begin
      cover(1'h1);
    end
    //
    if (_waddr_T) begin
      cover(1'h1);
    end
    //
    if (io_in_b_valid) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T_1) begin
      cover(1'h1);
    end
    //
    if (_waddr_T) begin
      cover(1'h1);
    end
    //
    if (_waddr_T) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (_len_T) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (rdata_REG_1) begin
      cover(1'h1);
    end
  end
endmodule
module LatencyPipe(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [7:0]  io_in_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [7:0]  io_out_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [2:0]  io_out_bits_size // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_len = io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module LatencyPipe_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_out_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4Delayer(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
);
  wire  io_out_ar_pipe_clock; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_reset; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_clock; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_reset; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  LatencyPipe io_out_ar_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .clock(io_out_ar_pipe_clock),
    .reset(io_out_ar_pipe_reset),
    .io_in_valid(io_out_ar_pipe_io_in_valid),
    .io_in_bits_addr(io_out_ar_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_ar_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_ar_pipe_io_in_bits_size),
    .io_out_valid(io_out_ar_pipe_io_out_valid),
    .io_out_bits_addr(io_out_ar_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_ar_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_ar_pipe_io_out_bits_size)
  );
  LatencyPipe_1 io_out_aw_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .clock(io_out_aw_pipe_clock),
    .reset(io_out_aw_pipe_reset),
    .io_in_ready(io_out_aw_pipe_io_in_ready),
    .io_in_valid(io_out_aw_pipe_io_in_valid),
    .io_in_bits_addr(io_out_aw_pipe_io_in_bits_addr),
    .io_out_ready(io_out_aw_pipe_io_out_ready),
    .io_out_valid(io_out_aw_pipe_io_out_valid),
    .io_out_bits_addr(io_out_aw_pipe_io_out_bits_addr)
  );
  assign io_in_aw_ready = io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_w_ready = io_out_w_ready; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_in_b_valid = io_out_b_valid; // @[src/main/scala/bus/axi4/Delayer.scala 18:13]
  assign io_in_r_valid = io_out_r_valid; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_data = io_out_r_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_last = io_out_r_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_out_aw_valid = io_out_aw_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_aw_bits_addr = io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_w_valid = io_in_w_valid; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_data = io_in_w_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_strb = io_in_w_bits_strb; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_last = io_in_w_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_ar_valid = io_out_ar_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_addr = io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_len = io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_size = io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_pipe_clock = clock;
  assign io_out_ar_pipe_reset = reset;
  assign io_out_ar_pipe_io_in_valid = io_in_ar_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_addr = io_in_ar_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_len = io_in_ar_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_size = io_in_ar_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_clock = clock;
  assign io_out_aw_pipe_reset = reset;
  assign io_out_aw_pipe_io_in_valid = io_in_aw_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_addr = io_in_aw_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_out_ready = io_out_aw_ready; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBusCrossbar1toN_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_4_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_4_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_4_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_4_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_4_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h40600010; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h50000000 & io_in_req_bits_addr < 32'h50400000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40001000 & io_in_req_bits_addr < 32'h40001008; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_3 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h40001000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_4 = io_in_req_bits_addr >= 32'h40002000 & io_in_req_bits_addr < 32'h40003000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [4:0] _outSelVec_enc_T = outMatchVec_4 ? 5'h10 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_1 = outMatchVec_3 ? 5'h8 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_2 = outMatchVec_2 ? 5'h4 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_3 = outMatchVec_1 ? 5'h2 : _outSelVec_enc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] outSelVec_enc = outMatchVec_0 ? 5'h1 : _outSelVec_enc_T_3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_3 = outSelVec_enc[3]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_4 = outSelVec_enc[4]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  line_1777_clock;
  wire  line_1777_reset;
  wire  line_1777_valid;
  reg  line_1777_valid_reg;
  wire [4:0] _reqInvalidAddr_T = {outSelVec_4,outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
  wire  line_1778_clock;
  wire  line_1778_reset;
  wire  line_1778_valid;
  reg  line_1778_valid_reg;
  wire  _T_3 = ~(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
  wire  line_1779_clock;
  wire  line_1779_reset;
  wire  line_1779_valid;
  reg  line_1779_valid_reg;
  wire  _T_4 = 2'h0 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1780_clock;
  wire  line_1780_reset;
  wire  line_1780_valid;
  reg  line_1780_valid_reg;
  wire  line_1781_clock;
  wire  line_1781_reset;
  wire  line_1781_valid;
  reg  line_1781_valid_reg;
  wire  line_1782_clock;
  wire  line_1782_reset;
  wire  line_1782_valid;
  reg  line_1782_valid_reg;
  wire  line_1783_clock;
  wire  line_1783_reset;
  wire  line_1783_valid;
  reg  line_1783_valid_reg;
  wire  _T_6 = 2'h1 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1784_clock;
  wire  line_1784_reset;
  wire  line_1784_valid;
  reg  line_1784_valid_reg;
  wire  _T_7 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1785_clock;
  wire  line_1785_reset;
  wire  line_1785_valid;
  reg  line_1785_valid_reg;
  wire [1:0] _GEN_19 = _T_7 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  line_1786_clock;
  wire  line_1786_reset;
  wire  line_1786_valid;
  reg  line_1786_valid_reg;
  wire  _T_8 = 2'h2 == state; // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
  wire  line_1787_clock;
  wire  line_1787_reset;
  wire  line_1787_valid;
  reg  line_1787_valid_reg;
  wire  line_1788_clock;
  wire  line_1788_reset;
  wire  line_1788_valid;
  reg  line_1788_valid_reg;
  wire  _io_in_req_ready_T_8 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready | outSelVec_3 & io_out_3_req_ready | outSelVec_4 & io_out_4_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_8 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid | outSelRespVec_3 & io_out_3_resp_valid | outSelRespVec_4 &
    io_out_4_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = outSelRespVec_3 ? io_out_3_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_4 = outSelRespVec_4 ? io_out_4_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_6 = _io_in_resp_bits_T | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_7 = _io_in_resp_bits_T_6 | _io_in_resp_bits_T_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_9 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_10 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_11 = outSelRespVec_2 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_12 = outSelRespVec_3 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_13 = outSelRespVec_4 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_14 = _io_in_resp_bits_T_9 | _io_in_resp_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_15 = _io_in_resp_bits_T_14 | _io_in_resp_bits_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_16 = _io_in_resp_bits_T_15 | _io_in_resp_bits_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  GEN_w1_line #(.COVER_INDEX(1777)) line_1777 (
    .clock(line_1777_clock),
    .reset(line_1777_reset),
    .valid(line_1777_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1778)) line_1778 (
    .clock(line_1778_clock),
    .reset(line_1778_reset),
    .valid(line_1778_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1779)) line_1779 (
    .clock(line_1779_clock),
    .reset(line_1779_reset),
    .valid(line_1779_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1780)) line_1780 (
    .clock(line_1780_clock),
    .reset(line_1780_reset),
    .valid(line_1780_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1781)) line_1781 (
    .clock(line_1781_clock),
    .reset(line_1781_reset),
    .valid(line_1781_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1782)) line_1782 (
    .clock(line_1782_clock),
    .reset(line_1782_reset),
    .valid(line_1782_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1783)) line_1783 (
    .clock(line_1783_clock),
    .reset(line_1783_reset),
    .valid(line_1783_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1784)) line_1784 (
    .clock(line_1784_clock),
    .reset(line_1784_reset),
    .valid(line_1784_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1785)) line_1785 (
    .clock(line_1785_clock),
    .reset(line_1785_reset),
    .valid(line_1785_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1786)) line_1786 (
    .clock(line_1786_clock),
    .reset(line_1786_reset),
    .valid(line_1786_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1787)) line_1787 (
    .clock(line_1787_clock),
    .reset(line_1787_reset),
    .valid(line_1787_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1788)) line_1788 (
    .clock(line_1788_clock),
    .reset(line_1788_reset),
    .valid(line_1788_valid)
  );
  assign line_1777_clock = clock;
  assign line_1777_reset = reset;
  assign line_1777_valid = _outSelRespVec_T_2 ^ line_1777_valid_reg;
  assign line_1778_clock = clock;
  assign line_1778_reset = reset;
  assign line_1778_valid = _T_2 ^ line_1778_valid_reg;
  assign line_1779_clock = clock;
  assign line_1779_reset = reset;
  assign line_1779_valid = _T_3 ^ line_1779_valid_reg;
  assign line_1780_clock = clock;
  assign line_1780_reset = reset;
  assign line_1780_valid = _T_4 ^ line_1780_valid_reg;
  assign line_1781_clock = clock;
  assign line_1781_reset = reset;
  assign line_1781_valid = _outSelRespVec_T ^ line_1781_valid_reg;
  assign line_1782_clock = clock;
  assign line_1782_reset = reset;
  assign line_1782_valid = reqInvalidAddr ^ line_1782_valid_reg;
  assign line_1783_clock = clock;
  assign line_1783_reset = reset;
  assign line_1783_valid = _T_4 ^ line_1783_valid_reg;
  assign line_1784_clock = clock;
  assign line_1784_reset = reset;
  assign line_1784_valid = _T_6 ^ line_1784_valid_reg;
  assign line_1785_clock = clock;
  assign line_1785_reset = reset;
  assign line_1785_valid = _T_7 ^ line_1785_valid_reg;
  assign line_1786_clock = clock;
  assign line_1786_reset = reset;
  assign line_1786_valid = _T_6 ^ line_1786_valid_reg;
  assign line_1787_clock = clock;
  assign line_1787_reset = reset;
  assign line_1787_valid = _T_8 ^ line_1787_valid_reg;
  assign line_1788_clock = clock;
  assign line_1788_reset = reset;
  assign line_1788_valid = _T_7 ^ line_1788_valid_reg;
  assign io_in_req_ready = _io_in_req_ready_T_8 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_8 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_16 | _io_in_resp_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_7 | _io_in_resp_bits_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_3_req_valid = outSelVec_3 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_3_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_resp_ready = outSelRespVec_3 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_4_req_valid = outSelVec_4 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_4_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_resp_ready = outSelRespVec_4 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_19;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_19;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= outSelVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= outSelVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    line_1777_valid_reg <= _outSelRespVec_T_2;
    line_1778_valid_reg <= _T_2;
    line_1779_valid_reg <= _T_3;
    line_1780_valid_reg <= _T_4;
    line_1781_valid_reg <= _outSelRespVec_T;
    line_1782_valid_reg <= reqInvalidAddr;
    line_1783_valid_reg <= _T_4;
    line_1784_valid_reg <= _T_6;
    line_1785_valid_reg <= _T_7;
    line_1786_valid_reg <= _T_6;
    line_1787_valid_reg <= _T_8;
    line_1788_valid_reg <= _T_7;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  outSelRespVec_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  outSelRespVec_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1777_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1778_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1779_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1780_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1781_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1782_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1783_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1784_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1785_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1786_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1787_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1788_valid_reg = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_outSelRespVec_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
    //
    if (_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_4 & _outSelRespVec_T) begin
      cover(1'h1);
    end
    //
    if (_T_4 & reqInvalidAddr) begin
      cover(1'h1);
    end
    //
    if (~_T_4) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & _T_6 & _T_7) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6 & _T_8) begin
      cover(1'h1);
    end
    //
    if (~_T_4 & ~_T_6 & _T_8 & _T_7) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4UART(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_out_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_out_ch, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_in_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_extra_in_ch // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1789_clock;
  wire  line_1789_reset;
  wire  line_1789_valid;
  reg  line_1789_valid_reg;
  wire  _GEN_11 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1790_clock;
  wire  line_1790_reset;
  wire  line_1790_valid;
  reg  line_1790_valid_reg;
  wire  _GEN_12 = _r_busy_T | _GEN_11; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1791_clock;
  wire  line_1791_reset;
  wire  line_1791_valid;
  reg  line_1791_valid_reg;
  wire  _GEN_13 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1792_clock;
  wire  line_1792_reset;
  wire  line_1792_valid;
  reg  line_1792_valid_reg;
  wire  _GEN_14 = _io_in_r_valid_T_2 | _GEN_13; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1793_clock;
  wire  line_1793_reset;
  wire  line_1793_valid;
  reg  line_1793_valid_reg;
  wire  _GEN_15 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1794_clock;
  wire  line_1794_reset;
  wire  line_1794_valid;
  reg  line_1794_valid_reg;
  wire  _GEN_16 = _w_busy_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1795_clock;
  wire  line_1795_reset;
  wire  line_1795_valid;
  reg  line_1795_valid_reg;
  wire  _GEN_17 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1796_clock;
  wire  line_1796_reset;
  wire  line_1796_valid;
  reg  line_1796_valid_reg;
  wire  _GEN_18 = _io_in_b_valid_T | _GEN_17; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] txfifo; // @[src/main/scala/device/AXI4UART.scala 29:19]
  reg [31:0] stat; // @[src/main/scala/device/AXI4UART.scala 30:21]
  reg [31:0] ctrl; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire  _io_extra_out_valid_T_1 = io_in_aw_bits_addr[3:0] == 4'h4; // @[src/main/scala/device/AXI4UART.scala 33:41]
  wire [7:0] _T_5 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4UART.scala 45:79]
  wire [7:0] _T_14 = _T_5[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_15 = _T_5[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_16 = _T_5[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_17 = _T_5[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_18 = _T_5[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_19 = _T_5[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_20 = _T_5[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_21 = _T_5[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_22 = {_T_21,_T_20,_T_19,_T_18,_T_17,_T_16,_T_15,_T_14}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 4'hc == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [7:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T ? io_extra_in_ch : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_1 ? txfifo : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_2 ? stat : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_3 ? ctrl : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_22 = {{24'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_8 = _GEN_22 | _io_in_r_bits_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_8 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_9 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_25 = _io_in_b_valid_T & _io_extra_out_valid_T_1; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1797_clock;
  wire  line_1797_reset;
  wire  line_1797_valid;
  reg  line_1797_valid_reg;
  wire [31:0] _txfifo_T = io_in_w_bits_data[31:0] & _T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _txfifo_T_1 = ~_T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _txfifo_T_2 = txfifo & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _txfifo_T_3 = _txfifo_T | _txfifo_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_27 = _io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1798_clock;
  wire  line_1798_reset;
  wire  line_1798_valid;
  reg  line_1798_valid_reg;
  wire [31:0] _stat_T_2 = stat & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _stat_T_3 = _txfifo_T | _stat_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_29 = _io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'hc; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1799_clock;
  wire  line_1799_reset;
  wire  line_1799_valid;
  reg  line_1799_valid_reg;
  wire [31:0] _ctrl_T_2 = ctrl & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _ctrl_T_3 = _txfifo_T | _ctrl_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  GEN_w1_line #(.COVER_INDEX(1789)) line_1789 (
    .clock(line_1789_clock),
    .reset(line_1789_reset),
    .valid(line_1789_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1790)) line_1790 (
    .clock(line_1790_clock),
    .reset(line_1790_reset),
    .valid(line_1790_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1791)) line_1791 (
    .clock(line_1791_clock),
    .reset(line_1791_reset),
    .valid(line_1791_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1792)) line_1792 (
    .clock(line_1792_clock),
    .reset(line_1792_reset),
    .valid(line_1792_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1793)) line_1793 (
    .clock(line_1793_clock),
    .reset(line_1793_reset),
    .valid(line_1793_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1794)) line_1794 (
    .clock(line_1794_clock),
    .reset(line_1794_reset),
    .valid(line_1794_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1795)) line_1795 (
    .clock(line_1795_clock),
    .reset(line_1795_reset),
    .valid(line_1795_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1796)) line_1796 (
    .clock(line_1796_clock),
    .reset(line_1796_reset),
    .valid(line_1796_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1797)) line_1797 (
    .clock(line_1797_clock),
    .reset(line_1797_reset),
    .valid(line_1797_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1798)) line_1798 (
    .clock(line_1798_clock),
    .reset(line_1798_reset),
    .valid(line_1798_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1799)) line_1799 (
    .clock(line_1799_clock),
    .reset(line_1799_reset),
    .valid(line_1799_valid)
  );
  assign line_1789_clock = clock;
  assign line_1789_reset = reset;
  assign line_1789_valid = _r_busy_T_1 ^ line_1789_valid_reg;
  assign line_1790_clock = clock;
  assign line_1790_reset = reset;
  assign line_1790_valid = _r_busy_T ^ line_1790_valid_reg;
  assign line_1791_clock = clock;
  assign line_1791_reset = reset;
  assign line_1791_valid = _r_busy_T_1 ^ line_1791_valid_reg;
  assign line_1792_clock = clock;
  assign line_1792_reset = reset;
  assign line_1792_valid = _io_in_r_valid_T_2 ^ line_1792_valid_reg;
  assign line_1793_clock = clock;
  assign line_1793_reset = reset;
  assign line_1793_valid = _w_busy_T_1 ^ line_1793_valid_reg;
  assign line_1794_clock = clock;
  assign line_1794_reset = reset;
  assign line_1794_valid = _w_busy_T ^ line_1794_valid_reg;
  assign line_1795_clock = clock;
  assign line_1795_reset = reset;
  assign line_1795_valid = _w_busy_T_1 ^ line_1795_valid_reg;
  assign line_1796_clock = clock;
  assign line_1796_reset = reset;
  assign line_1796_valid = _io_in_b_valid_T ^ line_1796_valid_reg;
  assign line_1797_clock = clock;
  assign line_1797_reset = reset;
  assign line_1797_valid = _T_25 ^ line_1797_valid_reg;
  assign line_1798_clock = clock;
  assign line_1798_reset = reset;
  assign line_1798_valid = _T_27 ^ line_1798_valid_reg;
  assign line_1799_clock = clock;
  assign line_1799_reset = reset;
  assign line_1799_valid = _T_29 ^ line_1799_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_10}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_out_valid = io_in_aw_bits_addr[3:0] == 4'h4 & _io_in_b_valid_T; // @[src/main/scala/device/AXI4UART.scala 33:49]
  assign io_extra_out_ch = io_in_w_bits_data[7:0]; // @[src/main/scala/device/AXI4UART.scala 34:40]
  assign io_extra_in_valid = io_in_ar_bits_addr[3:0] == 4'h0 & _r_busy_T_1; // @[src/main/scala/device/AXI4UART.scala 35:48]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_12;
    end
    line_1789_valid_reg <= _r_busy_T_1;
    line_1790_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_14;
    end
    line_1791_valid_reg <= _r_busy_T_1;
    line_1792_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_16;
    end
    line_1793_valid_reg <= _w_busy_T_1;
    line_1794_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_18;
    end
    line_1795_valid_reg <= _w_busy_T_1;
    line_1796_valid_reg <= _io_in_b_valid_T;
    if (_io_in_b_valid_T & _io_extra_out_valid_T_1) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      txfifo <= _txfifo_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 30:21]
      stat <= 32'h1; // @[src/main/scala/device/AXI4UART.scala 30:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      stat <= _stat_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 31:21]
      ctrl <= 32'h0; // @[src/main/scala/device/AXI4UART.scala 31:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'hc) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      ctrl <= _ctrl_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    line_1797_valid_reg <= _T_25;
    line_1798_valid_reg <= _T_27;
    line_1799_valid_reg <= _T_29;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1789_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1790_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1791_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1792_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1793_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1794_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1795_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1796_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  txfifo = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stat = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  ctrl = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  line_1797_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1798_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1799_valid_reg = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (_T_25) begin
      cover(1'h1);
    end
    //
    if (_T_27) begin
      cover(1'h1);
    end
    //
    if (_T_29) begin
      cover(1'h1);
    end
  end
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_sync // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1800_clock;
  wire  line_1800_reset;
  wire  line_1800_valid;
  reg  line_1800_valid_reg;
  wire  _GEN_8 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1801_clock;
  wire  line_1801_reset;
  wire  line_1801_valid;
  reg  line_1801_valid_reg;
  wire  _GEN_9 = _r_busy_T | _GEN_8; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1802_clock;
  wire  line_1802_reset;
  wire  line_1802_valid;
  reg  line_1802_valid_reg;
  wire  _GEN_10 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1803_clock;
  wire  line_1803_reset;
  wire  line_1803_valid;
  reg  line_1803_valid_reg;
  wire  _GEN_11 = _io_in_r_valid_T_2 | _GEN_10; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1804_clock;
  wire  line_1804_reset;
  wire  line_1804_valid;
  reg  line_1804_valid_reg;
  wire  _GEN_12 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1805_clock;
  wire  line_1805_reset;
  wire  line_1805_valid;
  reg  line_1805_valid_reg;
  wire  _GEN_13 = _w_busy_T | _GEN_12; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1806_clock;
  wire  line_1806_reset;
  wire  line_1806_valid;
  reg  line_1806_valid_reg;
  wire  _GEN_14 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1807_clock;
  wire  line_1807_reset;
  wire  line_1807_valid;
  reg  line_1807_valid_reg;
  wire  _GEN_15 = _io_in_b_valid_T | _GEN_14; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _io_in_r_bits_data_T_2 = _io_in_r_bits_data_T ? 32'h190012c : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_r_bits_data_T_3 = _io_in_r_bits_data_T_1 & _w_busy_T; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_16 = {{31'd0}, _io_in_r_bits_data_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T_2 | _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  GEN_w1_line #(.COVER_INDEX(1800)) line_1800 (
    .clock(line_1800_clock),
    .reset(line_1800_reset),
    .valid(line_1800_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1801)) line_1801 (
    .clock(line_1801_clock),
    .reset(line_1801_reset),
    .valid(line_1801_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1802)) line_1802 (
    .clock(line_1802_clock),
    .reset(line_1802_reset),
    .valid(line_1802_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1803)) line_1803 (
    .clock(line_1803_clock),
    .reset(line_1803_reset),
    .valid(line_1803_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1804)) line_1804 (
    .clock(line_1804_clock),
    .reset(line_1804_reset),
    .valid(line_1804_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1805)) line_1805 (
    .clock(line_1805_clock),
    .reset(line_1805_reset),
    .valid(line_1805_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1806)) line_1806 (
    .clock(line_1806_clock),
    .reset(line_1806_reset),
    .valid(line_1806_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1807)) line_1807 (
    .clock(line_1807_clock),
    .reset(line_1807_reset),
    .valid(line_1807_valid)
  );
  assign line_1800_clock = clock;
  assign line_1800_reset = reset;
  assign line_1800_valid = _r_busy_T_1 ^ line_1800_valid_reg;
  assign line_1801_clock = clock;
  assign line_1801_reset = reset;
  assign line_1801_valid = _r_busy_T ^ line_1801_valid_reg;
  assign line_1802_clock = clock;
  assign line_1802_reset = reset;
  assign line_1802_valid = _r_busy_T_1 ^ line_1802_valid_reg;
  assign line_1803_clock = clock;
  assign line_1803_reset = reset;
  assign line_1803_valid = _io_in_r_valid_T_2 ^ line_1803_valid_reg;
  assign line_1804_clock = clock;
  assign line_1804_reset = reset;
  assign line_1804_valid = _w_busy_T_1 ^ line_1804_valid_reg;
  assign line_1805_clock = clock;
  assign line_1805_reset = reset;
  assign line_1805_valid = _w_busy_T ^ line_1805_valid_reg;
  assign line_1806_clock = clock;
  assign line_1806_reset = reset;
  assign line_1806_valid = _w_busy_T_1 ^ line_1806_valid_reg;
  assign line_1807_clock = clock;
  assign line_1807_reset = reset;
  assign line_1807_valid = _io_in_b_valid_T ^ line_1807_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_sync = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_9;
    end
    line_1800_valid_reg <= _r_busy_T_1;
    line_1801_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_11;
    end
    line_1802_valid_reg <= _r_busy_T_1;
    line_1803_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_13;
    end
    line_1804_valid_reg <= _w_busy_T_1;
    line_1805_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_15;
    end
    line_1806_valid_reg <= _w_busy_T_1;
    line_1807_valid_reg <= _io_in_b_valid_T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1800_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1801_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1802_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1803_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1804_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1805_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1806_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1807_valid_reg = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4RAM_1(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] rdata_mem_0 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_1 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_2 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_3 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_4 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_5 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_6 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_7 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1808_clock;
  wire  line_1808_reset;
  wire  line_1808_valid;
  reg  line_1808_valid_reg;
  wire  _GEN_18 = io_in_r_valid ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1809_clock;
  wire  line_1809_reset;
  wire  line_1809_valid;
  reg  line_1809_valid_reg;
  wire  _GEN_19 = _r_busy_T | _GEN_18; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1810_clock;
  wire  line_1810_reset;
  wire  line_1810_valid;
  reg  line_1810_valid_reg;
  wire  _GEN_20 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1811_clock;
  wire  line_1811_reset;
  wire  line_1811_valid;
  reg  line_1811_valid_reg;
  wire  _GEN_21 = _io_in_r_valid_T_2 | _GEN_20; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1812_clock;
  wire  line_1812_reset;
  wire  line_1812_valid;
  reg  line_1812_valid_reg;
  wire  _GEN_22 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1813_clock;
  wire  line_1813_reset;
  wire  line_1813_valid;
  reg  line_1813_valid_reg;
  wire  _GEN_23 = _w_busy_T | _GEN_22; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1814_clock;
  wire  line_1814_reset;
  wire  line_1814_valid;
  reg  line_1814_valid_reg;
  wire  _GEN_24 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1815_clock;
  wire  line_1815_reset;
  wire  line_1815_valid;
  reg  line_1815_valid_reg;
  wire  _GEN_25 = _io_in_b_valid_T | _GEN_24; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = io_in_aw_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _wIdx_T_2 = {{1'd0}, _wIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [31:0] _rIdx_T = io_in_ar_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _rIdx_T_2 = {{1'd0}, _rIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [28:0] rIdx = _rIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'hea60; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire  wen = _io_in_b_valid_T & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 37:25]
  wire  line_1816_clock;
  wire  line_1816_reset;
  wire  line_1816_valid;
  reg  line_1816_valid_reg;
  wire  line_1817_clock;
  wire  line_1817_reset;
  wire  line_1817_valid;
  reg  line_1817_valid_reg;
  wire  line_1818_clock;
  wire  line_1818_reset;
  wire  line_1818_valid;
  reg  line_1818_valid_reg;
  wire  line_1819_clock;
  wire  line_1819_reset;
  wire  line_1819_valid;
  reg  line_1819_valid_reg;
  wire  line_1820_clock;
  wire  line_1820_reset;
  wire  line_1820_valid;
  reg  line_1820_valid_reg;
  wire  line_1821_clock;
  wire  line_1821_reset;
  wire  line_1821_valid;
  reg  line_1821_valid_reg;
  wire  line_1822_clock;
  wire  line_1822_reset;
  wire  line_1822_valid;
  reg  line_1822_valid_reg;
  wire  line_1823_clock;
  wire  line_1823_reset;
  wire  line_1823_valid;
  reg  line_1823_valid_reg;
  wire  line_1824_clock;
  wire  line_1824_reset;
  wire  line_1824_valid;
  reg  line_1824_valid_reg;
  wire [63:0] _rdata_T_12 = {rdata_mem_7_rdata_MPORT_1_data,rdata_mem_6_rdata_MPORT_1_data,
    rdata_mem_5_rdata_MPORT_1_data,rdata_mem_4_rdata_MPORT_1_data,rdata_mem_3_rdata_MPORT_1_data,
    rdata_mem_2_rdata_MPORT_1_data,rdata_mem_1_rdata_MPORT_1_data,rdata_mem_0_rdata_MPORT_1_data}; // @[src/main/scala/device/AXI4RAM.scala 55:18]
  reg [63:0] rdata; // @[src/main/scala/device/AXI4RAM.scala 55:14]
  wire  line_1825_clock;
  wire  line_1825_reset;
  wire  line_1825_valid;
  reg  line_1825_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1808)) line_1808 (
    .clock(line_1808_clock),
    .reset(line_1808_reset),
    .valid(line_1808_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1809)) line_1809 (
    .clock(line_1809_clock),
    .reset(line_1809_reset),
    .valid(line_1809_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1810)) line_1810 (
    .clock(line_1810_clock),
    .reset(line_1810_reset),
    .valid(line_1810_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1811)) line_1811 (
    .clock(line_1811_clock),
    .reset(line_1811_reset),
    .valid(line_1811_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1812)) line_1812 (
    .clock(line_1812_clock),
    .reset(line_1812_reset),
    .valid(line_1812_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1813)) line_1813 (
    .clock(line_1813_clock),
    .reset(line_1813_reset),
    .valid(line_1813_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1814)) line_1814 (
    .clock(line_1814_clock),
    .reset(line_1814_reset),
    .valid(line_1814_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1815)) line_1815 (
    .clock(line_1815_clock),
    .reset(line_1815_reset),
    .valid(line_1815_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1816)) line_1816 (
    .clock(line_1816_clock),
    .reset(line_1816_reset),
    .valid(line_1816_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1817)) line_1817 (
    .clock(line_1817_clock),
    .reset(line_1817_reset),
    .valid(line_1817_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1818)) line_1818 (
    .clock(line_1818_clock),
    .reset(line_1818_reset),
    .valid(line_1818_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1819)) line_1819 (
    .clock(line_1819_clock),
    .reset(line_1819_reset),
    .valid(line_1819_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1820)) line_1820 (
    .clock(line_1820_clock),
    .reset(line_1820_reset),
    .valid(line_1820_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1821)) line_1821 (
    .clock(line_1821_clock),
    .reset(line_1821_reset),
    .valid(line_1821_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1822)) line_1822 (
    .clock(line_1822_clock),
    .reset(line_1822_reset),
    .valid(line_1822_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1823)) line_1823 (
    .clock(line_1823_clock),
    .reset(line_1823_reset),
    .valid(line_1823_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1824)) line_1824 (
    .clock(line_1824_clock),
    .reset(line_1824_reset),
    .valid(line_1824_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1825)) line_1825 (
    .clock(line_1825_clock),
    .reset(line_1825_reset),
    .valid(line_1825_valid)
  );
  assign rdata_mem_0_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_0_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_1[7:0] :
    rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_data = io_in_w_bits_data[7:0];
  assign rdata_mem_0_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_0_rdata_MPORT_mask = io_in_w_bits_strb[0];
  assign rdata_mem_0_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_1_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_1_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_3[7:0] :
    rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_data = io_in_w_bits_data[15:8];
  assign rdata_mem_1_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_1_rdata_MPORT_mask = io_in_w_bits_strb[1];
  assign rdata_mem_1_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_2_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_2_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_5[7:0] :
    rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_data = io_in_w_bits_data[23:16];
  assign rdata_mem_2_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_2_rdata_MPORT_mask = io_in_w_bits_strb[2];
  assign rdata_mem_2_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_3_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_3_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_7[7:0] :
    rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_data = io_in_w_bits_data[31:24];
  assign rdata_mem_3_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_3_rdata_MPORT_mask = io_in_w_bits_strb[3];
  assign rdata_mem_3_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_4_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_4_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_9[7:0] :
    rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_data = io_in_w_bits_data[39:32];
  assign rdata_mem_4_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_4_rdata_MPORT_mask = io_in_w_bits_strb[4];
  assign rdata_mem_4_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_5_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_5_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_11[7:0] :
    rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_data = io_in_w_bits_data[47:40];
  assign rdata_mem_5_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_5_rdata_MPORT_mask = io_in_w_bits_strb[5];
  assign rdata_mem_5_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_6_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_6_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_13[7:0] :
    rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_data = io_in_w_bits_data[55:48];
  assign rdata_mem_6_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_6_rdata_MPORT_mask = io_in_w_bits_strb[6];
  assign rdata_mem_6_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_7_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_7_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_15[7:0] :
    rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_data = io_in_w_bits_data[63:56];
  assign rdata_mem_7_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_7_rdata_MPORT_mask = io_in_w_bits_strb[7];
  assign rdata_mem_7_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign line_1808_clock = clock;
  assign line_1808_reset = reset;
  assign line_1808_valid = io_in_r_valid ^ line_1808_valid_reg;
  assign line_1809_clock = clock;
  assign line_1809_reset = reset;
  assign line_1809_valid = _r_busy_T ^ line_1809_valid_reg;
  assign line_1810_clock = clock;
  assign line_1810_reset = reset;
  assign line_1810_valid = io_in_r_valid ^ line_1810_valid_reg;
  assign line_1811_clock = clock;
  assign line_1811_reset = reset;
  assign line_1811_valid = _io_in_r_valid_T_2 ^ line_1811_valid_reg;
  assign line_1812_clock = clock;
  assign line_1812_reset = reset;
  assign line_1812_valid = _w_busy_T_1 ^ line_1812_valid_reg;
  assign line_1813_clock = clock;
  assign line_1813_reset = reset;
  assign line_1813_valid = _w_busy_T ^ line_1813_valid_reg;
  assign line_1814_clock = clock;
  assign line_1814_reset = reset;
  assign line_1814_valid = _w_busy_T_1 ^ line_1814_valid_reg;
  assign line_1815_clock = clock;
  assign line_1815_reset = reset;
  assign line_1815_valid = _io_in_b_valid_T ^ line_1815_valid_reg;
  assign line_1816_clock = clock;
  assign line_1816_reset = reset;
  assign line_1816_valid = wen ^ line_1816_valid_reg;
  assign line_1817_clock = clock;
  assign line_1817_reset = reset;
  assign line_1817_valid = io_in_w_bits_strb[0] ^ line_1817_valid_reg;
  assign line_1818_clock = clock;
  assign line_1818_reset = reset;
  assign line_1818_valid = io_in_w_bits_strb[1] ^ line_1818_valid_reg;
  assign line_1819_clock = clock;
  assign line_1819_reset = reset;
  assign line_1819_valid = io_in_w_bits_strb[2] ^ line_1819_valid_reg;
  assign line_1820_clock = clock;
  assign line_1820_reset = reset;
  assign line_1820_valid = io_in_w_bits_strb[3] ^ line_1820_valid_reg;
  assign line_1821_clock = clock;
  assign line_1821_reset = reset;
  assign line_1821_valid = io_in_w_bits_strb[4] ^ line_1821_valid_reg;
  assign line_1822_clock = clock;
  assign line_1822_reset = reset;
  assign line_1822_valid = io_in_w_bits_strb[5] ^ line_1822_valid_reg;
  assign line_1823_clock = clock;
  assign line_1823_reset = reset;
  assign line_1823_valid = io_in_w_bits_strb[6] ^ line_1823_valid_reg;
  assign line_1824_clock = clock;
  assign line_1824_reset = reset;
  assign line_1824_valid = io_in_w_bits_strb[7] ^ line_1824_valid_reg;
  assign line_1825_clock = clock;
  assign line_1825_reset = reset;
  assign line_1825_valid = ren_REG ^ line_1825_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = rdata; // @[src/main/scala/device/AXI4RAM.scala 58:18]
  always @(posedge clock) begin
    if (rdata_mem_0_rdata_MPORT_en & rdata_mem_0_rdata_MPORT_mask) begin
      rdata_mem_0[rdata_mem_0_rdata_MPORT_addr] <= rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_1_rdata_MPORT_en & rdata_mem_1_rdata_MPORT_mask) begin
      rdata_mem_1[rdata_mem_1_rdata_MPORT_addr] <= rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_2_rdata_MPORT_en & rdata_mem_2_rdata_MPORT_mask) begin
      rdata_mem_2[rdata_mem_2_rdata_MPORT_addr] <= rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_3_rdata_MPORT_en & rdata_mem_3_rdata_MPORT_mask) begin
      rdata_mem_3[rdata_mem_3_rdata_MPORT_addr] <= rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_4_rdata_MPORT_en & rdata_mem_4_rdata_MPORT_mask) begin
      rdata_mem_4[rdata_mem_4_rdata_MPORT_addr] <= rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_5_rdata_MPORT_en & rdata_mem_5_rdata_MPORT_mask) begin
      rdata_mem_5[rdata_mem_5_rdata_MPORT_addr] <= rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_6_rdata_MPORT_en & rdata_mem_6_rdata_MPORT_mask) begin
      rdata_mem_6[rdata_mem_6_rdata_MPORT_addr] <= rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_7_rdata_MPORT_en & rdata_mem_7_rdata_MPORT_mask) begin
      rdata_mem_7[rdata_mem_7_rdata_MPORT_addr] <= rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_19;
    end
    line_1808_valid_reg <= io_in_r_valid;
    line_1809_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_21;
    end
    line_1810_valid_reg <= io_in_r_valid;
    line_1811_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_23;
    end
    line_1812_valid_reg <= _w_busy_T_1;
    line_1813_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_25;
    end
    line_1814_valid_reg <= _w_busy_T_1;
    line_1815_valid_reg <= _io_in_b_valid_T;
    line_1816_valid_reg <= wen;
    line_1817_valid_reg <= io_in_w_bits_strb[0];
    line_1818_valid_reg <= io_in_w_bits_strb[1];
    line_1819_valid_reg <= io_in_w_bits_strb[2];
    line_1820_valid_reg <= io_in_w_bits_strb[3];
    line_1821_valid_reg <= io_in_w_bits_strb[4];
    line_1822_valid_reg <= io_in_w_bits_strb[5];
    line_1823_valid_reg <= io_in_w_bits_strb[6];
    line_1824_valid_reg <= io_in_w_bits_strb[7];
    if (ren_REG) begin // @[src/main/scala/device/AXI4RAM.scala 55:14]
      rdata <= _rdata_T_12; // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    line_1825_valid_reg <= ren_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1808_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1809_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ren_REG = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_1810_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_1811_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  w_busy = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_1812_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_1813_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_1814_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_1815_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_1816_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_1817_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_1818_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_1819_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_1820_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_1821_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_1822_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_1823_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_1824_valid_reg = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  rdata = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  line_1825_valid_reg = _RAND_39[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (io_in_r_valid) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (io_in_r_valid) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (wen) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[0]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[1]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[2]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[3]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[4]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[5]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[6]) begin
      cover(1'h1);
    end
    //
    if (wen & io_in_w_bits_strb[7]) begin
      cover(1'h1);
    end
    //
    if (ren_REG) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_fb_aw_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [63:0] io_in_fb_w_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [7:0]  io_in_fb_w_bits_strb, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_ctrl_ar_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output [63:0] io_in_ctrl_r_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_vga_valid // @[src/main/scala/device/AXI4VGA.scala 117:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  fb_clock; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_reset; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fbHelper_clk; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_valid; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire [31:0] fbHelper_pixel; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_sync; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  _io_in_fb_r_valid_T = io_in_fb_ar_ready & io_in_fb_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _io_in_fb_r_valid_T_1 = io_in_fb_r_ready & io_in_fb_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1826_clock;
  wire  line_1826_reset;
  wire  line_1826_valid;
  reg  line_1826_valid_reg;
  wire  _GEN_11 = _io_in_fb_r_valid_T_1 ? 1'h0 : io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1827_clock;
  wire  line_1827_reset;
  wire  line_1827_valid;
  reg  line_1827_valid_reg;
  wire  _GEN_12 = _io_in_fb_r_valid_T | _GEN_11; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [10:0] hCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = hCounter == 11'h41f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [10:0] _wrap_value_T_1 = hCounter + 11'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1828_clock;
  wire  line_1828_reset;
  wire  line_1828_valid;
  reg  line_1828_valid_reg;
  reg [9:0] vCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_1829_clock;
  wire  line_1829_reset;
  wire  line_1829_valid;
  reg  line_1829_valid_reg;
  wire  wrap_wrap_1 = vCounter == 10'h273; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [9:0] _wrap_value_T_3 = vCounter + 10'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1830_clock;
  wire  line_1830_reset;
  wire  line_1830_valid;
  reg  line_1830_valid_reg;
  wire  hInRange = hCounter >= 11'ha8 & hCounter < 11'h3c8; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  vInRange = vCounter >= 10'h5 & vCounter < 10'h25d; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[src/main/scala/device/AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 152:31]
  wire  _nextPixel_T_2 = hCounter >= 11'ha7 & hCounter < 11'h3c7; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  nextPixel = _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
  wire  _fbPixelAddrV0_T_1 = nextPixel & ~vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_1831_clock;
  wire  line_1831_reset;
  wire  line_1831_valid;
  reg  line_1831_valid_reg;
  wire  fbPixelAddrV0_wrap_wrap = fbPixelAddrV0 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV0_wrap_value_T_1 = fbPixelAddrV0 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1832_clock;
  wire  line_1832_reset;
  wire  line_1832_valid;
  reg  line_1832_valid_reg;
  wire  _fbPixelAddrV1_T = nextPixel & vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  line_1833_clock;
  wire  line_1833_reset;
  wire  line_1833_valid;
  reg  line_1833_valid_reg;
  wire  fbPixelAddrV1_wrap_wrap = fbPixelAddrV1 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV1_wrap_value_T_1 = fbPixelAddrV1 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_1834_clock;
  wire  line_1834_reset;
  wire  line_1834_valid;
  reg  line_1834_valid_reg;
  wire [16:0] _fb_io_in_ar_bits_addr_T = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[src/main/scala/device/AXI4VGA.scala 161:35]
  wire [18:0] _fb_io_in_ar_bits_addr_T_1 = {_fb_io_in_ar_bits_addr_T,2'h0}; // @[src/main/scala/device/AXI4VGA.scala 161:31]
  reg  fb_io_in_ar_valid_REG; // @[src/main/scala/device/AXI4VGA.scala 162:31]
  wire  _data_T = fb_io_in_r_ready & fb_io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] data_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  line_1835_clock;
  wire  line_1835_reset;
  wire  line_1835_valid;
  reg  line_1835_valid_reg;
  wire [63:0] _GEN_25 = _data_T ? fb_io_in_r_bits_data : data_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  VGACtrl ctrl ( // @[src/main/scala/device/AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_aw_ready(ctrl_io_in_aw_ready),
    .io_in_aw_valid(ctrl_io_in_aw_valid),
    .io_in_w_ready(ctrl_io_in_w_ready),
    .io_in_w_valid(ctrl_io_in_w_valid),
    .io_in_b_ready(ctrl_io_in_b_ready),
    .io_in_b_valid(ctrl_io_in_b_valid),
    .io_in_ar_ready(ctrl_io_in_ar_ready),
    .io_in_ar_valid(ctrl_io_in_ar_valid),
    .io_in_ar_bits_addr(ctrl_io_in_ar_bits_addr),
    .io_in_r_ready(ctrl_io_in_r_ready),
    .io_in_r_valid(ctrl_io_in_r_valid),
    .io_in_r_bits_data(ctrl_io_in_r_bits_data),
    .io_extra_sync(ctrl_io_extra_sync)
  );
  AXI4RAM_1 fb ( // @[src/main/scala/device/AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_aw_ready(fb_io_in_aw_ready),
    .io_in_aw_valid(fb_io_in_aw_valid),
    .io_in_aw_bits_addr(fb_io_in_aw_bits_addr),
    .io_in_w_ready(fb_io_in_w_ready),
    .io_in_w_valid(fb_io_in_w_valid),
    .io_in_w_bits_data(fb_io_in_w_bits_data),
    .io_in_w_bits_strb(fb_io_in_w_bits_strb),
    .io_in_b_ready(fb_io_in_b_ready),
    .io_in_b_valid(fb_io_in_b_valid),
    .io_in_ar_ready(fb_io_in_ar_ready),
    .io_in_ar_valid(fb_io_in_ar_valid),
    .io_in_ar_bits_addr(fb_io_in_ar_bits_addr),
    .io_in_r_ready(fb_io_in_r_ready),
    .io_in_r_valid(fb_io_in_r_valid),
    .io_in_r_bits_data(fb_io_in_r_bits_data)
  );
  FBHelper fbHelper ( // @[src/main/scala/device/AXI4VGA.scala 171:26]
    .clk(fbHelper_clk),
    .valid(fbHelper_valid),
    .pixel(fbHelper_pixel),
    .sync(fbHelper_sync)
  );
  GEN_w1_line #(.COVER_INDEX(1826)) line_1826 (
    .clock(line_1826_clock),
    .reset(line_1826_reset),
    .valid(line_1826_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1827)) line_1827 (
    .clock(line_1827_clock),
    .reset(line_1827_reset),
    .valid(line_1827_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1828)) line_1828 (
    .clock(line_1828_clock),
    .reset(line_1828_reset),
    .valid(line_1828_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1829)) line_1829 (
    .clock(line_1829_clock),
    .reset(line_1829_reset),
    .valid(line_1829_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1830)) line_1830 (
    .clock(line_1830_clock),
    .reset(line_1830_reset),
    .valid(line_1830_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1831)) line_1831 (
    .clock(line_1831_clock),
    .reset(line_1831_reset),
    .valid(line_1831_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1832)) line_1832 (
    .clock(line_1832_clock),
    .reset(line_1832_reset),
    .valid(line_1832_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1833)) line_1833 (
    .clock(line_1833_clock),
    .reset(line_1833_reset),
    .valid(line_1833_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1834)) line_1834 (
    .clock(line_1834_clock),
    .reset(line_1834_reset),
    .valid(line_1834_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1835)) line_1835 (
    .clock(line_1835_clock),
    .reset(line_1835_reset),
    .valid(line_1835_valid)
  );
  assign line_1826_clock = clock;
  assign line_1826_reset = reset;
  assign line_1826_valid = _io_in_fb_r_valid_T_1 ^ line_1826_valid_reg;
  assign line_1827_clock = clock;
  assign line_1827_reset = reset;
  assign line_1827_valid = _io_in_fb_r_valid_T ^ line_1827_valid_reg;
  assign line_1828_clock = clock;
  assign line_1828_reset = reset;
  assign line_1828_valid = wrap_wrap ^ line_1828_valid_reg;
  assign line_1829_clock = clock;
  assign line_1829_reset = reset;
  assign line_1829_valid = wrap_wrap ^ line_1829_valid_reg;
  assign line_1830_clock = clock;
  assign line_1830_reset = reset;
  assign line_1830_valid = wrap_wrap_1 ^ line_1830_valid_reg;
  assign line_1831_clock = clock;
  assign line_1831_reset = reset;
  assign line_1831_valid = _fbPixelAddrV0_T_1 ^ line_1831_valid_reg;
  assign line_1832_clock = clock;
  assign line_1832_reset = reset;
  assign line_1832_valid = fbPixelAddrV0_wrap_wrap ^ line_1832_valid_reg;
  assign line_1833_clock = clock;
  assign line_1833_reset = reset;
  assign line_1833_valid = _fbPixelAddrV1_T ^ line_1833_valid_reg;
  assign line_1834_clock = clock;
  assign line_1834_reset = reset;
  assign line_1834_valid = fbPixelAddrV1_wrap_wrap ^ line_1834_valid_reg;
  assign line_1835_clock = clock;
  assign line_1835_reset = reset;
  assign line_1835_valid = _data_T ^ line_1835_valid_reg;
  assign io_in_fb_aw_ready = fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign io_in_fb_w_ready = fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign io_in_fb_b_valid = fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign io_in_fb_ar_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 133:21]
  assign io_in_fb_r_valid = io_in_fb_r_valid_r; // @[src/main/scala/device/AXI4VGA.scala 136:20]
  assign io_in_ctrl_aw_ready = ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_w_ready = ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_b_valid = ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_ar_ready = ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_valid = ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_bits_data = ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_vga_valid = hInRange & vInRange; // @[src/main/scala/device/AXI4VGA.scala 148:28]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_aw_valid = io_in_ctrl_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_w_valid = io_in_ctrl_w_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_b_ready = io_in_ctrl_b_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_valid = io_in_ctrl_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_bits_addr = io_in_ctrl_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_r_ready = io_in_ctrl_r_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_aw_valid = io_in_fb_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_aw_bits_addr = io_in_fb_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_w_valid = io_in_fb_w_valid; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_data = io_in_fb_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_strb = io_in_fb_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_b_ready = io_in_fb_b_ready; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign fb_io_in_ar_valid = fb_io_in_ar_valid_REG & hCounterIs2; // @[src/main/scala/device/AXI4VGA.scala 162:43]
  assign fb_io_in_ar_bits_addr = {{13'd0}, _fb_io_in_ar_bits_addr_T_1}; // @[src/main/scala/device/AXI4VGA.scala 161:25]
  assign fb_io_in_r_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 164:20]
  assign fbHelper_clk = clock; // @[src/main/scala/device/AXI4VGA.scala 172:21]
  assign fbHelper_valid = io_vga_valid; // @[src/main/scala/device/AXI4VGA.scala 173:23]
  assign fbHelper_pixel = hCounter[1] ? _GEN_25[63:32] : _GEN_25[31:0]; // @[src/main/scala/device/AXI4VGA.scala 167:23]
  assign fbHelper_sync = ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 175:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_fb_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_fb_r_valid_r <= _GEN_12;
    end
    line_1826_valid_reg <= _io_in_fb_r_valid_T_1;
    line_1827_valid_reg <= _io_in_fb_r_valid_T;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
    end else begin
      hCounter <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    line_1828_valid_reg <= wrap_wrap;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (wrap_wrap_1) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        vCounter <= _wrap_value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    line_1829_valid_reg <= wrap_wrap;
    line_1830_valid_reg <= wrap_wrap_1;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV0_T_1) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV0_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV0 <= _fbPixelAddrV0_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    line_1831_valid_reg <= _fbPixelAddrV0_T_1;
    line_1832_valid_reg <= fbPixelAddrV0_wrap_wrap;
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV1_T) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV1_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV1 <= _fbPixelAddrV1_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    line_1833_valid_reg <= _fbPixelAddrV1_T;
    line_1834_valid_reg <= fbPixelAddrV1_wrap_wrap;
    fb_io_in_ar_valid_REG <= _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_data_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= fb_io_in_r_bits_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    line_1835_valid_reg <= _data_T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_in_fb_r_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1826_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1827_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  hCounter = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  line_1828_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vCounter = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  line_1829_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1830_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  line_1831_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1832_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  line_1833_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1834_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fb_io_in_ar_valid_REG = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  data_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  line_1835_valid_reg = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_io_in_fb_r_valid_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_fb_r_valid_T) begin
      cover(1'h1);
    end
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (wrap_wrap) begin
      cover(1'h1);
    end
    //
    if (wrap_wrap) begin
      cover(1'h1);
    end
    //
    if (wrap_wrap & wrap_wrap_1) begin
      cover(1'h1);
    end
    //
    if (_fbPixelAddrV0_T_1) begin
      cover(1'h1);
    end
    //
    if (_fbPixelAddrV0_T_1 & fbPixelAddrV0_wrap_wrap) begin
      cover(1'h1);
    end
    //
    if (_fbPixelAddrV1_T) begin
      cover(1'h1);
    end
    //
    if (_fbPixelAddrV1_T & fbPixelAddrV1_wrap_wrap) begin
      cover(1'h1);
    end
    //
    if (_data_T) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4Flash(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1836_clock;
  wire  line_1836_reset;
  wire  line_1836_valid;
  reg  line_1836_valid_reg;
  wire  _GEN_9 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1837_clock;
  wire  line_1837_reset;
  wire  line_1837_valid;
  reg  line_1837_valid_reg;
  wire  _GEN_10 = _r_busy_T | _GEN_9; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1838_clock;
  wire  line_1838_reset;
  wire  line_1838_valid;
  reg  line_1838_valid_reg;
  wire  _GEN_11 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1839_clock;
  wire  line_1839_reset;
  wire  line_1839_valid;
  reg  line_1839_valid_reg;
  wire  _GEN_12 = _io_in_r_valid_T_2 | _GEN_11; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1840_clock;
  wire  line_1840_reset;
  wire  line_1840_valid;
  reg  line_1840_valid_reg;
  wire  _GEN_13 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1841_clock;
  wire  line_1841_reset;
  wire  line_1841_valid;
  reg  line_1841_valid_reg;
  wire  _GEN_14 = _w_busy_T | _GEN_13; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1842_clock;
  wire  line_1842_reset;
  wire  line_1842_valid;
  reg  line_1842_valid_reg;
  wire  _GEN_15 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1843_clock;
  wire  line_1843_reset;
  wire  line_1843_valid;
  reg  line_1843_valid_reg;
  wire  _GEN_16 = _io_in_b_valid_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _rdata_T = 11'h0 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 11'h1 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 11'h2 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [20:0] _rdata_T_3 = _rdata_T ? 21'h10029b : 21'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_4 = _rdata_T_1 ? 25'h1f29293 : 25'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [17:0] _rdata_T_5 = _rdata_T_2 ? 18'h28067 : 18'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_18 = {{4'd0}, _rdata_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_6 = _GEN_18 | _rdata_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_19 = {{7'd0}, _rdata_T_5}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_7 = _rdata_T_6 | _GEN_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = {{39'd0}, _rdata_T_7}; // @[src/main/scala/device/AXI4Flash.scala 37:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  wire  line_1844_clock;
  wire  line_1844_reset;
  wire  line_1844_valid;
  reg  line_1844_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1836)) line_1836 (
    .clock(line_1836_clock),
    .reset(line_1836_reset),
    .valid(line_1836_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1837)) line_1837 (
    .clock(line_1837_clock),
    .reset(line_1837_reset),
    .valid(line_1837_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1838)) line_1838 (
    .clock(line_1838_clock),
    .reset(line_1838_reset),
    .valid(line_1838_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1839)) line_1839 (
    .clock(line_1839_clock),
    .reset(line_1839_reset),
    .valid(line_1839_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1840)) line_1840 (
    .clock(line_1840_clock),
    .reset(line_1840_reset),
    .valid(line_1840_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1841)) line_1841 (
    .clock(line_1841_clock),
    .reset(line_1841_reset),
    .valid(line_1841_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1842)) line_1842 (
    .clock(line_1842_clock),
    .reset(line_1842_reset),
    .valid(line_1842_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1843)) line_1843 (
    .clock(line_1843_clock),
    .reset(line_1843_reset),
    .valid(line_1843_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1844)) line_1844 (
    .clock(line_1844_clock),
    .reset(line_1844_reset),
    .valid(line_1844_valid)
  );
  assign line_1836_clock = clock;
  assign line_1836_reset = reset;
  assign line_1836_valid = _r_busy_T_1 ^ line_1836_valid_reg;
  assign line_1837_clock = clock;
  assign line_1837_reset = reset;
  assign line_1837_valid = _r_busy_T ^ line_1837_valid_reg;
  assign line_1838_clock = clock;
  assign line_1838_reset = reset;
  assign line_1838_valid = _r_busy_T_1 ^ line_1838_valid_reg;
  assign line_1839_clock = clock;
  assign line_1839_reset = reset;
  assign line_1839_valid = _io_in_r_valid_T_2 ^ line_1839_valid_reg;
  assign line_1840_clock = clock;
  assign line_1840_reset = reset;
  assign line_1840_valid = _w_busy_T_1 ^ line_1840_valid_reg;
  assign line_1841_clock = clock;
  assign line_1841_reset = reset;
  assign line_1841_valid = _w_busy_T ^ line_1841_valid_reg;
  assign line_1842_clock = clock;
  assign line_1842_reset = reset;
  assign line_1842_valid = _w_busy_T_1 ^ line_1842_valid_reg;
  assign line_1843_clock = clock;
  assign line_1843_reset = reset;
  assign line_1843_valid = _io_in_b_valid_T ^ line_1843_valid_reg;
  assign line_1844_clock = clock;
  assign line_1844_reset = reset;
  assign line_1844_valid = ren_REG ^ line_1844_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_10;
    end
    line_1836_valid_reg <= _r_busy_T_1;
    line_1837_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_12;
    end
    line_1838_valid_reg <= _r_busy_T_1;
    line_1839_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_14;
    end
    line_1840_valid_reg <= _w_busy_T_1;
    line_1841_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_16;
    end
    line_1842_valid_reg <= _w_busy_T_1;
    line_1843_valid_reg <= _io_in_b_valid_T;
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4Flash.scala 41:43]
    if (ren_REG) begin // @[src/main/scala/device/AXI4Flash.scala 41:30]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    line_1844_valid_reg <= ren_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1836_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1837_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1838_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1839_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1840_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1841_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1842_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1843_valid_reg = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  line_1844_valid_reg = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (ren_REG) begin
      cover(1'h1);
    end
  end
endmodule
module AXI4DummySD(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  sdHelper_clk; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_ren; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_data; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_setAddr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_addr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1845_clock;
  wire  line_1845_reset;
  wire  line_1845_valid;
  reg  line_1845_valid_reg;
  wire  _GEN_23 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1846_clock;
  wire  line_1846_reset;
  wire  line_1846_valid;
  reg  line_1846_valid_reg;
  wire  _GEN_24 = _r_busy_T | _GEN_23; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1847_clock;
  wire  line_1847_reset;
  wire  line_1847_valid;
  reg  line_1847_valid_reg;
  wire  _GEN_25 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1848_clock;
  wire  line_1848_reset;
  wire  line_1848_valid;
  reg  line_1848_valid_reg;
  wire  _GEN_26 = _io_in_r_valid_T_2 | _GEN_25; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1849_clock;
  wire  line_1849_reset;
  wire  line_1849_valid;
  reg  line_1849_valid_reg;
  wire  _GEN_27 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1850_clock;
  wire  line_1850_reset;
  wire  line_1850_valid;
  reg  line_1850_valid_reg;
  wire  _GEN_28 = _w_busy_T | _GEN_27; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1851_clock;
  wire  line_1851_reset;
  wire  line_1851_valid;
  reg  line_1851_valid_reg;
  wire  _GEN_29 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  line_1852_clock;
  wire  line_1852_reset;
  wire  line_1852_valid;
  reg  line_1852_valid_reg;
  wire  _GEN_30 = _io_in_b_valid_T | _GEN_29; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] regs_0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_1; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_4; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_5; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_6; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_7; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_8; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_15; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_20; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [3:0] strb = io_in_aw_bits_addr[2] ? io_in_w_bits_strb[7:4] : io_in_w_bits_strb[3:0]; // @[src/main/scala/device/AXI4DummySD.scala 138:22]
  wire [7:0] _T_8 = strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_9 = strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_10 = strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_11 = strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [31:0] _T_12 = {_T_11,_T_10,_T_9,_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T = 13'h0 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 13'h38 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 13'h18 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 13'h34 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 13'h14 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_5 = 13'h1c == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_6 = 13'h50 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_7 = 13'h10 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_8 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_9 = 13'h20 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_10 = 13'h40 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_11 = _rdata_T ? regs_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_1 ? regs_15 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_13 = _rdata_T_2 ? regs_6 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdata_T_14 = _rdata_T_3 ? 8'h80 : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_15 = _rdata_T_4 ? regs_5 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_16 = _rdata_T_5 ? regs_7 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_17 = _rdata_T_6 ? regs_20 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_18 = _rdata_T_7 ? regs_4 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_19 = _rdata_T_8 ? regs_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_20 = _rdata_T_9 ? regs_8 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_21 = _rdata_T_10 ? sdHelper_data : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_22 = _rdata_T_11 | _rdata_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_23 = _rdata_T_22 | _rdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_63 = {{24'd0}, _rdata_T_14}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_24 = _rdata_T_23 | _GEN_63; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_25 = _rdata_T_24 | _rdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_26 = _rdata_T_25 | _rdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_27 = _rdata_T_26 | _rdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_28 = _rdata_T_27 | _rdata_T_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_29 = _rdata_T_28 | _rdata_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_30 = _rdata_T_29 | _rdata_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_31 = _rdata_T_30 | _rdata_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_14 = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1853_clock;
  wire  line_1853_reset;
  wire  line_1853_valid;
  reg  line_1853_valid_reg;
  wire [31:0] _regs_0_T = io_in_w_bits_data[31:0] & _T_12; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _regs_0_T_1 = ~_T_12; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _regs_0_T_2 = regs_0 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_0_T_3 = _regs_0_T | _regs_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [5:0] regs_0_cmd = _regs_0_T_3[5:0]; // @[src/main/scala/device/AXI4DummySD.scala 84:20]
  wire  _regs_0_T_4 = 6'h1 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18]
  wire  line_1854_clock;
  wire  line_1854_reset;
  wire  line_1854_valid;
  reg  line_1854_valid_reg;
  wire  line_1855_clock;
  wire  line_1855_reset;
  wire  line_1855_valid;
  reg  line_1855_valid_reg;
  wire  _regs_0_T_5 = 6'h2 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18]
  wire  line_1856_clock;
  wire  line_1856_reset;
  wire  line_1856_valid;
  reg  line_1856_valid_reg;
  wire  line_1857_clock;
  wire  line_1857_reset;
  wire  line_1857_valid;
  reg  line_1857_valid_reg;
  wire  _regs_0_T_6 = 6'h9 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18]
  wire  line_1858_clock;
  wire  line_1858_reset;
  wire  line_1858_valid;
  reg  line_1858_valid_reg;
  wire  line_1859_clock;
  wire  line_1859_reset;
  wire  line_1859_valid;
  reg  line_1859_valid_reg;
  wire  _regs_0_T_7 = 6'hd == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18]
  wire  line_1860_clock;
  wire  line_1860_reset;
  wire  line_1860_valid;
  reg  line_1860_valid_reg;
  wire  line_1861_clock;
  wire  line_1861_reset;
  wire  line_1861_valid;
  reg  line_1861_valid_reg;
  wire  _regs_0_T_8 = 6'h12 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18]
  wire  line_1862_clock;
  wire  line_1862_reset;
  wire  line_1862_valid;
  reg  line_1862_valid_reg;
  wire [31:0] _GEN_32 = 6'hd == regs_0_cmd ? 32'h0 : regs_4; // @[src/main/scala/device/AXI4DummySD.scala 85:18 102:22 72:43]
  wire [31:0] _GEN_33 = 6'hd == regs_0_cmd ? 32'h0 : regs_5; // @[src/main/scala/device/AXI4DummySD.scala 85:18 103:22 72:43]
  wire [31:0] _GEN_34 = 6'hd == regs_0_cmd ? 32'h0 : regs_6; // @[src/main/scala/device/AXI4DummySD.scala 85:18 104:22 72:43]
  wire [31:0] _GEN_35 = 6'hd == regs_0_cmd ? 32'h0 : regs_7; // @[src/main/scala/device/AXI4DummySD.scala 85:18 105:22 72:43]
  wire  _GEN_36 = 6'hd == regs_0_cmd ? 1'h0 : 6'h12 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire [31:0] _GEN_37 = 6'h9 == regs_0_cmd ? 32'h92404001 : _GEN_32; // @[src/main/scala/device/AXI4DummySD.scala 85:18 96:22]
  wire [31:0] _GEN_38 = 6'h9 == regs_0_cmd ? 32'hd24b97e3 : _GEN_33; // @[src/main/scala/device/AXI4DummySD.scala 85:18 97:22]
  wire [31:0] _GEN_39 = 6'h9 == regs_0_cmd ? 32'hf5f803f : _GEN_34; // @[src/main/scala/device/AXI4DummySD.scala 85:18 98:22]
  wire [31:0] _GEN_40 = 6'h9 == regs_0_cmd ? 32'h8c26012a : _GEN_35; // @[src/main/scala/device/AXI4DummySD.scala 85:18 99:22]
  wire  _GEN_41 = 6'h9 == regs_0_cmd ? 1'h0 : _GEN_36; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_46 = 6'h2 == regs_0_cmd ? 1'h0 : _GEN_41; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_51 = 6'h1 == regs_0_cmd ? 1'h0 : _GEN_46; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _T_16 = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h38; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1863_clock;
  wire  line_1863_reset;
  wire  line_1863_valid;
  reg  line_1863_valid_reg;
  wire [31:0] _regs_15_T_2 = regs_15 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_15_T_3 = _regs_0_T | _regs_15_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_18 = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h50; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1864_clock;
  wire  line_1864_reset;
  wire  line_1864_valid;
  reg  line_1864_valid_reg;
  wire [31:0] _regs_20_T_2 = regs_20 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_20_T_3 = _regs_0_T | _regs_20_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_20 = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h4; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1865_clock;
  wire  line_1865_reset;
  wire  line_1865_valid;
  reg  line_1865_valid_reg;
  wire [31:0] _regs_1_T_2 = regs_1 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_1_T_3 = _regs_0_T | _regs_1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_22 = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h20; // @[src/main/scala/utils/RegMap.scala 32:32]
  wire  line_1866_clock;
  wire  line_1866_reset;
  wire  line_1866_valid;
  reg  line_1866_valid_reg;
  wire [31:0] _regs_8_T_2 = regs_8 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_8_T_3 = _regs_0_T | _regs_8_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] rdata = {{32'd0}, _rdata_T_31}; // @[src/main/scala/device/AXI4DummySD.scala 139:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
  wire  line_1867_clock;
  wire  line_1867_reset;
  wire  line_1867_valid;
  reg  line_1867_valid_reg;
  SDHelper sdHelper ( // @[src/main/scala/device/AXI4DummySD.scala 114:24]
    .clk(sdHelper_clk),
    .ren(sdHelper_ren),
    .data(sdHelper_data),
    .setAddr(sdHelper_setAddr),
    .addr(sdHelper_addr)
  );
  GEN_w1_line #(.COVER_INDEX(1845)) line_1845 (
    .clock(line_1845_clock),
    .reset(line_1845_reset),
    .valid(line_1845_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1846)) line_1846 (
    .clock(line_1846_clock),
    .reset(line_1846_reset),
    .valid(line_1846_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1847)) line_1847 (
    .clock(line_1847_clock),
    .reset(line_1847_reset),
    .valid(line_1847_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1848)) line_1848 (
    .clock(line_1848_clock),
    .reset(line_1848_reset),
    .valid(line_1848_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1849)) line_1849 (
    .clock(line_1849_clock),
    .reset(line_1849_reset),
    .valid(line_1849_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1850)) line_1850 (
    .clock(line_1850_clock),
    .reset(line_1850_reset),
    .valid(line_1850_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1851)) line_1851 (
    .clock(line_1851_clock),
    .reset(line_1851_reset),
    .valid(line_1851_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1852)) line_1852 (
    .clock(line_1852_clock),
    .reset(line_1852_reset),
    .valid(line_1852_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1853)) line_1853 (
    .clock(line_1853_clock),
    .reset(line_1853_reset),
    .valid(line_1853_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1854)) line_1854 (
    .clock(line_1854_clock),
    .reset(line_1854_reset),
    .valid(line_1854_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1855)) line_1855 (
    .clock(line_1855_clock),
    .reset(line_1855_reset),
    .valid(line_1855_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1856)) line_1856 (
    .clock(line_1856_clock),
    .reset(line_1856_reset),
    .valid(line_1856_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1857)) line_1857 (
    .clock(line_1857_clock),
    .reset(line_1857_reset),
    .valid(line_1857_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1858)) line_1858 (
    .clock(line_1858_clock),
    .reset(line_1858_reset),
    .valid(line_1858_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1859)) line_1859 (
    .clock(line_1859_clock),
    .reset(line_1859_reset),
    .valid(line_1859_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1860)) line_1860 (
    .clock(line_1860_clock),
    .reset(line_1860_reset),
    .valid(line_1860_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1861)) line_1861 (
    .clock(line_1861_clock),
    .reset(line_1861_reset),
    .valid(line_1861_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1862)) line_1862 (
    .clock(line_1862_clock),
    .reset(line_1862_reset),
    .valid(line_1862_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1863)) line_1863 (
    .clock(line_1863_clock),
    .reset(line_1863_reset),
    .valid(line_1863_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1864)) line_1864 (
    .clock(line_1864_clock),
    .reset(line_1864_reset),
    .valid(line_1864_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1865)) line_1865 (
    .clock(line_1865_clock),
    .reset(line_1865_reset),
    .valid(line_1865_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1866)) line_1866 (
    .clock(line_1866_clock),
    .reset(line_1866_reset),
    .valid(line_1866_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1867)) line_1867 (
    .clock(line_1867_clock),
    .reset(line_1867_reset),
    .valid(line_1867_valid)
  );
  assign line_1845_clock = clock;
  assign line_1845_reset = reset;
  assign line_1845_valid = _r_busy_T_1 ^ line_1845_valid_reg;
  assign line_1846_clock = clock;
  assign line_1846_reset = reset;
  assign line_1846_valid = _r_busy_T ^ line_1846_valid_reg;
  assign line_1847_clock = clock;
  assign line_1847_reset = reset;
  assign line_1847_valid = _r_busy_T_1 ^ line_1847_valid_reg;
  assign line_1848_clock = clock;
  assign line_1848_reset = reset;
  assign line_1848_valid = _io_in_r_valid_T_2 ^ line_1848_valid_reg;
  assign line_1849_clock = clock;
  assign line_1849_reset = reset;
  assign line_1849_valid = _w_busy_T_1 ^ line_1849_valid_reg;
  assign line_1850_clock = clock;
  assign line_1850_reset = reset;
  assign line_1850_valid = _w_busy_T ^ line_1850_valid_reg;
  assign line_1851_clock = clock;
  assign line_1851_reset = reset;
  assign line_1851_valid = _w_busy_T_1 ^ line_1851_valid_reg;
  assign line_1852_clock = clock;
  assign line_1852_reset = reset;
  assign line_1852_valid = _io_in_b_valid_T ^ line_1852_valid_reg;
  assign line_1853_clock = clock;
  assign line_1853_reset = reset;
  assign line_1853_valid = _T_14 ^ line_1853_valid_reg;
  assign line_1854_clock = clock;
  assign line_1854_reset = reset;
  assign line_1854_valid = _regs_0_T_4 ^ line_1854_valid_reg;
  assign line_1855_clock = clock;
  assign line_1855_reset = reset;
  assign line_1855_valid = _regs_0_T_4 ^ line_1855_valid_reg;
  assign line_1856_clock = clock;
  assign line_1856_reset = reset;
  assign line_1856_valid = _regs_0_T_5 ^ line_1856_valid_reg;
  assign line_1857_clock = clock;
  assign line_1857_reset = reset;
  assign line_1857_valid = _regs_0_T_5 ^ line_1857_valid_reg;
  assign line_1858_clock = clock;
  assign line_1858_reset = reset;
  assign line_1858_valid = _regs_0_T_6 ^ line_1858_valid_reg;
  assign line_1859_clock = clock;
  assign line_1859_reset = reset;
  assign line_1859_valid = _regs_0_T_6 ^ line_1859_valid_reg;
  assign line_1860_clock = clock;
  assign line_1860_reset = reset;
  assign line_1860_valid = _regs_0_T_7 ^ line_1860_valid_reg;
  assign line_1861_clock = clock;
  assign line_1861_reset = reset;
  assign line_1861_valid = _regs_0_T_7 ^ line_1861_valid_reg;
  assign line_1862_clock = clock;
  assign line_1862_reset = reset;
  assign line_1862_valid = _regs_0_T_8 ^ line_1862_valid_reg;
  assign line_1863_clock = clock;
  assign line_1863_reset = reset;
  assign line_1863_valid = _T_16 ^ line_1863_valid_reg;
  assign line_1864_clock = clock;
  assign line_1864_reset = reset;
  assign line_1864_valid = _T_18 ^ line_1864_valid_reg;
  assign line_1865_clock = clock;
  assign line_1865_reset = reset;
  assign line_1865_valid = _T_20 ^ line_1865_valid_reg;
  assign line_1866_clock = clock;
  assign line_1866_reset = reset;
  assign line_1866_valid = _T_22 ^ line_1866_valid_reg;
  assign line_1867_clock = clock;
  assign line_1867_reset = reset;
  assign line_1867_valid = ren_REG ^ line_1867_valid_reg;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 143:18]
  assign sdHelper_clk = clock; // @[src/main/scala/device/AXI4DummySD.scala 115:19]
  assign sdHelper_ren = io_in_ar_bits_addr[12:0] == 13'h40 & _r_busy_T; // @[src/main/scala/device/AXI4DummySD.scala 116:51]
  assign sdHelper_setAddr = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0 & _GEN_51; // @[src/main/scala/utils/RegMap.scala 32:48 src/main/scala/device/AXI4DummySD.scala 81:25]
  assign sdHelper_addr = regs_1; // @[src/main/scala/device/AXI4DummySD.scala 118:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_24;
    end
    line_1845_valid_reg <= _r_busy_T_1;
    line_1846_valid_reg <= _r_busy_T;
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_26;
    end
    line_1847_valid_reg <= _r_busy_T_1;
    line_1848_valid_reg <= _io_in_r_valid_T_2;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_28;
    end
    line_1849_valid_reg <= _w_busy_T_1;
    line_1850_valid_reg <= _w_busy_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_30;
    end
    line_1851_valid_reg <= _w_busy_T_1;
    line_1852_valid_reg <= _io_in_b_valid_T;
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_0 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_0 <= _regs_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_1 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_1 <= _regs_1_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_4 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (6'h1 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h80ff8000; // @[src/main/scala/device/AXI4DummySD.scala 87:22]
      end else if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h1; // @[src/main/scala/device/AXI4DummySD.scala 90:22]
      end else begin
        regs_4 <= _GEN_37;
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 91:22]
        end else begin
          regs_5 <= _GEN_38;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 92:22]
        end else begin
          regs_6 <= _GEN_39;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_7 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_7 <= 32'h15000000; // @[src/main/scala/device/AXI4DummySD.scala 93:22]
        end else begin
          regs_7 <= _GEN_40;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_8 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h20) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_8 <= _regs_8_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_15 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h38) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_15 <= _regs_15_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_20 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h50) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_20 <= _regs_20_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    line_1853_valid_reg <= _T_14;
    line_1854_valid_reg <= _regs_0_T_4;
    line_1855_valid_reg <= _regs_0_T_4;
    line_1856_valid_reg <= _regs_0_T_5;
    line_1857_valid_reg <= _regs_0_T_5;
    line_1858_valid_reg <= _regs_0_T_6;
    line_1859_valid_reg <= _regs_0_T_6;
    line_1860_valid_reg <= _regs_0_T_7;
    line_1861_valid_reg <= _regs_0_T_7;
    line_1862_valid_reg <= _regs_0_T_8;
    line_1863_valid_reg <= _T_16;
    line_1864_valid_reg <= _T_18;
    line_1865_valid_reg <= _T_20;
    line_1866_valid_reg <= _T_22;
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4DummySD.scala 144:49]
    if (ren_REG) begin // @[src/main/scala/device/AXI4DummySD.scala 144:36]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    line_1867_valid_reg <= ren_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1845_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1846_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ren_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1847_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1848_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  w_busy = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1849_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1850_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1851_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1852_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regs_0 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_4 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_5 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_6 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_7 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_8 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_15 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_20 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  line_1853_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_1854_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_1855_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_1856_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_1857_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_1858_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_1859_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_1860_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_1861_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_1862_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_1863_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_1864_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_1865_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_1866_valid_reg = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  line_1867_valid_reg = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T) begin
      cover(1'h1);
    end
    //
    if (_r_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_r_valid_T_2) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T) begin
      cover(1'h1);
    end
    //
    if (_w_busy_T_1) begin
      cover(1'h1);
    end
    //
    if (_io_in_b_valid_T) begin
      cover(1'h1);
    end
    //
    if (_T_14) begin
      cover(1'h1);
    end
    //
    if (_T_14 & _regs_0_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & _regs_0_T_5) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5 & _regs_0_T_6) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5 & ~_regs_0_T_6) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5 & ~_regs_0_T_6 & _regs_0_T_7) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5 & ~_regs_0_T_6 & ~_regs_0_T_7) begin
      cover(1'h1);
    end
    //
    if (_T_14 & ~_regs_0_T_4 & ~_regs_0_T_5 & ~_regs_0_T_6 & ~_regs_0_T_7 & _regs_0_T_8) begin
      cover(1'h1);
    end
    //
    if (_T_16) begin
      cover(1'h1);
    end
    //
    if (_T_18) begin
      cover(1'h1);
    end
    //
    if (_T_20) begin
      cover(1'h1);
    end
    //
    if (_T_22) begin
      cover(1'h1);
    end
    //
    if (ren_REG) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_3(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1868_clock;
  wire  line_1868_reset;
  wire  line_1868_valid;
  reg  line_1868_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1869_clock;
  wire  line_1869_reset;
  wire  line_1869_valid;
  reg  line_1869_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1870_clock;
  wire  line_1870_reset;
  wire  line_1870_valid;
  reg  line_1870_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1871_clock;
  wire  line_1871_reset;
  wire  line_1871_valid;
  reg  line_1871_valid_reg;
  wire  line_1872_clock;
  wire  line_1872_reset;
  wire  line_1872_valid;
  reg  line_1872_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1873_clock;
  wire  line_1873_reset;
  wire  line_1873_valid;
  reg  line_1873_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1874_clock;
  wire  line_1874_reset;
  wire  line_1874_valid;
  reg  line_1874_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1868)) line_1868 (
    .clock(line_1868_clock),
    .reset(line_1868_reset),
    .valid(line_1868_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1869)) line_1869 (
    .clock(line_1869_clock),
    .reset(line_1869_reset),
    .valid(line_1869_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1870)) line_1870 (
    .clock(line_1870_clock),
    .reset(line_1870_reset),
    .valid(line_1870_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1871)) line_1871 (
    .clock(line_1871_clock),
    .reset(line_1871_reset),
    .valid(line_1871_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1872)) line_1872 (
    .clock(line_1872_clock),
    .reset(line_1872_reset),
    .valid(line_1872_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1873)) line_1873 (
    .clock(line_1873_clock),
    .reset(line_1873_reset),
    .valid(line_1873_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1874)) line_1874 (
    .clock(line_1874_clock),
    .reset(line_1874_reset),
    .valid(line_1874_valid)
  );
  assign line_1868_clock = clock;
  assign line_1868_reset = reset;
  assign line_1868_valid = _T_2 ^ line_1868_valid_reg;
  assign line_1869_clock = clock;
  assign line_1869_reset = reset;
  assign line_1869_valid = _T_3 ^ line_1869_valid_reg;
  assign line_1870_clock = clock;
  assign line_1870_reset = reset;
  assign line_1870_valid = _awAck_T ^ line_1870_valid_reg;
  assign line_1871_clock = clock;
  assign line_1871_reset = reset;
  assign line_1871_valid = wSend ^ line_1871_valid_reg;
  assign line_1872_clock = clock;
  assign line_1872_reset = reset;
  assign line_1872_valid = _wSend_T_1 ^ line_1872_valid_reg;
  assign line_1873_clock = clock;
  assign line_1873_reset = reset;
  assign line_1873_valid = wSend ^ line_1873_valid_reg;
  assign line_1874_clock = clock;
  assign line_1874_reset = reset;
  assign line_1874_valid = _wen_T_1 ^ line_1874_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1868_valid_reg <= _T_2;
    line_1869_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1870_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1871_valid_reg <= wSend;
    line_1872_valid_reg <= _wSend_T_1;
    line_1873_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1874_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1868_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1869_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1870_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1871_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1872_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1873_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1874_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_4(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1875_clock;
  wire  line_1875_reset;
  wire  line_1875_valid;
  reg  line_1875_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1876_clock;
  wire  line_1876_reset;
  wire  line_1876_valid;
  reg  line_1876_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1877_clock;
  wire  line_1877_reset;
  wire  line_1877_valid;
  reg  line_1877_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1878_clock;
  wire  line_1878_reset;
  wire  line_1878_valid;
  reg  line_1878_valid_reg;
  wire  line_1879_clock;
  wire  line_1879_reset;
  wire  line_1879_valid;
  reg  line_1879_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1880_clock;
  wire  line_1880_reset;
  wire  line_1880_valid;
  reg  line_1880_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1881_clock;
  wire  line_1881_reset;
  wire  line_1881_valid;
  reg  line_1881_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1875)) line_1875 (
    .clock(line_1875_clock),
    .reset(line_1875_reset),
    .valid(line_1875_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1876)) line_1876 (
    .clock(line_1876_clock),
    .reset(line_1876_reset),
    .valid(line_1876_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1877)) line_1877 (
    .clock(line_1877_clock),
    .reset(line_1877_reset),
    .valid(line_1877_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1878)) line_1878 (
    .clock(line_1878_clock),
    .reset(line_1878_reset),
    .valid(line_1878_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1879)) line_1879 (
    .clock(line_1879_clock),
    .reset(line_1879_reset),
    .valid(line_1879_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1880)) line_1880 (
    .clock(line_1880_clock),
    .reset(line_1880_reset),
    .valid(line_1880_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1881)) line_1881 (
    .clock(line_1881_clock),
    .reset(line_1881_reset),
    .valid(line_1881_valid)
  );
  assign line_1875_clock = clock;
  assign line_1875_reset = reset;
  assign line_1875_valid = _T_2 ^ line_1875_valid_reg;
  assign line_1876_clock = clock;
  assign line_1876_reset = reset;
  assign line_1876_valid = _T_3 ^ line_1876_valid_reg;
  assign line_1877_clock = clock;
  assign line_1877_reset = reset;
  assign line_1877_valid = _awAck_T ^ line_1877_valid_reg;
  assign line_1878_clock = clock;
  assign line_1878_reset = reset;
  assign line_1878_valid = wSend ^ line_1878_valid_reg;
  assign line_1879_clock = clock;
  assign line_1879_reset = reset;
  assign line_1879_valid = _wSend_T_1 ^ line_1879_valid_reg;
  assign line_1880_clock = clock;
  assign line_1880_reset = reset;
  assign line_1880_valid = wSend ^ line_1880_valid_reg;
  assign line_1881_clock = clock;
  assign line_1881_reset = reset;
  assign line_1881_valid = _wen_T_1 ^ line_1881_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : 1'h1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1875_valid_reg <= _T_2;
    line_1876_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1877_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1878_valid_reg <= wSend;
    line_1879_valid_reg <= _wSend_T_1;
    line_1880_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1881_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1875_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1876_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1877_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1878_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1879_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1880_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1881_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_5(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1882_clock;
  wire  line_1882_reset;
  wire  line_1882_valid;
  reg  line_1882_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1883_clock;
  wire  line_1883_reset;
  wire  line_1883_valid;
  reg  line_1883_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1884_clock;
  wire  line_1884_reset;
  wire  line_1884_valid;
  reg  line_1884_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1885_clock;
  wire  line_1885_reset;
  wire  line_1885_valid;
  reg  line_1885_valid_reg;
  wire  line_1886_clock;
  wire  line_1886_reset;
  wire  line_1886_valid;
  reg  line_1886_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1887_clock;
  wire  line_1887_reset;
  wire  line_1887_valid;
  reg  line_1887_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1888_clock;
  wire  line_1888_reset;
  wire  line_1888_valid;
  reg  line_1888_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1882)) line_1882 (
    .clock(line_1882_clock),
    .reset(line_1882_reset),
    .valid(line_1882_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1883)) line_1883 (
    .clock(line_1883_clock),
    .reset(line_1883_reset),
    .valid(line_1883_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1884)) line_1884 (
    .clock(line_1884_clock),
    .reset(line_1884_reset),
    .valid(line_1884_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1885)) line_1885 (
    .clock(line_1885_clock),
    .reset(line_1885_reset),
    .valid(line_1885_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1886)) line_1886 (
    .clock(line_1886_clock),
    .reset(line_1886_reset),
    .valid(line_1886_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1887)) line_1887 (
    .clock(line_1887_clock),
    .reset(line_1887_reset),
    .valid(line_1887_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1888)) line_1888 (
    .clock(line_1888_clock),
    .reset(line_1888_reset),
    .valid(line_1888_valid)
  );
  assign line_1882_clock = clock;
  assign line_1882_reset = reset;
  assign line_1882_valid = _T_2 ^ line_1882_valid_reg;
  assign line_1883_clock = clock;
  assign line_1883_reset = reset;
  assign line_1883_valid = _T_3 ^ line_1883_valid_reg;
  assign line_1884_clock = clock;
  assign line_1884_reset = reset;
  assign line_1884_valid = _awAck_T ^ line_1884_valid_reg;
  assign line_1885_clock = clock;
  assign line_1885_reset = reset;
  assign line_1885_valid = wSend ^ line_1885_valid_reg;
  assign line_1886_clock = clock;
  assign line_1886_reset = reset;
  assign line_1886_valid = _wSend_T_1 ^ line_1886_valid_reg;
  assign line_1887_clock = clock;
  assign line_1887_reset = reset;
  assign line_1887_valid = wSend ^ line_1887_valid_reg;
  assign line_1888_clock = clock;
  assign line_1888_reset = reset;
  assign line_1888_valid = _wen_T_1 ^ line_1888_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1882_valid_reg <= _T_2;
    line_1883_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1884_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1885_valid_reg <= wSend;
    line_1886_valid_reg <= _wSend_T_1;
    line_1887_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1888_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1882_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1883_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1884_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1885_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1886_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1887_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1888_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_6(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1889_clock;
  wire  line_1889_reset;
  wire  line_1889_valid;
  reg  line_1889_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1890_clock;
  wire  line_1890_reset;
  wire  line_1890_valid;
  reg  line_1890_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1891_clock;
  wire  line_1891_reset;
  wire  line_1891_valid;
  reg  line_1891_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1892_clock;
  wire  line_1892_reset;
  wire  line_1892_valid;
  reg  line_1892_valid_reg;
  wire  line_1893_clock;
  wire  line_1893_reset;
  wire  line_1893_valid;
  reg  line_1893_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1894_clock;
  wire  line_1894_reset;
  wire  line_1894_valid;
  reg  line_1894_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1895_clock;
  wire  line_1895_reset;
  wire  line_1895_valid;
  reg  line_1895_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1889)) line_1889 (
    .clock(line_1889_clock),
    .reset(line_1889_reset),
    .valid(line_1889_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1890)) line_1890 (
    .clock(line_1890_clock),
    .reset(line_1890_reset),
    .valid(line_1890_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1891)) line_1891 (
    .clock(line_1891_clock),
    .reset(line_1891_reset),
    .valid(line_1891_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1892)) line_1892 (
    .clock(line_1892_clock),
    .reset(line_1892_reset),
    .valid(line_1892_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1893)) line_1893 (
    .clock(line_1893_clock),
    .reset(line_1893_reset),
    .valid(line_1893_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1894)) line_1894 (
    .clock(line_1894_clock),
    .reset(line_1894_reset),
    .valid(line_1894_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1895)) line_1895 (
    .clock(line_1895_clock),
    .reset(line_1895_reset),
    .valid(line_1895_valid)
  );
  assign line_1889_clock = clock;
  assign line_1889_reset = reset;
  assign line_1889_valid = _T_2 ^ line_1889_valid_reg;
  assign line_1890_clock = clock;
  assign line_1890_reset = reset;
  assign line_1890_valid = _T_3 ^ line_1890_valid_reg;
  assign line_1891_clock = clock;
  assign line_1891_reset = reset;
  assign line_1891_valid = _awAck_T ^ line_1891_valid_reg;
  assign line_1892_clock = clock;
  assign line_1892_reset = reset;
  assign line_1892_valid = wSend ^ line_1892_valid_reg;
  assign line_1893_clock = clock;
  assign line_1893_reset = reset;
  assign line_1893_valid = _wSend_T_1 ^ line_1893_valid_reg;
  assign line_1894_clock = clock;
  assign line_1894_reset = reset;
  assign line_1894_valid = wSend ^ line_1894_valid_reg;
  assign line_1895_clock = clock;
  assign line_1895_reset = reset;
  assign line_1895_valid = _wen_T_1 ^ line_1895_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1889_valid_reg <= _T_2;
    line_1890_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1891_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1892_valid_reg <= wSend;
    line_1893_valid_reg <= _wSend_T_1;
    line_1894_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1895_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1889_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1890_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1891_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1892_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1893_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1894_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1895_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimpleBus2AXI4Converter_7(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _T_2 = ~reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1896_clock;
  wire  line_1896_reset;
  wire  line_1896_valid;
  reg  line_1896_valid_reg;
  wire  _T_3 = ~toAXI4Lite; // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
  wire  line_1897_clock;
  wire  line_1897_reset;
  wire  line_1897_valid;
  reg  line_1897_valid_reg;
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  line_1898_clock;
  wire  line_1898_reset;
  wire  line_1898_valid;
  reg  line_1898_valid_reg;
  wire  _GEN_7 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  line_1899_clock;
  wire  line_1899_reset;
  wire  line_1899_valid;
  reg  line_1899_valid_reg;
  wire  line_1900_clock;
  wire  line_1900_reset;
  wire  line_1900_valid;
  reg  line_1900_valid_reg;
  wire  _GEN_9 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  line_1901_clock;
  wire  line_1901_reset;
  wire  line_1901_valid;
  reg  line_1901_valid_reg;
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  line_1902_clock;
  wire  line_1902_reset;
  wire  line_1902_valid;
  reg  line_1902_valid_reg;
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  GEN_w1_line #(.COVER_INDEX(1896)) line_1896 (
    .clock(line_1896_clock),
    .reset(line_1896_reset),
    .valid(line_1896_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1897)) line_1897 (
    .clock(line_1897_clock),
    .reset(line_1897_reset),
    .valid(line_1897_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1898)) line_1898 (
    .clock(line_1898_clock),
    .reset(line_1898_reset),
    .valid(line_1898_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1899)) line_1899 (
    .clock(line_1899_clock),
    .reset(line_1899_reset),
    .valid(line_1899_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1900)) line_1900 (
    .clock(line_1900_clock),
    .reset(line_1900_reset),
    .valid(line_1900_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1901)) line_1901 (
    .clock(line_1901_clock),
    .reset(line_1901_reset),
    .valid(line_1901_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1902)) line_1902 (
    .clock(line_1902_clock),
    .reset(line_1902_reset),
    .valid(line_1902_valid)
  );
  assign line_1896_clock = clock;
  assign line_1896_reset = reset;
  assign line_1896_valid = _T_2 ^ line_1896_valid_reg;
  assign line_1897_clock = clock;
  assign line_1897_reset = reset;
  assign line_1897_valid = _T_3 ^ line_1897_valid_reg;
  assign line_1898_clock = clock;
  assign line_1898_reset = reset;
  assign line_1898_valid = _awAck_T ^ line_1898_valid_reg;
  assign line_1899_clock = clock;
  assign line_1899_reset = reset;
  assign line_1899_valid = wSend ^ line_1899_valid_reg;
  assign line_1900_clock = clock;
  assign line_1900_reset = reset;
  assign line_1900_valid = _wSend_T_1 ^ line_1900_valid_reg;
  assign line_1901_clock = clock;
  assign line_1901_reset = reset;
  assign line_1901_valid = wSend ^ line_1901_valid_reg;
  assign line_1902_clock = clock;
  assign line_1902_reset = reset;
  assign line_1902_valid = _wen_T_1 ^ line_1902_valid_reg;
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    line_1896_valid_reg <= _T_2;
    line_1897_valid_reg <= _T_3;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_7;
    end
    line_1898_valid_reg <= _awAck_T;
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_9;
    end
    line_1899_valid_reg <= wSend;
    line_1900_valid_reg <= _wSend_T_1;
    line_1901_valid_reg <= wSend;
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    line_1902_valid_reg <= _wen_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1896_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1897_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  awAck = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1898_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wAck = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1899_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1900_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1901_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wen = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1902_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_2) begin
      cover(1'h1);
    end
    //
    if (_T_2 & _T_3) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (_awAck_T) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wSend_T_1) begin
      cover(1'h1);
    end
    //
    if (wSend) begin
      cover(1'h1);
    end
    //
    if (_wen_T_1) begin
      cover(1'h1);
    end
  end
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_rw_req_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_req_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [31:0] io_rw_req_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [3:0]  io_rw_req_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_rw_req_bits_wmask, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [63:0] io_rw_req_bits_wdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_resp_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_rw_resp_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [3:0]  io_rw_resp_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [63:0] io_rw_resp_bits_rdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_out_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_uart_out_ch, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_in_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_uart_in_ch // @[src/main/scala/sim/SimMMIO.scala 28:14]
);
  wire  xbar_clock; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_reset; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_in_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_in_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_0_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_0_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_0_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_1_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_1_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_1_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_2_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_2_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_3_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_3_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_4_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_4_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_4_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  uart_clock; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_reset; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_in_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  vga_clock; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_reset; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_fb_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_fb_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [7:0] vga_io_in_fb_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_ctrl_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_vga_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  flash_clock; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_reset; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [31:0] flash_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [63:0] flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  sd_clock; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_reset; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [7:0] sd_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  uart_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] uart_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_fb_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_ctrl_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] flash_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] sd_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  SimpleBusCrossbar1toN_1 xbar ( // @[src/main/scala/sim/SimMMIO.scala 45:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_req_ready(xbar_io_in_req_ready),
    .io_in_req_valid(xbar_io_in_req_valid),
    .io_in_req_bits_addr(xbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(xbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(xbar_io_in_req_bits_wdata),
    .io_in_resp_ready(xbar_io_in_resp_ready),
    .io_in_resp_valid(xbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(xbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(xbar_io_out_0_req_ready),
    .io_out_0_req_valid(xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(xbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(xbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(xbar_io_out_1_req_ready),
    .io_out_1_req_valid(xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(xbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(xbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(xbar_io_out_1_resp_valid),
    .io_out_2_req_ready(xbar_io_out_2_req_ready),
    .io_out_2_req_valid(xbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(xbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(xbar_io_out_2_req_bits_cmd),
    .io_out_2_resp_ready(xbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(xbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(xbar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(xbar_io_out_3_req_ready),
    .io_out_3_req_valid(xbar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(xbar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_cmd(xbar_io_out_3_req_bits_cmd),
    .io_out_3_resp_ready(xbar_io_out_3_resp_ready),
    .io_out_3_resp_valid(xbar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(xbar_io_out_3_resp_bits_rdata),
    .io_out_4_req_ready(xbar_io_out_4_req_ready),
    .io_out_4_req_valid(xbar_io_out_4_req_valid),
    .io_out_4_req_bits_addr(xbar_io_out_4_req_bits_addr),
    .io_out_4_req_bits_cmd(xbar_io_out_4_req_bits_cmd),
    .io_out_4_req_bits_wmask(xbar_io_out_4_req_bits_wmask),
    .io_out_4_req_bits_wdata(xbar_io_out_4_req_bits_wdata),
    .io_out_4_resp_ready(xbar_io_out_4_resp_ready),
    .io_out_4_resp_valid(xbar_io_out_4_resp_valid),
    .io_out_4_resp_bits_rdata(xbar_io_out_4_resp_bits_rdata)
  );
  AXI4UART uart ( // @[src/main/scala/sim/SimMMIO.scala 48:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in_aw_ready(uart_io_in_aw_ready),
    .io_in_aw_valid(uart_io_in_aw_valid),
    .io_in_aw_bits_addr(uart_io_in_aw_bits_addr),
    .io_in_w_ready(uart_io_in_w_ready),
    .io_in_w_valid(uart_io_in_w_valid),
    .io_in_w_bits_data(uart_io_in_w_bits_data),
    .io_in_w_bits_strb(uart_io_in_w_bits_strb),
    .io_in_b_ready(uart_io_in_b_ready),
    .io_in_b_valid(uart_io_in_b_valid),
    .io_in_ar_ready(uart_io_in_ar_ready),
    .io_in_ar_valid(uart_io_in_ar_valid),
    .io_in_ar_bits_addr(uart_io_in_ar_bits_addr),
    .io_in_r_ready(uart_io_in_r_ready),
    .io_in_r_valid(uart_io_in_r_valid),
    .io_in_r_bits_data(uart_io_in_r_bits_data),
    .io_extra_out_valid(uart_io_extra_out_valid),
    .io_extra_out_ch(uart_io_extra_out_ch),
    .io_extra_in_valid(uart_io_extra_in_valid),
    .io_extra_in_ch(uart_io_extra_in_ch)
  );
  AXI4VGA vga ( // @[src/main/scala/sim/SimMMIO.scala 49:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_aw_ready(vga_io_in_fb_aw_ready),
    .io_in_fb_aw_valid(vga_io_in_fb_aw_valid),
    .io_in_fb_aw_bits_addr(vga_io_in_fb_aw_bits_addr),
    .io_in_fb_w_ready(vga_io_in_fb_w_ready),
    .io_in_fb_w_valid(vga_io_in_fb_w_valid),
    .io_in_fb_w_bits_data(vga_io_in_fb_w_bits_data),
    .io_in_fb_w_bits_strb(vga_io_in_fb_w_bits_strb),
    .io_in_fb_b_ready(vga_io_in_fb_b_ready),
    .io_in_fb_b_valid(vga_io_in_fb_b_valid),
    .io_in_fb_ar_ready(vga_io_in_fb_ar_ready),
    .io_in_fb_ar_valid(vga_io_in_fb_ar_valid),
    .io_in_fb_r_ready(vga_io_in_fb_r_ready),
    .io_in_fb_r_valid(vga_io_in_fb_r_valid),
    .io_in_ctrl_aw_ready(vga_io_in_ctrl_aw_ready),
    .io_in_ctrl_aw_valid(vga_io_in_ctrl_aw_valid),
    .io_in_ctrl_w_ready(vga_io_in_ctrl_w_ready),
    .io_in_ctrl_w_valid(vga_io_in_ctrl_w_valid),
    .io_in_ctrl_b_ready(vga_io_in_ctrl_b_ready),
    .io_in_ctrl_b_valid(vga_io_in_ctrl_b_valid),
    .io_in_ctrl_ar_ready(vga_io_in_ctrl_ar_ready),
    .io_in_ctrl_ar_valid(vga_io_in_ctrl_ar_valid),
    .io_in_ctrl_ar_bits_addr(vga_io_in_ctrl_ar_bits_addr),
    .io_in_ctrl_r_ready(vga_io_in_ctrl_r_ready),
    .io_in_ctrl_r_valid(vga_io_in_ctrl_r_valid),
    .io_in_ctrl_r_bits_data(vga_io_in_ctrl_r_bits_data),
    .io_vga_valid(vga_io_vga_valid)
  );
  AXI4Flash flash ( // @[src/main/scala/sim/SimMMIO.scala 50:21]
    .clock(flash_clock),
    .reset(flash_reset),
    .io_in_aw_ready(flash_io_in_aw_ready),
    .io_in_aw_valid(flash_io_in_aw_valid),
    .io_in_w_ready(flash_io_in_w_ready),
    .io_in_w_valid(flash_io_in_w_valid),
    .io_in_b_ready(flash_io_in_b_ready),
    .io_in_b_valid(flash_io_in_b_valid),
    .io_in_ar_ready(flash_io_in_ar_ready),
    .io_in_ar_valid(flash_io_in_ar_valid),
    .io_in_ar_bits_addr(flash_io_in_ar_bits_addr),
    .io_in_r_ready(flash_io_in_r_ready),
    .io_in_r_valid(flash_io_in_r_valid),
    .io_in_r_bits_data(flash_io_in_r_bits_data)
  );
  AXI4DummySD sd ( // @[src/main/scala/sim/SimMMIO.scala 51:18]
    .clock(sd_clock),
    .reset(sd_reset),
    .io_in_aw_ready(sd_io_in_aw_ready),
    .io_in_aw_valid(sd_io_in_aw_valid),
    .io_in_aw_bits_addr(sd_io_in_aw_bits_addr),
    .io_in_w_ready(sd_io_in_w_ready),
    .io_in_w_valid(sd_io_in_w_valid),
    .io_in_w_bits_data(sd_io_in_w_bits_data),
    .io_in_w_bits_strb(sd_io_in_w_bits_strb),
    .io_in_b_ready(sd_io_in_b_ready),
    .io_in_b_valid(sd_io_in_b_valid),
    .io_in_ar_ready(sd_io_in_ar_ready),
    .io_in_ar_valid(sd_io_in_ar_valid),
    .io_in_ar_bits_addr(sd_io_in_ar_bits_addr),
    .io_in_r_ready(sd_io_in_r_ready),
    .io_in_r_valid(sd_io_in_r_valid),
    .io_in_r_bits_data(sd_io_in_r_bits_data)
  );
  SimpleBus2AXI4Converter_3 uart_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(uart_io_in_bridge_clock),
    .reset(uart_io_in_bridge_reset),
    .io_in_req_ready(uart_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(uart_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(uart_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(uart_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(uart_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(uart_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(uart_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(uart_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(uart_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(uart_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(uart_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(uart_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(uart_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(uart_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(uart_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(uart_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(uart_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(uart_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(uart_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(uart_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(uart_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(uart_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(uart_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(uart_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_4 vga_io_in_fb_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_fb_bridge_clock),
    .reset(vga_io_in_fb_bridge_reset),
    .io_in_req_ready(vga_io_in_fb_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_fb_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_fb_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_fb_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(vga_io_in_fb_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(vga_io_in_fb_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(vga_io_in_fb_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_fb_bridge_io_in_resp_valid),
    .io_out_aw_ready(vga_io_in_fb_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_fb_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(vga_io_in_fb_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(vga_io_in_fb_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_fb_bridge_io_out_w_valid),
    .io_out_w_bits_data(vga_io_in_fb_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(vga_io_in_fb_bridge_io_out_w_bits_strb),
    .io_out_b_ready(vga_io_in_fb_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_fb_bridge_io_out_b_valid),
    .io_out_ar_valid(vga_io_in_fb_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_fb_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_fb_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_fb_bridge_io_out_r_valid)
  );
  SimpleBus2AXI4Converter_5 vga_io_in_ctrl_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_ctrl_bridge_clock),
    .reset(vga_io_in_ctrl_bridge_reset),
    .io_in_req_ready(vga_io_in_ctrl_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_ctrl_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_ctrl_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_ctrl_bridge_io_in_req_bits_cmd),
    .io_in_resp_ready(vga_io_in_ctrl_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_ctrl_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(vga_io_in_ctrl_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(vga_io_in_ctrl_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_ctrl_bridge_io_out_aw_valid),
    .io_out_w_ready(vga_io_in_ctrl_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_ctrl_bridge_io_out_w_valid),
    .io_out_b_ready(vga_io_in_ctrl_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_ctrl_bridge_io_out_b_valid),
    .io_out_ar_ready(vga_io_in_ctrl_bridge_io_out_ar_ready),
    .io_out_ar_valid(vga_io_in_ctrl_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_ctrl_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_ctrl_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_ctrl_bridge_io_out_r_valid),
    .io_out_r_bits_data(vga_io_in_ctrl_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_6 flash_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(flash_io_in_bridge_clock),
    .reset(flash_io_in_bridge_reset),
    .io_in_req_ready(flash_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(flash_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(flash_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(flash_io_in_bridge_io_in_req_bits_cmd),
    .io_in_resp_ready(flash_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(flash_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(flash_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(flash_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(flash_io_in_bridge_io_out_aw_valid),
    .io_out_w_ready(flash_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(flash_io_in_bridge_io_out_w_valid),
    .io_out_b_ready(flash_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(flash_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(flash_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(flash_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(flash_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(flash_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(flash_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(flash_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_7 sd_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(sd_io_in_bridge_clock),
    .reset(sd_io_in_bridge_reset),
    .io_in_req_ready(sd_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(sd_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(sd_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(sd_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(sd_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(sd_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(sd_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(sd_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(sd_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(sd_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(sd_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(sd_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(sd_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(sd_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(sd_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(sd_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(sd_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(sd_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(sd_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(sd_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(sd_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(sd_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(sd_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(sd_io_in_bridge_io_out_r_bits_data)
  );
  assign io_rw_req_ready = xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_valid = xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_cmd = xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_rdata = xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_uart_out_valid = uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_out_ch = uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_in_valid = uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_req_valid = io_rw_req_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_addr = io_rw_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_cmd = io_rw_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wmask = io_rw_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wdata = io_rw_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_resp_ready = io_rw_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_out_0_req_ready = uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_valid = uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_bits_rdata = uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_req_ready = vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_valid = vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_req_ready = vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_valid = vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_bits_rdata = vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_req_ready = flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_valid = flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_bits_rdata = flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_req_ready = sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_valid = sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_bits_rdata = sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in_aw_valid = uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_aw_bits_addr = uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_valid = uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_data = uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_strb = uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_b_ready = uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_valid = uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_bits_addr = uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_r_ready = uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_extra_in_ch = io_uart_in_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_aw_valid = vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_aw_bits_addr = vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_valid = vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_data = vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_strb = vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_b_ready = vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_ar_valid = vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_r_ready = vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_aw_valid = vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_w_valid = vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_b_ready = vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_valid = vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_bits_addr = vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_r_ready = vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_clock = clock;
  assign flash_reset = reset;
  assign flash_io_in_aw_valid = flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_w_valid = flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_b_ready = flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_valid = flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_bits_addr = flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_r_ready = flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_clock = clock;
  assign sd_reset = reset;
  assign sd_io_in_aw_valid = sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_aw_bits_addr = sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_valid = sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_data = sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_strb = sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_b_ready = sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_valid = sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_bits_addr = sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_r_ready = sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign uart_io_in_bridge_clock = clock;
  assign uart_io_in_bridge_reset = reset;
  assign uart_io_in_bridge_io_in_req_valid = xbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_addr = xbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_resp_ready = xbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_out_aw_ready = uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_w_ready = uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_b_valid = uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_ar_ready = uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_valid = uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_bits_data = uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign vga_io_in_fb_bridge_clock = clock;
  assign vga_io_in_fb_bridge_reset = reset;
  assign vga_io_in_fb_bridge_io_in_req_valid = xbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_addr = xbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_cmd = xbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wmask = xbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wdata = xbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_resp_ready = xbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_out_aw_ready = vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_w_ready = vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_b_valid = vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_r_valid = vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_bridge_clock = clock;
  assign vga_io_in_ctrl_bridge_reset = reset;
  assign vga_io_in_ctrl_bridge_io_in_req_valid = xbar_io_out_2_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_addr = xbar_io_out_2_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_cmd = xbar_io_out_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_resp_ready = xbar_io_out_2_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_out_aw_ready = vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_w_ready = vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_b_valid = vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_ar_ready = vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_valid = vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_bits_data = vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_io_in_bridge_clock = clock;
  assign flash_io_in_bridge_reset = reset;
  assign flash_io_in_bridge_io_in_req_valid = xbar_io_out_3_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_addr = xbar_io_out_3_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_resp_ready = xbar_io_out_3_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_out_aw_ready = flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_w_ready = flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_b_valid = flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_ar_ready = flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_valid = flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_bits_data = flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_io_in_bridge_clock = clock;
  assign sd_io_in_bridge_reset = reset;
  assign sd_io_in_bridge_io_in_req_valid = xbar_io_out_4_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_addr = xbar_io_out_4_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_4_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_4_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_4_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_resp_ready = xbar_io_out_4_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_out_aw_ready = sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_w_ready = sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_b_valid = sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_ar_ready = sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_valid = sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_bits_data = sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
  end
endmodule
module SimTop(
  input         clock,
  input         reset,
  output [63:0] difftest_exit, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [63:0] difftest_step, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_clean, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_dump, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_begin, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_end, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_level, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_out_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [7:0]  difftest_uart_out_ch, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_in_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [7:0]  difftest_uart_in_ch // @[difftest/src/main/scala/Difftest.scala 496:22]
);
initial assume(reset);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  soc_clock; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_reset; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_b_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [2:0] soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  mem_clock; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_reset; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [2:0] mem_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  memdelay_clock; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_reset; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  mmio_clock; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_reset; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [31:0] mmio_io_rw_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_rw_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  reg [63:0] difftest_timer; // @[difftest/src/main/scala/Difftest.scala 501:24]
  wire [63:0] _difftest_timer_T_1 = difftest_timer + 64'h1; // @[difftest/src/main/scala/Difftest.scala 502:20]
  wire  _T_1 = ~reset; // @[src/main/scala/sim/NutShellSim.scala 57:9]
  wire  line_1903_clock;
  wire  line_1903_reset;
  wire  line_1903_valid;
  reg  line_1903_valid_reg;
  wire  _T_2 = ~(difftest_logCtrl_begin <= difftest_logCtrl_end); // @[src/main/scala/sim/NutShellSim.scala 57:9]
  wire  line_1904_clock;
  wire  line_1904_reset;
  wire  line_1904_valid;
  reg  line_1904_valid_reg;
  wire  difftest_log_enable = difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end; // @[difftest/src/main/scala/Difftest.scala 650:26]
  NutShell soc ( // @[src/main/scala/sim/NutShellSim.scala 34:19]
    .clock(soc_clock),
    .reset(soc_reset),
    .io_mem_aw_ready(soc_io_mem_aw_ready),
    .io_mem_aw_valid(soc_io_mem_aw_valid),
    .io_mem_aw_bits_addr(soc_io_mem_aw_bits_addr),
    .io_mem_w_ready(soc_io_mem_w_ready),
    .io_mem_w_valid(soc_io_mem_w_valid),
    .io_mem_w_bits_data(soc_io_mem_w_bits_data),
    .io_mem_w_bits_strb(soc_io_mem_w_bits_strb),
    .io_mem_w_bits_last(soc_io_mem_w_bits_last),
    .io_mem_b_valid(soc_io_mem_b_valid),
    .io_mem_ar_valid(soc_io_mem_ar_valid),
    .io_mem_ar_bits_addr(soc_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(soc_io_mem_ar_bits_len),
    .io_mem_ar_bits_size(soc_io_mem_ar_bits_size),
    .io_mem_r_valid(soc_io_mem_r_valid),
    .io_mem_r_bits_data(soc_io_mem_r_bits_data),
    .io_mem_r_bits_last(soc_io_mem_r_bits_last),
    .io_mmio_req_ready(soc_io_mmio_req_ready),
    .io_mmio_req_valid(soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr(soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(soc_io_mmio_resp_ready),
    .io_mmio_resp_valid(soc_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(soc_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(soc_io_mmio_resp_bits_rdata)
  );
  AXI4RAM mem ( // @[src/main/scala/sim/NutShellSim.scala 35:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_aw_ready(mem_io_in_aw_ready),
    .io_in_aw_valid(mem_io_in_aw_valid),
    .io_in_aw_bits_addr(mem_io_in_aw_bits_addr),
    .io_in_w_ready(mem_io_in_w_ready),
    .io_in_w_valid(mem_io_in_w_valid),
    .io_in_w_bits_data(mem_io_in_w_bits_data),
    .io_in_w_bits_strb(mem_io_in_w_bits_strb),
    .io_in_w_bits_last(mem_io_in_w_bits_last),
    .io_in_b_valid(mem_io_in_b_valid),
    .io_in_ar_ready(mem_io_in_ar_ready),
    .io_in_ar_valid(mem_io_in_ar_valid),
    .io_in_ar_bits_addr(mem_io_in_ar_bits_addr),
    .io_in_ar_bits_len(mem_io_in_ar_bits_len),
    .io_in_ar_bits_size(mem_io_in_ar_bits_size),
    .io_in_r_valid(mem_io_in_r_valid),
    .io_in_r_bits_data(mem_io_in_r_bits_data),
    .io_in_r_bits_last(mem_io_in_r_bits_last)
  );
  AXI4Delayer memdelay ( // @[src/main/scala/sim/NutShellSim.scala 38:24]
    .clock(memdelay_clock),
    .reset(memdelay_reset),
    .io_in_aw_ready(memdelay_io_in_aw_ready),
    .io_in_aw_valid(memdelay_io_in_aw_valid),
    .io_in_aw_bits_addr(memdelay_io_in_aw_bits_addr),
    .io_in_w_ready(memdelay_io_in_w_ready),
    .io_in_w_valid(memdelay_io_in_w_valid),
    .io_in_w_bits_data(memdelay_io_in_w_bits_data),
    .io_in_w_bits_strb(memdelay_io_in_w_bits_strb),
    .io_in_w_bits_last(memdelay_io_in_w_bits_last),
    .io_in_b_valid(memdelay_io_in_b_valid),
    .io_in_ar_valid(memdelay_io_in_ar_valid),
    .io_in_ar_bits_addr(memdelay_io_in_ar_bits_addr),
    .io_in_ar_bits_len(memdelay_io_in_ar_bits_len),
    .io_in_ar_bits_size(memdelay_io_in_ar_bits_size),
    .io_in_r_valid(memdelay_io_in_r_valid),
    .io_in_r_bits_data(memdelay_io_in_r_bits_data),
    .io_in_r_bits_last(memdelay_io_in_r_bits_last),
    .io_out_aw_ready(memdelay_io_out_aw_ready),
    .io_out_aw_valid(memdelay_io_out_aw_valid),
    .io_out_aw_bits_addr(memdelay_io_out_aw_bits_addr),
    .io_out_w_ready(memdelay_io_out_w_ready),
    .io_out_w_valid(memdelay_io_out_w_valid),
    .io_out_w_bits_data(memdelay_io_out_w_bits_data),
    .io_out_w_bits_strb(memdelay_io_out_w_bits_strb),
    .io_out_w_bits_last(memdelay_io_out_w_bits_last),
    .io_out_b_valid(memdelay_io_out_b_valid),
    .io_out_ar_valid(memdelay_io_out_ar_valid),
    .io_out_ar_bits_addr(memdelay_io_out_ar_bits_addr),
    .io_out_ar_bits_len(memdelay_io_out_ar_bits_len),
    .io_out_ar_bits_size(memdelay_io_out_ar_bits_size),
    .io_out_r_valid(memdelay_io_out_r_valid),
    .io_out_r_bits_data(memdelay_io_out_r_bits_data),
    .io_out_r_bits_last(memdelay_io_out_r_bits_last)
  );
  SimMMIO mmio ( // @[src/main/scala/sim/NutShellSim.scala 39:20]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_rw_req_ready(mmio_io_rw_req_ready),
    .io_rw_req_valid(mmio_io_rw_req_valid),
    .io_rw_req_bits_addr(mmio_io_rw_req_bits_addr),
    .io_rw_req_bits_cmd(mmio_io_rw_req_bits_cmd),
    .io_rw_req_bits_wmask(mmio_io_rw_req_bits_wmask),
    .io_rw_req_bits_wdata(mmio_io_rw_req_bits_wdata),
    .io_rw_resp_ready(mmio_io_rw_resp_ready),
    .io_rw_resp_valid(mmio_io_rw_resp_valid),
    .io_rw_resp_bits_cmd(mmio_io_rw_resp_bits_cmd),
    .io_rw_resp_bits_rdata(mmio_io_rw_resp_bits_rdata),
    .io_uart_out_valid(mmio_io_uart_out_valid),
    .io_uart_out_ch(mmio_io_uart_out_ch),
    .io_uart_in_valid(mmio_io_uart_in_valid),
    .io_uart_in_ch(mmio_io_uart_in_ch)
  );
  GEN_w1_line #(.COVER_INDEX(1903)) line_1903 (
    .clock(line_1903_clock),
    .reset(line_1903_reset),
    .valid(line_1903_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1904)) line_1904 (
    .clock(line_1904_clock),
    .reset(line_1904_reset),
    .valid(line_1904_valid)
  );
  assign line_1903_clock = clock;
  assign line_1903_reset = reset;
  assign line_1903_valid = _T_1 ^ line_1903_valid_reg;
  assign line_1904_clock = clock;
  assign line_1904_reset = reset;
  assign line_1904_valid = _T_2 ^ line_1904_valid_reg;
  assign difftest_exit = 64'h0; // @[difftest/src/main/scala/Difftest.scala 498:19]
  assign difftest_step = 64'h1; // @[difftest/src/main/scala/Difftest.scala 499:19]
  assign difftest_uart_out_valid = mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_out_ch = mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_in_valid = mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign soc_clock = clock;
  assign soc_reset = reset;
  assign soc_io_mem_aw_ready = memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_w_ready = memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_b_valid = memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_valid = memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_data = memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_last = memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mmio_req_ready = mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_valid = mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_cmd = mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_rdata = mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_aw_valid = memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_aw_bits_addr = memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_valid = memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_data = memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_strb = memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_last = memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_valid = memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_addr = memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_len = memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_size = memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_clock = clock;
  assign memdelay_reset = reset;
  assign memdelay_io_in_aw_valid = soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_addr = soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_valid = soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_data = soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_strb = soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_last = soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_valid = soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_addr = soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_len = soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_size = soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_out_aw_ready = mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_w_ready = mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_b_valid = mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_valid = mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_data = mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_last = mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_rw_req_valid = soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_addr = soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_cmd = soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wmask = soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wdata = soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_resp_ready = soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_uart_in_ch = difftest_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/Difftest.scala 501:24]
      difftest_timer <= 64'h0; // @[difftest/src/main/scala/Difftest.scala 501:24]
    end else begin
      difftest_timer <= _difftest_timer_T_1; // @[difftest/src/main/scala/Difftest.scala 502:11]
    end
    line_1903_valid_reg <= _T_1;
    line_1904_valid_reg <= _T_2;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(difftest_logCtrl_begin <= difftest_logCtrl_end)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutShellSim.scala:57 assert(log_begin <= log_end)\n"); // @[src/main/scala/sim/NutShellSim.scala 57:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_timer = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  line_1903_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1904_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (1'h1) begin
      cover(1'h1);
    end
    //
    if (_T_1) begin
      cover(1'h1);
    end
    //
    if (_T_1 & _T_2) begin
      cover(1'h1);
    end
    //
    if (~reset) begin
      assert(difftest_logCtrl_begin <= difftest_logCtrl_end); // @[src/main/scala/sim/NutShellSim.scala 57:9]
    end
  end
endmodule
module array_0(
  input  [8:0]  R0_addr,
  input         R0_en,
  input         R0_clk,
  output [73:0] R0_data,
  input  [8:0]  W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [73:0] W0_data
);
  wire [8:0] array_0_ext_R0_addr;
  wire  array_0_ext_R0_en;
  wire  array_0_ext_R0_clk;
  wire [73:0] array_0_ext_R0_data;
  wire [8:0] array_0_ext_W0_addr;
  wire  array_0_ext_W0_en;
  wire  array_0_ext_W0_clk;
  wire [73:0] array_0_ext_W0_data;
  array_0_ext array_0_ext (
    .R0_addr(array_0_ext_R0_addr),
    .R0_en(array_0_ext_R0_en),
    .R0_clk(array_0_ext_R0_clk),
    .R0_data(array_0_ext_R0_data),
    .W0_addr(array_0_ext_W0_addr),
    .W0_en(array_0_ext_W0_en),
    .W0_clk(array_0_ext_W0_clk),
    .W0_data(array_0_ext_W0_data)
  );
  assign array_0_ext_R0_clk = R0_clk;
  assign array_0_ext_R0_en = R0_en;
  assign array_0_ext_R0_addr = R0_addr;
  assign R0_data = array_0_ext_R0_data[73:0];
  assign array_0_ext_W0_clk = W0_clk;
  assign array_0_ext_W0_en = W0_en;
  assign array_0_ext_W0_addr = W0_addr;
  assign array_0_ext_W0_data = W0_data;
endmodule
