module IntXbar(
  input   clock,
  input   reset
);
endmodule
module InterruptBusWrapper(
  input   auto_clock_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_clock_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output  reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  int_bus_clock; // @[src/main/scala/subsystem/InterruptBus.scala 14:27]
  wire  int_bus_reset; // @[src/main/scala/subsystem/InterruptBus.scala 14:27]
  IntXbar int_bus ( // @[src/main/scala/subsystem/InterruptBus.scala 14:27]
    .clock(int_bus_clock),
    .reset(int_bus_reset)
  );
  assign clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign int_bus_clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign int_bus_reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module SimpleClockGroupSource(
  input   clock,
  input   reset,
  output  auto_out_member_subsystem_sbus_5_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_5_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_4_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_4_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_3_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_3_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_2_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_2_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_sbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_member_subsystem_sbus_5_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_5_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
  assign auto_out_member_subsystem_sbus_4_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_4_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
  assign auto_out_member_subsystem_sbus_3_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_3_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
  assign auto_out_member_subsystem_sbus_2_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_2_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
  assign auto_out_member_subsystem_sbus_1_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_1_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
  assign auto_out_member_subsystem_sbus_0_clock = clock; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:17]
  assign auto_out_member_subsystem_sbus_0_reset = reset; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/prci/ClockGroup.scala 75:35]
endmodule
module ClockGroupAggregator(
  input   auto_in_member_subsystem_sbus_5_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_5_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_4_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_4_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_3_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_3_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_2_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_2_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_3_member_subsystem_l2_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_3_member_subsystem_l2_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_3_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_3_member_subsystem_l2_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_2_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_2_member_subsystem_fbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_cbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_cbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_cbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_sbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_sbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_3_member_subsystem_l2_1_clock = auto_in_member_subsystem_sbus_5_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_3_member_subsystem_l2_1_reset = auto_in_member_subsystem_sbus_5_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_3_member_subsystem_l2_0_clock = auto_in_member_subsystem_sbus_4_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_3_member_subsystem_l2_0_reset = auto_in_member_subsystem_sbus_4_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_2_member_subsystem_fbus_0_clock = auto_in_member_subsystem_sbus_3_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_2_member_subsystem_fbus_0_reset = auto_in_member_subsystem_sbus_3_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_cbus_1_clock = auto_in_member_subsystem_sbus_2_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_cbus_1_reset = auto_in_member_subsystem_sbus_2_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_cbus_0_clock = auto_in_member_subsystem_sbus_1_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_cbus_0_reset = auto_in_member_subsystem_sbus_1_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_sbus_0_clock = auto_in_member_subsystem_sbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_sbus_0_reset = auto_in_member_subsystem_sbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup(
  input   auto_in_member_subsystem_sbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_sbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_sbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_sbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_2_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_2_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_2_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_2_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus(
  input   clock,
  input   reset
);
endmodule
module TLXbar(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_1_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_1_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_1_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_1_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_1_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_1_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_1_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_1_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_1_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_1_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_1_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_1_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_1_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_1_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_1_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_1_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_1_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_1_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_1_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_1_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_1_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_1_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_1_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_0_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_0_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_0_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_0_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_0_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_0_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_0_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_0_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_0_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_0_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_0_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_0_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_0_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_0_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_0_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_0_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] beatsLeft; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
  wire  idle = beatsLeft == 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 61:28]
  wire [1:0] readys_valid = {auto_out_1_d_valid,auto_out_0_d_valid}; // @[src/main/scala/tilelink/Arbiter.scala 68:51]
  reg [1:0] readys_mask; // @[src/main/scala/tilelink/Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[src/main/scala/tilelink/Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[src/main/scala/tilelink/Arbiter.scala 24:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,auto_out_1_d_valid,auto_out_0_d_valid}; // @[src/main/scala/tilelink/Arbiter.scala 24:21]
  wire [3:0] _GEN_8 = {{1'd0}, readys_filter[3:1]}; // @[src/main/scala/util/package.scala 254:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_8; // @[src/main/scala/util/package.scala 254:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[src/main/scala/tilelink/Arbiter.scala 25:66]
  wire [3:0] _GEN_9 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[src/main/scala/tilelink/Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_9 | _readys_unready_T_4; // @[src/main/scala/tilelink/Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[src/main/scala/tilelink/Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[src/main/scala/tilelink/Arbiter.scala 26:18]
  wire  readys_0 = readys_readys[0]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  winner_0 = readys_0 & auto_out_0_d_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  reg  state_0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  muxState_0 = idle ? winner_0 : state_0; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire [1:0] _in_0_d_bits_T_12 = muxState_0 ? auto_out_0_d_bits_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  readys_1 = readys_readys[1]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  winner_1 = readys_1 & auto_out_1_d_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  reg  state_1; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  muxState_1 = idle ? winner_1 : state_1; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire [1:0] _in_0_d_bits_T_13 = muxState_1 ? auto_out_1_d_bits_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [32:0] _requestAIO_T_1 = {1'b0,$signed(auto_in_a_bits_address)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [32:0] _requestAIO_T_3 = $signed(_requestAIO_T_1) & 33'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  requestAIO_0_0 = $signed(_requestAIO_T_3) == 33'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire [31:0] _requestAIO_T_5 = auto_in_a_bits_address ^ 32'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [32:0] _requestAIO_T_6 = {1'b0,$signed(_requestAIO_T_5)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [32:0] _requestAIO_T_8 = $signed(_requestAIO_T_6) & 33'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  requestAIO_0_1 = $signed(_requestAIO_T_8) == 33'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire [11:0] _beatsDO_decode_T_1 = 12'h1f << auto_out_0_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beatsDO_decode_T_3 = ~_beatsDO_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beatsDO_decode = _beatsDO_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire [11:0] _beatsDO_decode_T_5 = 12'h1f << auto_out_1_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beatsDO_decode_T_7 = ~_beatsDO_decode_T_5[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beatsDO_decode_1 = _beatsDO_decode_T_7[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  beatsDO_opdata_1 = auto_out_1_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  wire [1:0] beatsDO_1 = beatsDO_opdata_1 ? beatsDO_decode_1 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire  latch = idle & auto_in_d_ready; // @[src/main/scala/tilelink/Arbiter.scala 62:24]
  wire  _readys_T_3 = ~reset; // @[src/main/scala/tilelink/Arbiter.scala 22:12]
  wire  line_0_clock;
  wire  line_0_reset;
  wire  line_0_valid;
  reg  line_0_valid_reg;
  wire  _readys_T_6 = latch & |readys_valid; // @[src/main/scala/tilelink/Arbiter.scala 27:18]
  wire  line_1_clock;
  wire  line_1_reset;
  wire  line_1_valid;
  reg  line_1_valid_reg;
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[src/main/scala/tilelink/Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[src/main/scala/util/package.scala 245:43]
  wire  _prefixOR_T = winner_0 | winner_1; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  line_2_clock;
  wire  line_2_reset;
  wire  line_2_valid;
  reg  line_2_valid_reg;
  wire  _T_9 = ~(~winner_0 | ~winner_1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
  wire  line_3_clock;
  wire  line_3_reset;
  wire  line_3_valid;
  reg  line_3_valid_reg;
  wire  _T_10 = auto_out_0_d_valid | auto_out_1_d_valid; // @[src/main/scala/tilelink/Arbiter.scala 79:31]
  wire  line_4_clock;
  wire  line_4_reset;
  wire  line_4_valid;
  reg  line_4_valid_reg;
  wire  _T_16 = ~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
  wire  line_5_clock;
  wire  line_5_reset;
  wire  line_5_valid;
  reg  line_5_valid_reg;
  wire [1:0] maskedBeats_0 = winner_0 ? beatsDO_decode : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] maskedBeats_1 = winner_1 ? beatsDO_1 : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] initBeats = maskedBeats_0 | maskedBeats_1; // @[src/main/scala/tilelink/Arbiter.scala 84:44]
  wire  _in_0_d_valid_T_3 = state_0 & auto_out_0_d_valid | state_1 & auto_out_1_d_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  in_0_d_valid = idle ? _T_10 : _in_0_d_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  wire  _beatsLeft_T = auto_in_d_ready & in_0_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_10 = {{1'd0}, _beatsLeft_T}; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire [1:0] _beatsLeft_T_2 = beatsLeft - _GEN_10; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire [63:0] _in_0_d_bits_T_3 = muxState_0 ? auto_out_0_d_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _in_0_d_bits_T_4 = muxState_1 ? auto_out_1_d_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] out_0_d_bits_sink = {{1'd0}, auto_out_0_d_bits_sink}; // @[src/main/scala/tilelink/Xbar.scala 213:19 248:28]
  wire [1:0] _in_0_d_bits_T_9 = muxState_0 ? out_0_d_bits_sink : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _in_0_d_bits_T_10 = muxState_1 ? auto_out_1_d_bits_sink : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _in_0_d_bits_T_15 = muxState_0 ? auto_out_0_d_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _in_0_d_bits_T_16 = muxState_1 ? auto_out_1_d_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _in_0_d_bits_T_18 = muxState_0 ? auto_out_0_d_bits_param : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _in_0_d_bits_T_19 = muxState_1 ? auto_out_1_d_bits_param : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _in_0_d_bits_T_21 = muxState_0 ? auto_out_0_d_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _in_0_d_bits_T_22 = muxState_1 ? auto_out_1_d_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  GEN_w1_line #(.COVER_INDEX(0)) line_0 (
    .clock(line_0_clock),
    .reset(line_0_reset),
    .valid(line_0_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1)) line_1 (
    .clock(line_1_clock),
    .reset(line_1_reset),
    .valid(line_1_valid)
  );
  GEN_w1_line #(.COVER_INDEX(2)) line_2 (
    .clock(line_2_clock),
    .reset(line_2_reset),
    .valid(line_2_valid)
  );
  GEN_w1_line #(.COVER_INDEX(3)) line_3 (
    .clock(line_3_clock),
    .reset(line_3_reset),
    .valid(line_3_valid)
  );
  GEN_w1_line #(.COVER_INDEX(4)) line_4 (
    .clock(line_4_clock),
    .reset(line_4_reset),
    .valid(line_4_valid)
  );
  GEN_w1_line #(.COVER_INDEX(5)) line_5 (
    .clock(line_5_clock),
    .reset(line_5_reset),
    .valid(line_5_valid)
  );
  assign line_0_clock = clock;
  assign line_0_reset = reset;
  assign line_0_valid = _readys_T_3 ^ line_0_valid_reg;
  assign line_1_clock = clock;
  assign line_1_reset = reset;
  assign line_1_valid = _readys_T_6 ^ line_1_valid_reg;
  assign line_2_clock = clock;
  assign line_2_reset = reset;
  assign line_2_valid = _readys_T_3 ^ line_2_valid_reg;
  assign line_3_clock = clock;
  assign line_3_reset = reset;
  assign line_3_valid = _T_9 ^ line_3_valid_reg;
  assign line_4_clock = clock;
  assign line_4_reset = reset;
  assign line_4_valid = _readys_T_3 ^ line_4_valid_reg;
  assign line_5_clock = clock;
  assign line_5_reset = reset;
  assign line_5_valid = _T_16 ^ line_5_valid_reg;
  assign auto_in_a_ready = requestAIO_0_0 & auto_out_0_a_ready | requestAIO_0_1 & auto_out_1_a_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_b_valid = auto_out_1_b_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_b_bits_param = auto_out_1_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_1_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_1_c_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_valid = idle ? _T_10 : _in_0_d_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  assign auto_in_d_bits_opcode = _in_0_d_bits_T_21 | _in_0_d_bits_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_param = _in_0_d_bits_T_18 | _in_0_d_bits_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_size = _in_0_d_bits_T_15 | _in_0_d_bits_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_source = _in_0_d_bits_T_12 | _in_0_d_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_sink = _in_0_d_bits_T_9 | _in_0_d_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_denied = muxState_0 & auto_out_0_d_bits_denied | muxState_1 & auto_out_1_d_bits_denied; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_data = _in_0_d_bits_T_3 | _in_0_d_bits_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_corrupt = muxState_0 & auto_out_0_d_bits_corrupt | muxState_1 & auto_out_1_d_bits_corrupt; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_1_a_valid = auto_in_a_valid & requestAIO_0_1; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_1_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_1_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_c_valid = auto_in_c_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_1_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/tilelink/Xbar.scala 184:55]
  assign auto_out_1_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_d_ready = auto_in_d_ready & allowed_1; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign auto_out_1_e_valid = auto_in_e_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_1_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_out_0_a_valid = auto_in_a_valid & requestAIO_0_0; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_0_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_0_a_bits_address = auto_in_a_bits_address[28:0]; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Xbar.scala 218:41]
  assign auto_out_0_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_d_ready = auto_in_d_ready & allowed_0; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 60:30]
      beatsLeft <= 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
    end else if (latch) begin // @[src/main/scala/tilelink/Arbiter.scala 85:23]
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= _beatsLeft_T_2;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[src/main/scala/tilelink/Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin // @[src/main/scala/tilelink/Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_3; // @[src/main/scala/tilelink/Arbiter.scala 28:12]
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_0 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_0 <= winner_0;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1 <= winner_1;
    end
    line_0_valid_reg <= _readys_T_3;
    line_1_valid_reg <= _readys_T_6;
    line_2_valid_reg <= _readys_T_3;
    line_3_valid_reg <= _T_9;
    line_4_valid_reg <= _readys_T_3;
    line_5_valid_reg <= _T_16;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~winner_0 | ~winner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  readys_mask = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_0_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_2_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_3_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_4_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_5_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/tilelink/Arbiter.scala 22:12]
    end
    //
    if (_readys_T_3) begin
      assert(~winner_0 | ~winner_1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
    end
    //
    if (_readys_T_3) begin
      assert(~(auto_out_0_d_valid | auto_out_1_d_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
    end
  end
endmodule
module TLFIFOFixer(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _a_first_T = auto_out_a_ready & auto_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _a_first_beats1_decode_T_1 = 12'h1f << auto_in_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  reg [1:0] a_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] a_first_counter1 = a_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_6_clock;
  wire  line_6_reset;
  wire  line_6_valid;
  reg  line_6_valid_reg;
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _d_first_beats1_decode_T_1 = 12'h1f << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  reg [1:0] d_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] d_first_counter1 = d_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  d_first_first = d_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_7_clock;
  wire  line_7_reset;
  wire  line_7_valid;
  reg  line_7_valid_reg;
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[src/main/scala/tilelink/FIFOFixer.scala 69:42]
  wire  _T_1 = a_first & _a_first_T; // @[src/main/scala/tilelink/FIFOFixer.scala 74:21]
  wire  line_8_clock;
  wire  line_8_reset;
  wire  line_8_valid;
  reg  line_8_valid_reg;
  wire  line_9_clock;
  wire  line_9_reset;
  wire  line_9_valid;
  reg  line_9_valid_reg;
  wire  line_10_clock;
  wire  line_10_reset;
  wire  line_10_valid;
  reg  line_10_valid_reg;
  wire  line_11_clock;
  wire  line_11_reset;
  wire  line_11_valid;
  reg  line_11_valid_reg;
  wire  _T_3 = d_first & _d_first_T; // @[src/main/scala/tilelink/FIFOFixer.scala 75:21]
  wire  line_12_clock;
  wire  line_12_reset;
  wire  line_12_valid;
  reg  line_12_valid_reg;
  wire  line_13_clock;
  wire  line_13_reset;
  wire  line_13_valid;
  reg  line_13_valid_reg;
  wire  line_14_clock;
  wire  line_14_reset;
  wire  line_14_valid;
  reg  line_14_valid_reg;
  wire  line_15_clock;
  wire  line_15_reset;
  wire  line_15_valid;
  reg  line_15_valid_reg;
  wire  line_16_clock;
  wire  line_16_reset;
  wire  line_16_valid;
  reg  line_16_valid_reg;
  GEN_w1_line #(.COVER_INDEX(6)) line_6 (
    .clock(line_6_clock),
    .reset(line_6_reset),
    .valid(line_6_valid)
  );
  GEN_w1_line #(.COVER_INDEX(7)) line_7 (
    .clock(line_7_clock),
    .reset(line_7_reset),
    .valid(line_7_valid)
  );
  GEN_w1_line #(.COVER_INDEX(8)) line_8 (
    .clock(line_8_clock),
    .reset(line_8_reset),
    .valid(line_8_valid)
  );
  GEN_w1_line #(.COVER_INDEX(9)) line_9 (
    .clock(line_9_clock),
    .reset(line_9_reset),
    .valid(line_9_valid)
  );
  GEN_w1_line #(.COVER_INDEX(10)) line_10 (
    .clock(line_10_clock),
    .reset(line_10_reset),
    .valid(line_10_valid)
  );
  GEN_w1_line #(.COVER_INDEX(11)) line_11 (
    .clock(line_11_clock),
    .reset(line_11_reset),
    .valid(line_11_valid)
  );
  GEN_w1_line #(.COVER_INDEX(12)) line_12 (
    .clock(line_12_clock),
    .reset(line_12_reset),
    .valid(line_12_valid)
  );
  GEN_w1_line #(.COVER_INDEX(13)) line_13 (
    .clock(line_13_clock),
    .reset(line_13_reset),
    .valid(line_13_valid)
  );
  GEN_w1_line #(.COVER_INDEX(14)) line_14 (
    .clock(line_14_clock),
    .reset(line_14_reset),
    .valid(line_14_valid)
  );
  GEN_w1_line #(.COVER_INDEX(15)) line_15 (
    .clock(line_15_clock),
    .reset(line_15_reset),
    .valid(line_15_valid)
  );
  GEN_w1_line #(.COVER_INDEX(16)) line_16 (
    .clock(line_16_clock),
    .reset(line_16_reset),
    .valid(line_16_valid)
  );
  assign line_6_clock = clock;
  assign line_6_reset = reset;
  assign line_6_valid = _a_first_T ^ line_6_valid_reg;
  assign line_7_clock = clock;
  assign line_7_reset = reset;
  assign line_7_valid = _d_first_T ^ line_7_valid_reg;
  assign line_8_clock = clock;
  assign line_8_reset = reset;
  assign line_8_valid = _T_1 ^ line_8_valid_reg;
  assign line_9_clock = clock;
  assign line_9_reset = reset;
  assign line_9_valid = 2'h0 == auto_in_a_bits_source ^ line_9_valid_reg;
  assign line_10_clock = clock;
  assign line_10_reset = reset;
  assign line_10_valid = 2'h1 == auto_in_a_bits_source ^ line_10_valid_reg;
  assign line_11_clock = clock;
  assign line_11_reset = reset;
  assign line_11_valid = 2'h2 == auto_in_a_bits_source ^ line_11_valid_reg;
  assign line_12_clock = clock;
  assign line_12_reset = reset;
  assign line_12_valid = _T_3 ^ line_12_valid_reg;
  assign line_13_clock = clock;
  assign line_13_reset = reset;
  assign line_13_valid = 2'h0 == auto_out_d_bits_source ^ line_13_valid_reg;
  assign line_14_clock = clock;
  assign line_14_reset = reset;
  assign line_14_valid = 2'h1 == auto_out_d_bits_source ^ line_14_valid_reg;
  assign line_15_clock = clock;
  assign line_15_reset = reset;
  assign line_15_valid = 2'h2 == auto_out_d_bits_source ^ line_15_valid_reg;
  assign line_16_clock = clock;
  assign line_16_reset = reset;
  assign line_16_valid = _T_3 ^ line_16_valid_reg;
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 90:33]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 89:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      a_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_a_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (a_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (a_first_beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 2'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    line_6_valid_reg <= _a_first_T;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      d_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_d_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (d_first_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (d_first_beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 2'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    line_7_valid_reg <= _d_first_T;
    line_8_valid_reg <= _T_1;
    line_9_valid_reg <= 2'h0 == auto_in_a_bits_source;
    line_10_valid_reg <= 2'h1 == auto_in_a_bits_source;
    line_11_valid_reg <= 2'h2 == auto_in_a_bits_source;
    line_12_valid_reg <= _T_3;
    line_13_valid_reg <= 2'h0 == auto_out_d_bits_source;
    line_14_valid_reg <= 2'h1 == auto_out_d_bits_source;
    line_15_valid_reg <= 2'h2 == auto_out_d_bits_source;
    line_16_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_6_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  d_first_counter = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  line_7_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_8_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_9_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_10_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_11_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_12_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_13_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_14_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_15_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_16_valid_reg = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLInterconnectCoupler(
  input         clock,
  input         reset,
  output        auto_widget_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_widget_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_widget_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_bus_xing_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_bus_xing_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_bus_xing_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_bus_xing_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_bus_xing_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_bus_xing_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [28:0] widget_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [28:0] widget_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_out_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
  );
  assign auto_widget_in_a_ready = widget_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_valid = widget_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_param = widget_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_sink = widget_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bus_xing_out_a_valid = widget_auto_out_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_size = widget_auto_out_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_source = widget_auto_out_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_address = widget_auto_out_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_mask = widget_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_d_ready = widget_auto_out_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_d_ready = auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_out_a_ready = auto_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_valid = auto_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_opcode = auto_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_param = auto_bus_xing_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_size = auto_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_source = auto_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_sink = auto_bus_xing_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_denied = auto_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_data = auto_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_corrupt = auto_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
endmodule
module TLWidthWidget_1(
  input   clock,
  input   reset
);
endmodule
module TLInterconnectCoupler_1(
  input   clock,
  input   reset
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget_1 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset)
  );
  assign widget_clock = clock;
  assign widget_reset = reset;
endmodule
module TLWidthWidget_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLInterconnectCoupler_2(
  input         clock,
  input         reset,
  output        auto_widget_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_widget_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_widget_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_widget_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_widget_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_widget_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_widget_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_widget_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_widget_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_widget_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_widget_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_widget_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_widget_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_widget_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_b_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_b_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_b_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_b_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_c_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_c_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_c_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_c_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_c_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_e_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_e_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_out_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_b_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_b_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_b_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_b_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_c_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_c_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_c_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_c_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_c_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_e_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_e_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget_2 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_b_ready(widget_auto_in_b_ready),
    .auto_in_b_valid(widget_auto_in_b_valid),
    .auto_in_b_bits_param(widget_auto_in_b_bits_param),
    .auto_in_b_bits_address(widget_auto_in_b_bits_address),
    .auto_in_c_ready(widget_auto_in_c_ready),
    .auto_in_c_valid(widget_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_auto_in_c_bits_address),
    .auto_in_c_bits_data(widget_auto_in_c_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_in_e_valid(widget_auto_in_e_valid),
    .auto_in_e_bits_sink(widget_auto_in_e_bits_sink),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_b_ready(widget_auto_out_b_ready),
    .auto_out_b_valid(widget_auto_out_b_valid),
    .auto_out_b_bits_param(widget_auto_out_b_bits_param),
    .auto_out_b_bits_address(widget_auto_out_b_bits_address),
    .auto_out_c_ready(widget_auto_out_c_ready),
    .auto_out_c_valid(widget_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_auto_out_c_bits_address),
    .auto_out_c_bits_data(widget_auto_out_c_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt),
    .auto_out_e_valid(widget_auto_out_e_valid),
    .auto_out_e_bits_sink(widget_auto_out_e_bits_sink)
  );
  assign auto_widget_in_a_ready = widget_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_b_valid = widget_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_b_bits_param = widget_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_b_bits_address = widget_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_c_ready = widget_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_valid = widget_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_param = widget_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_sink = widget_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_out_a_valid = widget_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_param = widget_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_size = widget_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_source = widget_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_address = widget_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_mask = widget_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_a_bits_data = widget_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_b_ready = widget_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_valid = widget_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_opcode = widget_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_param = widget_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_size = widget_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_source = widget_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_address = widget_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_c_bits_data = widget_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_d_ready = widget_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_e_valid = widget_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_widget_out_e_bits_sink = widget_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_opcode = auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_param = auto_widget_in_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_data = auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_b_ready = auto_widget_in_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_valid = auto_widget_in_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_opcode = auto_widget_in_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_param = auto_widget_in_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_size = auto_widget_in_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_source = auto_widget_in_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_address = auto_widget_in_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_c_bits_data = auto_widget_in_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_d_ready = auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_e_valid = auto_widget_in_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_e_bits_sink = auto_widget_in_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_out_a_ready = auto_widget_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_b_valid = auto_widget_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_b_bits_param = auto_widget_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_b_bits_address = auto_widget_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_c_ready = auto_widget_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_valid = auto_widget_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_opcode = auto_widget_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_param = auto_widget_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_size = auto_widget_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_source = auto_widget_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_sink = auto_widget_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_denied = auto_widget_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_data = auto_widget_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_corrupt = auto_widget_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
endmodule
module TLInterconnectCoupler_3(
  input         clock,
  input         reset,
  output        auto_tl_master_clock_xing_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tl_master_clock_xing_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_tl_master_clock_xing_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_master_clock_xing_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_master_clock_xing_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tl_master_clock_xing_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_master_clock_xing_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_master_clock_xing_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_tl_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tl_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_tl_master_clock_xing_in_a_ready = auto_tl_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_b_valid = auto_tl_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_b_bits_param = auto_tl_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_b_bits_address = auto_tl_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_c_ready = auto_tl_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_valid = auto_tl_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_opcode = auto_tl_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_param = auto_tl_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_size = auto_tl_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_source = auto_tl_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_sink = auto_tl_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_denied = auto_tl_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_data = auto_tl_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_master_clock_xing_in_d_bits_corrupt = auto_tl_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_out_a_valid = auto_tl_master_clock_xing_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_opcode = auto_tl_master_clock_xing_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_param = auto_tl_master_clock_xing_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_size = auto_tl_master_clock_xing_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_source = auto_tl_master_clock_xing_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_address = auto_tl_master_clock_xing_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_mask = auto_tl_master_clock_xing_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_data = auto_tl_master_clock_xing_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_b_ready = auto_tl_master_clock_xing_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_valid = auto_tl_master_clock_xing_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_opcode = auto_tl_master_clock_xing_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_param = auto_tl_master_clock_xing_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_size = auto_tl_master_clock_xing_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_source = auto_tl_master_clock_xing_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_address = auto_tl_master_clock_xing_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_c_bits_data = auto_tl_master_clock_xing_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_d_ready = auto_tl_master_clock_xing_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_e_valid = auto_tl_master_clock_xing_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_e_bits_sink = auto_tl_master_clock_xing_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module SystemBus(
  output        auto_coupler_from_tile_tl_master_clock_xing_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_from_tile_tl_master_clock_xing_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_from_tile_tl_master_clock_xing_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_from_tile_tl_master_clock_xing_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_from_tile_tl_master_clock_xing_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_from_tile_tl_master_clock_xing_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_from_tile_tl_master_clock_xing_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_from_tile_tl_master_clock_xing_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_from_tile_tl_master_clock_xing_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_sbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_sbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_2_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_2_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_1_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_1_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_0_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_0_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  system_bus_xbar_clock; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_reset; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_a_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_a_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_in_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_in_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_a_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_b_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_b_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_b_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_in_b_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_c_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_c_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_c_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_c_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_c_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_c_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_in_c_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_c_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_in_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_in_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_in_e_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_in_e_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_a_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_a_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_out_1_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_out_1_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_1_a_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_b_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_b_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_b_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_out_1_b_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_c_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_c_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_c_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_c_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_c_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_c_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [31:0] system_bus_xbar_auto_out_1_c_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_1_c_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_1_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_1_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_1_e_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_1_e_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_0_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [28:0] system_bus_xbar_auto_out_0_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [7:0] system_bus_xbar_auto_out_0_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_0_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [2:0] system_bus_xbar_auto_out_0_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [1:0] system_bus_xbar_auto_out_0_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire [63:0] system_bus_xbar_auto_out_0_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  system_bus_xbar_auto_out_0_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 40:43]
  wire  fixer_clock; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_reset; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_a_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_a_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_a_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_in_a_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_b_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_b_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_b_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_in_b_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_c_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_c_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_c_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_c_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_c_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_c_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_in_c_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_in_c_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_d_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_d_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_d_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_d_bits_sink; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_in_d_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_e_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_in_e_bits_sink; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_a_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_a_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_a_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_out_a_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_b_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_b_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_b_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_out_b_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_c_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_c_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_c_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_c_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_c_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_c_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_out_c_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_out_c_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_d_bits_param; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_d_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_d_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_d_bits_sink; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_bits_denied; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_out_d_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_e_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [1:0] fixer_auto_out_e_bits_sink; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  coupler_to_bus_named_subsystem_cbus_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [28:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [28:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_bus_named_subsystem_fbus_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_bus_named_subsystem_fbus_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_in_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_in_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_l2_auto_widget_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bus_named_subsystem_l2_auto_widget_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_master_clock_xing_in_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_master_clock_xing_in_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_from_tile_auto_tl_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_from_tile_auto_tl_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_from_tile_auto_tl_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_from_tile_auto_tl_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_from_tile_auto_tl_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_from_tile_auto_tl_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  ClockGroupAggregator subsystem_sbus_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_sbus_5_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock),
    .auto_in_member_subsystem_sbus_5_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset),
    .auto_in_member_subsystem_sbus_4_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock),
    .auto_in_member_subsystem_sbus_4_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset),
    .auto_in_member_subsystem_sbus_3_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock),
    .auto_in_member_subsystem_sbus_3_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset),
    .auto_in_member_subsystem_sbus_2_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock),
    .auto_in_member_subsystem_sbus_2_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset),
    .auto_in_member_subsystem_sbus_1_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock),
    .auto_in_member_subsystem_sbus_1_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset),
    .auto_in_member_subsystem_sbus_0_clock(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock),
    .auto_in_member_subsystem_sbus_0_reset(subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset),
    .auto_out_3_member_subsystem_l2_1_clock(subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock),
    .auto_out_3_member_subsystem_l2_1_reset(subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset),
    .auto_out_3_member_subsystem_l2_0_clock(subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock),
    .auto_out_3_member_subsystem_l2_0_reset(subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset),
    .auto_out_2_member_subsystem_fbus_0_clock(subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock),
    .auto_out_2_member_subsystem_fbus_0_reset(subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset),
    .auto_out_1_member_subsystem_cbus_1_clock(subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock),
    .auto_out_1_member_subsystem_cbus_1_reset(subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset),
    .auto_out_1_member_subsystem_cbus_0_clock(subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock),
    .auto_out_1_member_subsystem_cbus_0_reset(subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset),
    .auto_out_0_member_subsystem_sbus_0_clock(subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock),
    .auto_out_0_member_subsystem_sbus_0_reset(subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset)
  );
  ClockGroup clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_sbus_0_clock(clockGroup_auto_in_member_subsystem_sbus_0_clock),
    .auto_in_member_subsystem_sbus_0_reset(clockGroup_auto_in_member_subsystem_sbus_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_2_clock(fixedClockNode_auto_out_2_clock),
    .auto_out_2_reset(fixedClockNode_auto_out_2_reset),
    .auto_out_1_clock(fixedClockNode_auto_out_1_clock),
    .auto_out_1_reset(fixedClockNode_auto_out_1_reset),
    .auto_out_0_clock(fixedClockNode_auto_out_0_clock),
    .auto_out_0_reset(fixedClockNode_auto_out_0_reset)
  );
  BundleBridgeNexus broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLXbar system_bus_xbar ( // @[src/main/scala/subsystem/SystemBus.scala 40:43]
    .clock(system_bus_xbar_clock),
    .reset(system_bus_xbar_reset),
    .auto_in_a_ready(system_bus_xbar_auto_in_a_ready),
    .auto_in_a_valid(system_bus_xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(system_bus_xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(system_bus_xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(system_bus_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(system_bus_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(system_bus_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(system_bus_xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(system_bus_xbar_auto_in_a_bits_data),
    .auto_in_b_ready(system_bus_xbar_auto_in_b_ready),
    .auto_in_b_valid(system_bus_xbar_auto_in_b_valid),
    .auto_in_b_bits_param(system_bus_xbar_auto_in_b_bits_param),
    .auto_in_b_bits_address(system_bus_xbar_auto_in_b_bits_address),
    .auto_in_c_ready(system_bus_xbar_auto_in_c_ready),
    .auto_in_c_valid(system_bus_xbar_auto_in_c_valid),
    .auto_in_c_bits_opcode(system_bus_xbar_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(system_bus_xbar_auto_in_c_bits_param),
    .auto_in_c_bits_size(system_bus_xbar_auto_in_c_bits_size),
    .auto_in_c_bits_source(system_bus_xbar_auto_in_c_bits_source),
    .auto_in_c_bits_address(system_bus_xbar_auto_in_c_bits_address),
    .auto_in_c_bits_data(system_bus_xbar_auto_in_c_bits_data),
    .auto_in_d_ready(system_bus_xbar_auto_in_d_ready),
    .auto_in_d_valid(system_bus_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(system_bus_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(system_bus_xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(system_bus_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(system_bus_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(system_bus_xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(system_bus_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(system_bus_xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(system_bus_xbar_auto_in_d_bits_corrupt),
    .auto_in_e_valid(system_bus_xbar_auto_in_e_valid),
    .auto_in_e_bits_sink(system_bus_xbar_auto_in_e_bits_sink),
    .auto_out_1_a_ready(system_bus_xbar_auto_out_1_a_ready),
    .auto_out_1_a_valid(system_bus_xbar_auto_out_1_a_valid),
    .auto_out_1_a_bits_opcode(system_bus_xbar_auto_out_1_a_bits_opcode),
    .auto_out_1_a_bits_param(system_bus_xbar_auto_out_1_a_bits_param),
    .auto_out_1_a_bits_size(system_bus_xbar_auto_out_1_a_bits_size),
    .auto_out_1_a_bits_source(system_bus_xbar_auto_out_1_a_bits_source),
    .auto_out_1_a_bits_address(system_bus_xbar_auto_out_1_a_bits_address),
    .auto_out_1_a_bits_mask(system_bus_xbar_auto_out_1_a_bits_mask),
    .auto_out_1_a_bits_data(system_bus_xbar_auto_out_1_a_bits_data),
    .auto_out_1_b_ready(system_bus_xbar_auto_out_1_b_ready),
    .auto_out_1_b_valid(system_bus_xbar_auto_out_1_b_valid),
    .auto_out_1_b_bits_param(system_bus_xbar_auto_out_1_b_bits_param),
    .auto_out_1_b_bits_address(system_bus_xbar_auto_out_1_b_bits_address),
    .auto_out_1_c_ready(system_bus_xbar_auto_out_1_c_ready),
    .auto_out_1_c_valid(system_bus_xbar_auto_out_1_c_valid),
    .auto_out_1_c_bits_opcode(system_bus_xbar_auto_out_1_c_bits_opcode),
    .auto_out_1_c_bits_param(system_bus_xbar_auto_out_1_c_bits_param),
    .auto_out_1_c_bits_size(system_bus_xbar_auto_out_1_c_bits_size),
    .auto_out_1_c_bits_source(system_bus_xbar_auto_out_1_c_bits_source),
    .auto_out_1_c_bits_address(system_bus_xbar_auto_out_1_c_bits_address),
    .auto_out_1_c_bits_data(system_bus_xbar_auto_out_1_c_bits_data),
    .auto_out_1_d_ready(system_bus_xbar_auto_out_1_d_ready),
    .auto_out_1_d_valid(system_bus_xbar_auto_out_1_d_valid),
    .auto_out_1_d_bits_opcode(system_bus_xbar_auto_out_1_d_bits_opcode),
    .auto_out_1_d_bits_param(system_bus_xbar_auto_out_1_d_bits_param),
    .auto_out_1_d_bits_size(system_bus_xbar_auto_out_1_d_bits_size),
    .auto_out_1_d_bits_source(system_bus_xbar_auto_out_1_d_bits_source),
    .auto_out_1_d_bits_sink(system_bus_xbar_auto_out_1_d_bits_sink),
    .auto_out_1_d_bits_denied(system_bus_xbar_auto_out_1_d_bits_denied),
    .auto_out_1_d_bits_data(system_bus_xbar_auto_out_1_d_bits_data),
    .auto_out_1_d_bits_corrupt(system_bus_xbar_auto_out_1_d_bits_corrupt),
    .auto_out_1_e_valid(system_bus_xbar_auto_out_1_e_valid),
    .auto_out_1_e_bits_sink(system_bus_xbar_auto_out_1_e_bits_sink),
    .auto_out_0_a_ready(system_bus_xbar_auto_out_0_a_ready),
    .auto_out_0_a_valid(system_bus_xbar_auto_out_0_a_valid),
    .auto_out_0_a_bits_size(system_bus_xbar_auto_out_0_a_bits_size),
    .auto_out_0_a_bits_source(system_bus_xbar_auto_out_0_a_bits_source),
    .auto_out_0_a_bits_address(system_bus_xbar_auto_out_0_a_bits_address),
    .auto_out_0_a_bits_mask(system_bus_xbar_auto_out_0_a_bits_mask),
    .auto_out_0_d_ready(system_bus_xbar_auto_out_0_d_ready),
    .auto_out_0_d_valid(system_bus_xbar_auto_out_0_d_valid),
    .auto_out_0_d_bits_opcode(system_bus_xbar_auto_out_0_d_bits_opcode),
    .auto_out_0_d_bits_param(system_bus_xbar_auto_out_0_d_bits_param),
    .auto_out_0_d_bits_size(system_bus_xbar_auto_out_0_d_bits_size),
    .auto_out_0_d_bits_source(system_bus_xbar_auto_out_0_d_bits_source),
    .auto_out_0_d_bits_sink(system_bus_xbar_auto_out_0_d_bits_sink),
    .auto_out_0_d_bits_denied(system_bus_xbar_auto_out_0_d_bits_denied),
    .auto_out_0_d_bits_data(system_bus_xbar_auto_out_0_d_bits_data),
    .auto_out_0_d_bits_corrupt(system_bus_xbar_auto_out_0_d_bits_corrupt)
  );
  TLFIFOFixer fixer ( // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fixer_auto_in_a_bits_param),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_b_ready(fixer_auto_in_b_ready),
    .auto_in_b_valid(fixer_auto_in_b_valid),
    .auto_in_b_bits_param(fixer_auto_in_b_bits_param),
    .auto_in_b_bits_address(fixer_auto_in_b_bits_address),
    .auto_in_c_ready(fixer_auto_in_c_ready),
    .auto_in_c_valid(fixer_auto_in_c_valid),
    .auto_in_c_bits_opcode(fixer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(fixer_auto_in_c_bits_param),
    .auto_in_c_bits_size(fixer_auto_in_c_bits_size),
    .auto_in_c_bits_source(fixer_auto_in_c_bits_source),
    .auto_in_c_bits_address(fixer_auto_in_c_bits_address),
    .auto_in_c_bits_data(fixer_auto_in_c_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fixer_auto_in_d_bits_param),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fixer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_in_e_valid(fixer_auto_in_e_valid),
    .auto_in_e_bits_sink(fixer_auto_in_e_bits_sink),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fixer_auto_out_a_bits_param),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_b_ready(fixer_auto_out_b_ready),
    .auto_out_b_valid(fixer_auto_out_b_valid),
    .auto_out_b_bits_param(fixer_auto_out_b_bits_param),
    .auto_out_b_bits_address(fixer_auto_out_b_bits_address),
    .auto_out_c_ready(fixer_auto_out_c_ready),
    .auto_out_c_valid(fixer_auto_out_c_valid),
    .auto_out_c_bits_opcode(fixer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(fixer_auto_out_c_bits_param),
    .auto_out_c_bits_size(fixer_auto_out_c_bits_size),
    .auto_out_c_bits_source(fixer_auto_out_c_bits_source),
    .auto_out_c_bits_address(fixer_auto_out_c_bits_address),
    .auto_out_c_bits_data(fixer_auto_out_c_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fixer_auto_out_d_bits_param),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fixer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt),
    .auto_out_e_valid(fixer_auto_out_e_valid),
    .auto_out_e_bits_sink(fixer_auto_out_e_bits_sink)
  );
  TLInterconnectCoupler coupler_to_bus_named_subsystem_cbus ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_bus_named_subsystem_cbus_clock),
    .reset(coupler_to_bus_named_subsystem_cbus_reset),
    .auto_widget_in_a_ready(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready),
    .auto_widget_in_a_valid(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid),
    .auto_widget_in_a_bits_size(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size),
    .auto_widget_in_a_bits_source(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source),
    .auto_widget_in_a_bits_address(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address),
    .auto_widget_in_a_bits_mask(coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask),
    .auto_widget_in_d_ready(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready),
    .auto_widget_in_d_valid(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid),
    .auto_widget_in_d_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode),
    .auto_widget_in_d_bits_param(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param),
    .auto_widget_in_d_bits_size(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size),
    .auto_widget_in_d_bits_source(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source),
    .auto_widget_in_d_bits_sink(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink),
    .auto_widget_in_d_bits_denied(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied),
    .auto_widget_in_d_bits_data(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data),
    .auto_widget_in_d_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt),
    .auto_bus_xing_out_a_ready(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready),
    .auto_bus_xing_out_a_valid(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid),
    .auto_bus_xing_out_a_bits_size(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size),
    .auto_bus_xing_out_a_bits_source(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source),
    .auto_bus_xing_out_a_bits_address(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address),
    .auto_bus_xing_out_a_bits_mask(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask),
    .auto_bus_xing_out_d_ready(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready),
    .auto_bus_xing_out_d_valid(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid),
    .auto_bus_xing_out_d_bits_opcode(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode),
    .auto_bus_xing_out_d_bits_param(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param),
    .auto_bus_xing_out_d_bits_size(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size),
    .auto_bus_xing_out_d_bits_source(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source),
    .auto_bus_xing_out_d_bits_sink(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink),
    .auto_bus_xing_out_d_bits_denied(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied),
    .auto_bus_xing_out_d_bits_data(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data),
    .auto_bus_xing_out_d_bits_corrupt(coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt)
  );
  TLInterconnectCoupler_1 coupler_from_bus_named_subsystem_fbus ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_from_bus_named_subsystem_fbus_clock),
    .reset(coupler_from_bus_named_subsystem_fbus_reset)
  );
  TLInterconnectCoupler_2 coupler_to_bus_named_subsystem_l2 ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_bus_named_subsystem_l2_clock),
    .reset(coupler_to_bus_named_subsystem_l2_reset),
    .auto_widget_in_a_ready(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready),
    .auto_widget_in_a_valid(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid),
    .auto_widget_in_a_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode),
    .auto_widget_in_a_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_param),
    .auto_widget_in_a_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size),
    .auto_widget_in_a_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source),
    .auto_widget_in_a_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address),
    .auto_widget_in_a_bits_mask(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask),
    .auto_widget_in_a_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data),
    .auto_widget_in_b_ready(coupler_to_bus_named_subsystem_l2_auto_widget_in_b_ready),
    .auto_widget_in_b_valid(coupler_to_bus_named_subsystem_l2_auto_widget_in_b_valid),
    .auto_widget_in_b_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_param),
    .auto_widget_in_b_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_address),
    .auto_widget_in_c_ready(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_ready),
    .auto_widget_in_c_valid(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_valid),
    .auto_widget_in_c_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_opcode),
    .auto_widget_in_c_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_param),
    .auto_widget_in_c_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_size),
    .auto_widget_in_c_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_source),
    .auto_widget_in_c_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_address),
    .auto_widget_in_c_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_data),
    .auto_widget_in_d_ready(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready),
    .auto_widget_in_d_valid(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid),
    .auto_widget_in_d_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode),
    .auto_widget_in_d_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_param),
    .auto_widget_in_d_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size),
    .auto_widget_in_d_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source),
    .auto_widget_in_d_bits_sink(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_sink),
    .auto_widget_in_d_bits_denied(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied),
    .auto_widget_in_d_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data),
    .auto_widget_in_d_bits_corrupt(coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt),
    .auto_widget_in_e_valid(coupler_to_bus_named_subsystem_l2_auto_widget_in_e_valid),
    .auto_widget_in_e_bits_sink(coupler_to_bus_named_subsystem_l2_auto_widget_in_e_bits_sink),
    .auto_widget_out_a_ready(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready),
    .auto_widget_out_a_valid(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid),
    .auto_widget_out_a_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode),
    .auto_widget_out_a_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_param),
    .auto_widget_out_a_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size),
    .auto_widget_out_a_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source),
    .auto_widget_out_a_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address),
    .auto_widget_out_a_bits_mask(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask),
    .auto_widget_out_a_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data),
    .auto_widget_out_b_ready(coupler_to_bus_named_subsystem_l2_auto_widget_out_b_ready),
    .auto_widget_out_b_valid(coupler_to_bus_named_subsystem_l2_auto_widget_out_b_valid),
    .auto_widget_out_b_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_param),
    .auto_widget_out_b_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_address),
    .auto_widget_out_c_ready(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_ready),
    .auto_widget_out_c_valid(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_valid),
    .auto_widget_out_c_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_opcode),
    .auto_widget_out_c_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_param),
    .auto_widget_out_c_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_size),
    .auto_widget_out_c_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_source),
    .auto_widget_out_c_bits_address(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_address),
    .auto_widget_out_c_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_data),
    .auto_widget_out_d_ready(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready),
    .auto_widget_out_d_valid(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid),
    .auto_widget_out_d_bits_opcode(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode),
    .auto_widget_out_d_bits_param(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_param),
    .auto_widget_out_d_bits_size(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size),
    .auto_widget_out_d_bits_source(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source),
    .auto_widget_out_d_bits_sink(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_sink),
    .auto_widget_out_d_bits_denied(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied),
    .auto_widget_out_d_bits_data(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data),
    .auto_widget_out_d_bits_corrupt(coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt),
    .auto_widget_out_e_valid(coupler_to_bus_named_subsystem_l2_auto_widget_out_e_valid),
    .auto_widget_out_e_bits_sink(coupler_to_bus_named_subsystem_l2_auto_widget_out_e_bits_sink)
  );
  TLInterconnectCoupler_3 coupler_from_tile ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_from_tile_clock),
    .reset(coupler_from_tile_reset),
    .auto_tl_master_clock_xing_in_a_ready(coupler_from_tile_auto_tl_master_clock_xing_in_a_ready),
    .auto_tl_master_clock_xing_in_a_valid(coupler_from_tile_auto_tl_master_clock_xing_in_a_valid),
    .auto_tl_master_clock_xing_in_a_bits_opcode(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode),
    .auto_tl_master_clock_xing_in_a_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param),
    .auto_tl_master_clock_xing_in_a_bits_size(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size),
    .auto_tl_master_clock_xing_in_a_bits_source(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source),
    .auto_tl_master_clock_xing_in_a_bits_address(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address),
    .auto_tl_master_clock_xing_in_a_bits_mask(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask),
    .auto_tl_master_clock_xing_in_a_bits_data(coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data),
    .auto_tl_master_clock_xing_in_b_ready(coupler_from_tile_auto_tl_master_clock_xing_in_b_ready),
    .auto_tl_master_clock_xing_in_b_valid(coupler_from_tile_auto_tl_master_clock_xing_in_b_valid),
    .auto_tl_master_clock_xing_in_b_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_param),
    .auto_tl_master_clock_xing_in_b_bits_address(coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_address),
    .auto_tl_master_clock_xing_in_c_ready(coupler_from_tile_auto_tl_master_clock_xing_in_c_ready),
    .auto_tl_master_clock_xing_in_c_valid(coupler_from_tile_auto_tl_master_clock_xing_in_c_valid),
    .auto_tl_master_clock_xing_in_c_bits_opcode(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_opcode),
    .auto_tl_master_clock_xing_in_c_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_param),
    .auto_tl_master_clock_xing_in_c_bits_size(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_size),
    .auto_tl_master_clock_xing_in_c_bits_source(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_source),
    .auto_tl_master_clock_xing_in_c_bits_address(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_address),
    .auto_tl_master_clock_xing_in_c_bits_data(coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_data),
    .auto_tl_master_clock_xing_in_d_ready(coupler_from_tile_auto_tl_master_clock_xing_in_d_ready),
    .auto_tl_master_clock_xing_in_d_valid(coupler_from_tile_auto_tl_master_clock_xing_in_d_valid),
    .auto_tl_master_clock_xing_in_d_bits_opcode(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode),
    .auto_tl_master_clock_xing_in_d_bits_param(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param),
    .auto_tl_master_clock_xing_in_d_bits_size(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size),
    .auto_tl_master_clock_xing_in_d_bits_source(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source),
    .auto_tl_master_clock_xing_in_d_bits_sink(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink),
    .auto_tl_master_clock_xing_in_d_bits_denied(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied),
    .auto_tl_master_clock_xing_in_d_bits_data(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data),
    .auto_tl_master_clock_xing_in_d_bits_corrupt(coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt),
    .auto_tl_master_clock_xing_in_e_valid(coupler_from_tile_auto_tl_master_clock_xing_in_e_valid),
    .auto_tl_master_clock_xing_in_e_bits_sink(coupler_from_tile_auto_tl_master_clock_xing_in_e_bits_sink),
    .auto_tl_out_a_ready(coupler_from_tile_auto_tl_out_a_ready),
    .auto_tl_out_a_valid(coupler_from_tile_auto_tl_out_a_valid),
    .auto_tl_out_a_bits_opcode(coupler_from_tile_auto_tl_out_a_bits_opcode),
    .auto_tl_out_a_bits_param(coupler_from_tile_auto_tl_out_a_bits_param),
    .auto_tl_out_a_bits_size(coupler_from_tile_auto_tl_out_a_bits_size),
    .auto_tl_out_a_bits_source(coupler_from_tile_auto_tl_out_a_bits_source),
    .auto_tl_out_a_bits_address(coupler_from_tile_auto_tl_out_a_bits_address),
    .auto_tl_out_a_bits_mask(coupler_from_tile_auto_tl_out_a_bits_mask),
    .auto_tl_out_a_bits_data(coupler_from_tile_auto_tl_out_a_bits_data),
    .auto_tl_out_b_ready(coupler_from_tile_auto_tl_out_b_ready),
    .auto_tl_out_b_valid(coupler_from_tile_auto_tl_out_b_valid),
    .auto_tl_out_b_bits_param(coupler_from_tile_auto_tl_out_b_bits_param),
    .auto_tl_out_b_bits_address(coupler_from_tile_auto_tl_out_b_bits_address),
    .auto_tl_out_c_ready(coupler_from_tile_auto_tl_out_c_ready),
    .auto_tl_out_c_valid(coupler_from_tile_auto_tl_out_c_valid),
    .auto_tl_out_c_bits_opcode(coupler_from_tile_auto_tl_out_c_bits_opcode),
    .auto_tl_out_c_bits_param(coupler_from_tile_auto_tl_out_c_bits_param),
    .auto_tl_out_c_bits_size(coupler_from_tile_auto_tl_out_c_bits_size),
    .auto_tl_out_c_bits_source(coupler_from_tile_auto_tl_out_c_bits_source),
    .auto_tl_out_c_bits_address(coupler_from_tile_auto_tl_out_c_bits_address),
    .auto_tl_out_c_bits_data(coupler_from_tile_auto_tl_out_c_bits_data),
    .auto_tl_out_d_ready(coupler_from_tile_auto_tl_out_d_ready),
    .auto_tl_out_d_valid(coupler_from_tile_auto_tl_out_d_valid),
    .auto_tl_out_d_bits_opcode(coupler_from_tile_auto_tl_out_d_bits_opcode),
    .auto_tl_out_d_bits_param(coupler_from_tile_auto_tl_out_d_bits_param),
    .auto_tl_out_d_bits_size(coupler_from_tile_auto_tl_out_d_bits_size),
    .auto_tl_out_d_bits_source(coupler_from_tile_auto_tl_out_d_bits_source),
    .auto_tl_out_d_bits_sink(coupler_from_tile_auto_tl_out_d_bits_sink),
    .auto_tl_out_d_bits_denied(coupler_from_tile_auto_tl_out_d_bits_denied),
    .auto_tl_out_d_bits_data(coupler_from_tile_auto_tl_out_d_bits_data),
    .auto_tl_out_d_bits_corrupt(coupler_from_tile_auto_tl_out_d_bits_corrupt),
    .auto_tl_out_e_valid(coupler_from_tile_auto_tl_out_e_valid),
    .auto_tl_out_e_bits_sink(coupler_from_tile_auto_tl_out_e_bits_sink)
  );
  assign auto_coupler_from_tile_tl_master_clock_xing_in_a_ready = coupler_from_tile_auto_tl_master_clock_xing_in_a_ready
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_b_valid = coupler_from_tile_auto_tl_master_clock_xing_in_b_valid
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param =
    coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address =
    coupler_from_tile_auto_tl_master_clock_xing_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_c_ready = coupler_from_tile_auto_tl_master_clock_xing_in_c_ready
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_valid = coupler_from_tile_auto_tl_master_clock_xing_in_d_valid
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt =
    coupler_from_tile_auto_tl_master_clock_xing_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink =
    coupler_to_bus_named_subsystem_l2_auto_widget_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_1_clock = fixedClockNode_auto_out_2_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_1_reset = fixedClockNode_auto_out_2_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_0_clock = fixedClockNode_auto_out_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_0_reset = fixedClockNode_auto_out_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset =
    subsystem_sbus_clock_groups_auto_out_3_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_2_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_1_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_5_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_4_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_3_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_2_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_1_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_clock =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_sbus_clock_groups_auto_in_member_subsystem_sbus_0_reset =
    auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_sbus_0_clock =
    subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_sbus_0_reset =
    subsystem_sbus_clock_groups_auto_out_0_member_subsystem_sbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_param = fixer_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_b_ready = fixer_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_valid = fixer_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_opcode = fixer_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_param = fixer_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_size = fixer_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_source = fixer_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_address = fixer_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_c_bits_data = fixer_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_e_valid = fixer_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_in_e_bits_sink = fixer_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign system_bus_xbar_auto_out_1_a_ready = coupler_to_bus_named_subsystem_l2_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_b_valid = coupler_to_bus_named_subsystem_l2_auto_widget_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_b_bits_param = coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_b_bits_address = coupler_to_bus_named_subsystem_l2_auto_widget_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_c_ready = coupler_to_bus_named_subsystem_l2_auto_widget_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_valid = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_opcode = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_param = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_size = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_source = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_sink = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_denied = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_data = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_1_d_bits_corrupt = coupler_to_bus_named_subsystem_l2_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_a_ready = coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_valid = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_opcode = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_param = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_size = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_source = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_sink = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_denied = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_data = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign system_bus_xbar_auto_out_0_d_bits_corrupt = coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_valid = coupler_from_tile_auto_tl_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_opcode = coupler_from_tile_auto_tl_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_param = coupler_from_tile_auto_tl_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_size = coupler_from_tile_auto_tl_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_source = coupler_from_tile_auto_tl_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_address = coupler_from_tile_auto_tl_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_mask = coupler_from_tile_auto_tl_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_data = coupler_from_tile_auto_tl_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_b_ready = coupler_from_tile_auto_tl_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_valid = coupler_from_tile_auto_tl_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_opcode = coupler_from_tile_auto_tl_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_param = coupler_from_tile_auto_tl_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_size = coupler_from_tile_auto_tl_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_source = coupler_from_tile_auto_tl_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_address = coupler_from_tile_auto_tl_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_c_bits_data = coupler_from_tile_auto_tl_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_d_ready = coupler_from_tile_auto_tl_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_e_valid = coupler_from_tile_auto_tl_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_e_bits_sink = coupler_from_tile_auto_tl_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_a_ready = system_bus_xbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_b_valid = system_bus_xbar_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_b_bits_param = system_bus_xbar_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_b_bits_address = system_bus_xbar_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_c_ready = system_bus_xbar_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_valid = system_bus_xbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_opcode = system_bus_xbar_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_param = system_bus_xbar_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_size = system_bus_xbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_source = system_bus_xbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_sink = system_bus_xbar_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_denied = system_bus_xbar_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_data = system_bus_xbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_corrupt = system_bus_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_cbus_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_cbus_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_valid = system_bus_xbar_auto_out_0_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_size = system_bus_xbar_auto_out_0_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_source = system_bus_xbar_auto_out_0_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_address = system_bus_xbar_auto_out_0_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_a_bits_mask = system_bus_xbar_auto_out_0_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_widget_in_d_ready = system_bus_xbar_auto_out_0_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_a_ready =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_valid =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_param =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_sink =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_cbus_auto_bus_xing_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_from_bus_named_subsystem_fbus_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_bus_named_subsystem_fbus_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_l2_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_l2_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_valid = system_bus_xbar_auto_out_1_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_opcode = system_bus_xbar_auto_out_1_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_param = system_bus_xbar_auto_out_1_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_size = system_bus_xbar_auto_out_1_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_source = system_bus_xbar_auto_out_1_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_address = system_bus_xbar_auto_out_1_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_mask = system_bus_xbar_auto_out_1_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_a_bits_data = system_bus_xbar_auto_out_1_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_b_ready = system_bus_xbar_auto_out_1_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_valid = system_bus_xbar_auto_out_1_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_opcode = system_bus_xbar_auto_out_1_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_param = system_bus_xbar_auto_out_1_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_size = system_bus_xbar_auto_out_1_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_source = system_bus_xbar_auto_out_1_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_address = system_bus_xbar_auto_out_1_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_c_bits_data = system_bus_xbar_auto_out_1_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_d_ready = system_bus_xbar_auto_out_1_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_e_valid = system_bus_xbar_auto_out_1_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_in_e_bits_sink = system_bus_xbar_auto_out_1_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_a_ready =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_b_valid =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_param =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_b_bits_address =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_c_ready =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_valid =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_param =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_sink =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_l2_auto_widget_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_from_tile_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_valid = auto_coupler_from_tile_tl_master_clock_xing_in_a_valid
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_opcode =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_param =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_size =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_source =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_address =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_mask =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_a_bits_data =
    auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_b_ready = auto_coupler_from_tile_tl_master_clock_xing_in_b_ready
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_valid = auto_coupler_from_tile_tl_master_clock_xing_in_c_valid
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_opcode =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_param =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_size =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_source =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_address =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_c_bits_data =
    auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_d_ready = auto_coupler_from_tile_tl_master_clock_xing_in_d_ready
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_e_valid = auto_coupler_from_tile_tl_master_clock_xing_in_e_valid
    ; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_master_clock_xing_in_e_bits_sink =
    auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coupler_from_tile_auto_tl_out_a_ready = fixer_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_b_valid = fixer_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_b_bits_param = fixer_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_b_bits_address = fixer_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_c_ready = fixer_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_valid = fixer_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_param = fixer_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_size = fixer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_source = fixer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_sink = fixer_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_data = fixer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_from_tile_auto_tl_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module ClockGroupAggregator_1(
  input   auto_in_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_pbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_pbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_member_subsystem_pbus_0_clock = auto_in_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_member_subsystem_pbus_0_reset = auto_in_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup_1(
  input   auto_in_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_pbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_1(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_1(
  input   clock,
  input   reset
);
endmodule
module TLFIFOFixer_1(
  input   clock,
  input   reset
);
endmodule
module TLXbar_1(
  input   clock,
  input   reset
);
endmodule
module TLXbar_2(
  input   clock,
  input   reset
);
endmodule
module TLBuffer(
  input   clock,
  input   reset
);
endmodule
module TLAtomicAutomata(
  input   clock,
  input   reset
);
endmodule
module TLBuffer_1(
  input   clock,
  input   reset
);
endmodule
module PeripheryBus(
  input   auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output  reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_pbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_pbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  fixer_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  in_xbar_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  out_xbar_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  atomics_clock; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_reset; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  buffer_1_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  ClockGroupAggregator_1 subsystem_pbus_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_pbus_0_clock(subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock),
    .auto_in_member_subsystem_pbus_0_reset(subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset),
    .auto_out_member_subsystem_pbus_0_clock(subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock),
    .auto_out_member_subsystem_pbus_0_reset(subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset)
  );
  ClockGroup_1 clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_pbus_0_clock(clockGroup_auto_in_member_subsystem_pbus_0_clock),
    .auto_in_member_subsystem_pbus_0_reset(clockGroup_auto_in_member_subsystem_pbus_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast_1 fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_clock(fixedClockNode_auto_out_clock),
    .auto_out_reset(fixedClockNode_auto_out_reset)
  );
  BundleBridgeNexus_1 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLFIFOFixer_1 fixer ( // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
    .clock(fixer_clock),
    .reset(fixer_reset)
  );
  TLXbar_1 in_xbar ( // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
    .clock(in_xbar_clock),
    .reset(in_xbar_reset)
  );
  TLXbar_2 out_xbar ( // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
    .clock(out_xbar_clock),
    .reset(out_xbar_reset)
  );
  TLBuffer buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset)
  );
  TLAtomicAutomata atomics ( // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
    .clock(atomics_clock),
    .reset(atomics_reset)
  );
  TLBuffer_1 buffer_1 ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset)
  );
  assign clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_clock =
    auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_pbus_clock_groups_auto_in_member_subsystem_pbus_0_reset =
    auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_pbus_0_clock =
    subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_pbus_0_reset =
    subsystem_pbus_clock_groups_auto_out_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign out_xbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign out_xbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module ClockGroupAggregator_2(
  input   auto_in_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_fbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_fbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_member_subsystem_fbus_0_clock = auto_in_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_member_subsystem_fbus_0_reset = auto_in_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup_2(
  input   auto_in_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_fbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_2(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_2(
  input   clock,
  input   reset
);
endmodule
module TLXbar_3(
  input   clock,
  input   reset
);
endmodule
module TLBuffer_2(
  input   clock,
  input   reset
);
endmodule
module FrontBus(
  input   auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output  reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_fbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_fbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  subsystem_fbus_xbar_clock; // @[src/main/scala/tilelink/BusWrapper.scala 221:32]
  wire  subsystem_fbus_xbar_reset; // @[src/main/scala/tilelink/BusWrapper.scala 221:32]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  ClockGroupAggregator_2 subsystem_fbus_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_fbus_0_clock(subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock),
    .auto_in_member_subsystem_fbus_0_reset(subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset),
    .auto_out_member_subsystem_fbus_0_clock(subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock),
    .auto_out_member_subsystem_fbus_0_reset(subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset)
  );
  ClockGroup_2 clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_fbus_0_clock(clockGroup_auto_in_member_subsystem_fbus_0_clock),
    .auto_in_member_subsystem_fbus_0_reset(clockGroup_auto_in_member_subsystem_fbus_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast_2 fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_clock(fixedClockNode_auto_out_clock),
    .auto_out_reset(fixedClockNode_auto_out_reset)
  );
  BundleBridgeNexus_2 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLXbar_3 subsystem_fbus_xbar ( // @[src/main/scala/tilelink/BusWrapper.scala 221:32]
    .clock(subsystem_fbus_xbar_clock),
    .reset(subsystem_fbus_xbar_reset)
  );
  TLBuffer_2 buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset)
  );
  assign clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_clock =
    auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_fbus_clock_groups_auto_in_member_subsystem_fbus_0_reset =
    auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_fbus_0_clock =
    subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_fbus_0_reset =
    subsystem_fbus_clock_groups_auto_out_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_fbus_xbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_fbus_xbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module ClockGroupAggregator_3(
  input   auto_in_member_subsystem_cbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_cbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_cbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_pbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_cbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_1_member_subsystem_pbus_0_clock = auto_in_member_subsystem_cbus_1_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_pbus_0_reset = auto_in_member_subsystem_cbus_1_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_cbus_0_clock = auto_in_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_cbus_0_reset = auto_in_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup_3(
  input   auto_in_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_cbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_3(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_1_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_3(
  input   clock,
  input   reset
);
endmodule
module TLFIFOFixer_2(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  a_first_done = auto_out_a_ready & auto_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [1:0] a_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] a_first_counter1 = a_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_17_clock;
  wire  line_17_reset;
  wire  line_17_valid;
  reg  line_17_valid_reg;
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _d_first_beats1_decode_T_1 = 12'h1f << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  reg [1:0] d_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] d_first_counter1 = d_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  d_first_first = d_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_18_clock;
  wire  line_18_reset;
  wire  line_18_valid;
  reg  line_18_valid_reg;
  wire  _T_1 = a_first & a_first_done; // @[src/main/scala/tilelink/FIFOFixer.scala 74:21]
  wire  line_19_clock;
  wire  line_19_reset;
  wire  line_19_valid;
  reg  line_19_valid_reg;
  wire  line_20_clock;
  wire  line_20_reset;
  wire  line_20_valid;
  reg  line_20_valid_reg;
  wire  line_21_clock;
  wire  line_21_reset;
  wire  line_21_valid;
  reg  line_21_valid_reg;
  wire  line_22_clock;
  wire  line_22_reset;
  wire  line_22_valid;
  reg  line_22_valid_reg;
  wire  _T_3 = d_first_first & _d_first_T; // @[src/main/scala/tilelink/FIFOFixer.scala 75:21]
  wire  line_23_clock;
  wire  line_23_reset;
  wire  line_23_valid;
  reg  line_23_valid_reg;
  wire  line_24_clock;
  wire  line_24_reset;
  wire  line_24_valid;
  reg  line_24_valid_reg;
  wire  line_25_clock;
  wire  line_25_reset;
  wire  line_25_valid;
  reg  line_25_valid_reg;
  wire  line_26_clock;
  wire  line_26_reset;
  wire  line_26_valid;
  reg  line_26_valid_reg;
  wire  line_27_clock;
  wire  line_27_reset;
  wire  line_27_valid;
  reg  line_27_valid_reg;
  wire  line_28_clock;
  wire  line_28_reset;
  wire  line_28_valid;
  reg  line_28_valid_reg;
  GEN_w1_line #(.COVER_INDEX(17)) line_17 (
    .clock(line_17_clock),
    .reset(line_17_reset),
    .valid(line_17_valid)
  );
  GEN_w1_line #(.COVER_INDEX(18)) line_18 (
    .clock(line_18_clock),
    .reset(line_18_reset),
    .valid(line_18_valid)
  );
  GEN_w1_line #(.COVER_INDEX(19)) line_19 (
    .clock(line_19_clock),
    .reset(line_19_reset),
    .valid(line_19_valid)
  );
  GEN_w1_line #(.COVER_INDEX(20)) line_20 (
    .clock(line_20_clock),
    .reset(line_20_reset),
    .valid(line_20_valid)
  );
  GEN_w1_line #(.COVER_INDEX(21)) line_21 (
    .clock(line_21_clock),
    .reset(line_21_reset),
    .valid(line_21_valid)
  );
  GEN_w1_line #(.COVER_INDEX(22)) line_22 (
    .clock(line_22_clock),
    .reset(line_22_reset),
    .valid(line_22_valid)
  );
  GEN_w1_line #(.COVER_INDEX(23)) line_23 (
    .clock(line_23_clock),
    .reset(line_23_reset),
    .valid(line_23_valid)
  );
  GEN_w1_line #(.COVER_INDEX(24)) line_24 (
    .clock(line_24_clock),
    .reset(line_24_reset),
    .valid(line_24_valid)
  );
  GEN_w1_line #(.COVER_INDEX(25)) line_25 (
    .clock(line_25_clock),
    .reset(line_25_reset),
    .valid(line_25_valid)
  );
  GEN_w1_line #(.COVER_INDEX(26)) line_26 (
    .clock(line_26_clock),
    .reset(line_26_reset),
    .valid(line_26_valid)
  );
  GEN_w1_line #(.COVER_INDEX(27)) line_27 (
    .clock(line_27_clock),
    .reset(line_27_reset),
    .valid(line_27_valid)
  );
  GEN_w1_line #(.COVER_INDEX(28)) line_28 (
    .clock(line_28_clock),
    .reset(line_28_reset),
    .valid(line_28_valid)
  );
  assign line_17_clock = clock;
  assign line_17_reset = reset;
  assign line_17_valid = a_first_done ^ line_17_valid_reg;
  assign line_18_clock = clock;
  assign line_18_reset = reset;
  assign line_18_valid = _d_first_T ^ line_18_valid_reg;
  assign line_19_clock = clock;
  assign line_19_reset = reset;
  assign line_19_valid = _T_1 ^ line_19_valid_reg;
  assign line_20_clock = clock;
  assign line_20_reset = reset;
  assign line_20_valid = 2'h0 == auto_in_a_bits_source ^ line_20_valid_reg;
  assign line_21_clock = clock;
  assign line_21_reset = reset;
  assign line_21_valid = 2'h1 == auto_in_a_bits_source ^ line_21_valid_reg;
  assign line_22_clock = clock;
  assign line_22_reset = reset;
  assign line_22_valid = 2'h2 == auto_in_a_bits_source ^ line_22_valid_reg;
  assign line_23_clock = clock;
  assign line_23_reset = reset;
  assign line_23_valid = _T_3 ^ line_23_valid_reg;
  assign line_24_clock = clock;
  assign line_24_reset = reset;
  assign line_24_valid = 2'h0 == auto_out_d_bits_source ^ line_24_valid_reg;
  assign line_25_clock = clock;
  assign line_25_reset = reset;
  assign line_25_valid = 2'h1 == auto_out_d_bits_source ^ line_25_valid_reg;
  assign line_26_clock = clock;
  assign line_26_reset = reset;
  assign line_26_valid = 2'h2 == auto_out_d_bits_source ^ line_26_valid_reg;
  assign line_27_clock = clock;
  assign line_27_reset = reset;
  assign line_27_valid = _T_1 ^ line_27_valid_reg;
  assign line_28_clock = clock;
  assign line_28_reset = reset;
  assign line_28_valid = _T_3 ^ line_28_valid_reg;
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 90:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 89:33]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      a_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (a_first_done) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (a_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        a_first_counter <= 2'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    line_17_valid_reg <= a_first_done;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      d_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_d_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (d_first_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        d_first_counter <= d_first_beats1_decode;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    line_18_valid_reg <= _d_first_T;
    line_19_valid_reg <= _T_1;
    line_20_valid_reg <= 2'h0 == auto_in_a_bits_source;
    line_21_valid_reg <= 2'h1 == auto_in_a_bits_source;
    line_22_valid_reg <= 2'h2 == auto_in_a_bits_source;
    line_23_valid_reg <= _T_3;
    line_24_valid_reg <= 2'h0 == auto_out_d_bits_source;
    line_25_valid_reg <= 2'h1 == auto_out_d_bits_source;
    line_26_valid_reg <= 2'h2 == auto_out_d_bits_source;
    line_27_valid_reg <= _T_1;
    line_28_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_17_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  d_first_counter = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  line_18_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_19_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_20_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_21_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_22_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_23_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_24_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_25_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_26_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_27_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_28_valid_reg = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_4(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 248:53]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLXbar_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [28:0] io_enq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [28:0] io_deq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [28:0] ram_address [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [28:0] ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_mask [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_29_clock;
  wire  line_29_reset;
  wire  line_29_valid;
  reg  line_29_valid_reg;
  wire  line_30_clock;
  wire  line_30_reset;
  wire  line_30_valid;
  reg  line_30_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_31_clock;
  wire  line_31_reset;
  wire  line_31_valid;
  reg  line_31_valid_reg;
  GEN_w1_line #(.COVER_INDEX(29)) line_29 (
    .clock(line_29_clock),
    .reset(line_29_reset),
    .valid(line_29_valid)
  );
  GEN_w1_line #(.COVER_INDEX(30)) line_30 (
    .clock(line_30_clock),
    .reset(line_30_reset),
    .valid(line_30_valid)
  );
  GEN_w1_line #(.COVER_INDEX(31)) line_31 (
    .clock(line_31_clock),
    .reset(line_31_reset),
    .valid(line_31_valid)
  );
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_29_clock = clock;
  assign line_29_reset = reset;
  assign line_29_valid = do_enq ^ line_29_valid_reg;
  assign line_30_clock = clock;
  assign line_30_reset = reset;
  assign line_30_valid = do_deq ^ line_30_valid_reg;
  assign line_31_clock = clock;
  assign line_31_reset = reset;
  assign line_31_valid = _T ^ line_31_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_29_valid_reg <= do_enq;
    line_30_valid_reg <= do_deq;
    line_31_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_2[28:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_3[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_29_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_30_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_31_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_sink, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_denied, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_corrupt // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_param [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_sink [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_denied [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_corrupt [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_32_clock;
  wire  line_32_reset;
  wire  line_32_valid;
  reg  line_32_valid_reg;
  wire  line_33_clock;
  wire  line_33_reset;
  wire  line_33_valid;
  reg  line_33_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_34_clock;
  wire  line_34_reset;
  wire  line_34_valid;
  reg  line_34_valid_reg;
  GEN_w1_line #(.COVER_INDEX(32)) line_32 (
    .clock(line_32_clock),
    .reset(line_32_reset),
    .valid(line_32_valid)
  );
  GEN_w1_line #(.COVER_INDEX(33)) line_33 (
    .clock(line_33_clock),
    .reset(line_33_reset),
    .valid(line_33_valid)
  );
  GEN_w1_line #(.COVER_INDEX(34)) line_34 (
    .clock(line_34_clock),
    .reset(line_34_reset),
    .valid(line_34_valid)
  );
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_opcode_MPORT_data = 3'h1;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = enq_ptr_value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sink_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = enq_ptr_value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = enq_ptr_value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = enq_ptr_value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_32_clock = clock;
  assign line_32_reset = reset;
  assign line_32_valid = do_enq ^ line_32_valid_reg;
  assign line_33_clock = clock;
  assign line_33_reset = reset;
  assign line_33_valid = do_deq ^ line_33_valid_reg;
  assign line_34_clock = clock;
  assign line_34_reset = reset;
  assign line_34_valid = _T ^ line_34_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_32_valid_reg <= do_enq;
    line_33_valid_reg <= do_deq;
    line_34_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_32_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_33_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_34_valid_reg = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_3(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  nodeOut_a_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_a_q_io_enq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [28:0] nodeOut_a_q_io_enq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_a_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_a_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [28:0] nodeOut_a_q_io_deq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_a_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_enq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_d_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_deq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_deq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_bits_sink; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_bits_denied; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_d_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_bits_corrupt; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  Queue nodeOut_a_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_a_q_clock),
    .reset(nodeOut_a_q_reset),
    .io_enq_ready(nodeOut_a_q_io_enq_ready),
    .io_enq_valid(nodeOut_a_q_io_enq_valid),
    .io_enq_bits_size(nodeOut_a_q_io_enq_bits_size),
    .io_enq_bits_source(nodeOut_a_q_io_enq_bits_source),
    .io_enq_bits_address(nodeOut_a_q_io_enq_bits_address),
    .io_enq_bits_mask(nodeOut_a_q_io_enq_bits_mask),
    .io_deq_ready(nodeOut_a_q_io_deq_ready),
    .io_deq_valid(nodeOut_a_q_io_deq_valid),
    .io_deq_bits_size(nodeOut_a_q_io_deq_bits_size),
    .io_deq_bits_source(nodeOut_a_q_io_deq_bits_source),
    .io_deq_bits_address(nodeOut_a_q_io_deq_bits_address),
    .io_deq_bits_mask(nodeOut_a_q_io_deq_bits_mask)
  );
  Queue_1 nodeIn_d_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeIn_d_q_clock),
    .reset(nodeIn_d_q_reset),
    .io_enq_ready(nodeIn_d_q_io_enq_ready),
    .io_enq_valid(nodeIn_d_q_io_enq_valid),
    .io_enq_bits_size(nodeIn_d_q_io_enq_bits_size),
    .io_enq_bits_source(nodeIn_d_q_io_enq_bits_source),
    .io_enq_bits_data(nodeIn_d_q_io_enq_bits_data),
    .io_deq_ready(nodeIn_d_q_io_deq_ready),
    .io_deq_valid(nodeIn_d_q_io_deq_valid),
    .io_deq_bits_opcode(nodeIn_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(nodeIn_d_q_io_deq_bits_param),
    .io_deq_bits_size(nodeIn_d_q_io_deq_bits_size),
    .io_deq_bits_source(nodeIn_d_q_io_deq_bits_source),
    .io_deq_bits_sink(nodeIn_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(nodeIn_d_q_io_deq_bits_denied),
    .io_deq_bits_data(nodeIn_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(nodeIn_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = nodeOut_a_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_d_valid = nodeIn_d_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_opcode = nodeIn_d_q_io_deq_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_param = nodeIn_d_q_io_deq_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_size = nodeIn_d_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_source = nodeIn_d_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_sink = nodeIn_d_q_io_deq_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_denied = nodeIn_d_q_io_deq_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_data = nodeIn_d_q_io_deq_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_corrupt = nodeIn_d_q_io_deq_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_out_a_valid = nodeOut_a_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_size = nodeOut_a_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_source = nodeOut_a_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_address = nodeOut_a_q_io_deq_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_mask = nodeOut_a_q_io_deq_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_d_ready = nodeIn_d_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign nodeOut_a_q_clock = clock;
  assign nodeOut_a_q_reset = reset;
  assign nodeOut_a_q_io_enq_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_deq_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_clock = clock;
  assign nodeIn_d_q_reset = reset;
  assign nodeIn_d_q_io_enq_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_deq_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLAtomicAutomata_1(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLBuffer_4(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLWidthWidget_3(
  input   clock,
  input   reset
);
endmodule
module TLInterconnectCoupler_4(
  input   clock,
  input   reset
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget_3 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset)
  );
  assign widget_clock = clock;
  assign widget_reset = reset;
endmodule
module TLWidthWidget_4(
  input   clock,
  input   reset
);
endmodule
module TLInterconnectCoupler_5(
  input   clock,
  input   reset
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget_4 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset)
  );
  assign widget_clock = clock;
  assign widget_reset = reset;
endmodule
module Repeater(
  input         clock,
  input         reset,
  input         io_repeat, // @[src/main/scala/util/Repeater.scala 12:14]
  output        io_full, // @[src/main/scala/util/Repeater.scala 12:14]
  output        io_enq_ready, // @[src/main/scala/util/Repeater.scala 12:14]
  input         io_enq_valid, // @[src/main/scala/util/Repeater.scala 12:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/util/Repeater.scala 12:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/util/Repeater.scala 12:14]
  input  [28:0] io_enq_bits_address, // @[src/main/scala/util/Repeater.scala 12:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/util/Repeater.scala 12:14]
  input         io_deq_ready, // @[src/main/scala/util/Repeater.scala 12:14]
  output        io_deq_valid, // @[src/main/scala/util/Repeater.scala 12:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/util/Repeater.scala 12:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/util/Repeater.scala 12:14]
  output [28:0] io_deq_bits_address, // @[src/main/scala/util/Repeater.scala 12:14]
  output [7:0]  io_deq_bits_mask // @[src/main/scala/util/Repeater.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[src/main/scala/util/Repeater.scala 19:21]
  reg [2:0] saved_size; // @[src/main/scala/util/Repeater.scala 20:18]
  reg [1:0] saved_source; // @[src/main/scala/util/Repeater.scala 20:18]
  reg [28:0] saved_address; // @[src/main/scala/util/Repeater.scala 20:18]
  reg [7:0] saved_mask; // @[src/main/scala/util/Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & io_repeat; // @[src/main/scala/util/Repeater.scala 28:21]
  wire  line_35_clock;
  wire  line_35_reset;
  wire  line_35_valid;
  reg  line_35_valid_reg;
  wire  _GEN_2 = _T & io_repeat | full; // @[src/main/scala/util/Repeater.scala 19:21 28:{36,43}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_4 = _T_2 & ~io_repeat; // @[src/main/scala/util/Repeater.scala 29:21]
  wire  line_36_clock;
  wire  line_36_reset;
  wire  line_36_valid;
  reg  line_36_valid_reg;
  GEN_w1_line #(.COVER_INDEX(35)) line_35 (
    .clock(line_35_clock),
    .reset(line_35_reset),
    .valid(line_35_valid)
  );
  GEN_w1_line #(.COVER_INDEX(36)) line_36 (
    .clock(line_36_clock),
    .reset(line_36_reset),
    .valid(line_36_valid)
  );
  assign line_35_clock = clock;
  assign line_35_reset = reset;
  assign line_35_valid = _T_1 ^ line_35_valid_reg;
  assign line_36_clock = clock;
  assign line_36_reset = reset;
  assign line_36_valid = _T_4 ^ line_36_valid_reg;
  assign io_full = full; // @[src/main/scala/util/Repeater.scala 26:11]
  assign io_enq_ready = io_deq_ready & ~full; // @[src/main/scala/util/Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[src/main/scala/util/Repeater.scala 23:32]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[src/main/scala/util/Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[src/main/scala/util/Repeater.scala 25:21]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[src/main/scala/util/Repeater.scala 25:21]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[src/main/scala/util/Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/util/Repeater.scala 19:21]
      full <= 1'h0; // @[src/main/scala/util/Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[src/main/scala/util/Repeater.scala 29:36]
      full <= 1'h0; // @[src/main/scala/util/Repeater.scala 29:43]
    end else begin
      full <= _GEN_2;
    end
    if (_T & io_repeat) begin // @[src/main/scala/util/Repeater.scala 28:36]
      saved_size <= io_enq_bits_size; // @[src/main/scala/util/Repeater.scala 28:60]
    end
    if (_T & io_repeat) begin // @[src/main/scala/util/Repeater.scala 28:36]
      saved_source <= io_enq_bits_source; // @[src/main/scala/util/Repeater.scala 28:60]
    end
    if (_T & io_repeat) begin // @[src/main/scala/util/Repeater.scala 28:36]
      saved_address <= io_enq_bits_address; // @[src/main/scala/util/Repeater.scala 28:60]
    end
    if (_T & io_repeat) begin // @[src/main/scala/util/Repeater.scala 28:36]
      saved_mask <= io_enq_bits_mask; // @[src/main/scala/util/Repeater.scala 28:60]
    end
    line_35_valid_reg <= _T_1;
    line_36_valid_reg <= _T_4;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_size = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_source = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  saved_address = _RAND_3[28:0];
  _RAND_4 = {1{`RANDOM}};
  saved_mask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  line_35_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_36_valid_reg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [4:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [4:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  repeater_clock; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_reset; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_repeat; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_full; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_enq_ready; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_enq_valid; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [2:0] repeater_io_enq_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [1:0] repeater_io_enq_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [28:0] repeater_io_enq_bits_address; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [7:0] repeater_io_enq_bits_mask; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_deq_ready; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire  repeater_io_deq_valid; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [2:0] repeater_io_deq_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [1:0] repeater_io_deq_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [28:0] repeater_io_deq_bits_address; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  wire [7:0] repeater_io_deq_bits_mask; // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
  reg [1:0] acknum; // @[src/main/scala/tilelink/Fragmenter.scala 191:29]
  reg [2:0] dOrig; // @[src/main/scala/tilelink/Fragmenter.scala 192:24]
  reg  dToggle; // @[src/main/scala/tilelink/Fragmenter.scala 193:30]
  wire [1:0] dFragnum = auto_out_d_bits_source[1:0]; // @[src/main/scala/tilelink/Fragmenter.scala 194:41]
  wire  dFirst = acknum == 2'h0; // @[src/main/scala/tilelink/Fragmenter.scala 195:29]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[src/main/scala/util/package.scala 235:46]
  wire  _T_5 = ~reset; // @[src/main/scala/tilelink/Fragmenter.scala 204:16]
  wire  line_37_clock;
  wire  line_37_reset;
  wire  line_37_valid;
  reg  line_37_valid_reg;
  wire [4:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[src/main/scala/tilelink/Fragmenter.scala 208:47]
  wire [4:0] _GEN_17 = {{2'd0}, dsizeOH1}; // @[src/main/scala/tilelink/Fragmenter.scala 208:69]
  wire [4:0] _dFirst_size_T_1 = _dFirst_size_T | _GEN_17; // @[src/main/scala/tilelink/Fragmenter.scala 208:69]
  wire [5:0] _dFirst_size_T_2 = {_dFirst_size_T_1, 1'h0}; // @[src/main/scala/util/package.scala 233:35]
  wire [5:0] _dFirst_size_T_3 = _dFirst_size_T_2 | 6'h1; // @[src/main/scala/util/package.scala 233:40]
  wire [5:0] _dFirst_size_T_4 = {1'h0,_dFirst_size_T_1}; // @[src/main/scala/util/package.scala 233:53]
  wire [5:0] _dFirst_size_T_5 = ~_dFirst_size_T_4; // @[src/main/scala/util/package.scala 233:49]
  wire [5:0] _dFirst_size_T_6 = _dFirst_size_T_3 & _dFirst_size_T_5; // @[src/main/scala/util/package.scala 233:47]
  wire [1:0] dFirst_size_hi = _dFirst_size_T_6[5:4]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [3:0] dFirst_size_lo = _dFirst_size_T_6[3:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [3:0] _GEN_18 = {{2'd0}, dFirst_size_hi}; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [3:0] _dFirst_size_T_8 = _GEN_18 | dFirst_size_lo; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [1:0] dFirst_size_hi_1 = _dFirst_size_T_8[3:2]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [1:0] dFirst_size_lo_1 = _dFirst_size_T_8[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [1:0] _dFirst_size_T_10 = dFirst_size_hi_1 | dFirst_size_lo_1; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [2:0] dFirst_size = {|dFirst_size_hi,|dFirst_size_hi_1,_dFirst_size_T_10[1]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:10]
  wire  _T_7 = auto_in_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_38_clock;
  wire  line_38_reset;
  wire  line_38_valid;
  reg  line_38_valid_reg;
  wire [1:0] _acknum_T_1 = acknum - 2'h1; // @[src/main/scala/tilelink/Fragmenter.scala 211:55]
  wire  line_39_clock;
  wire  line_39_reset;
  wire  line_39_valid;
  reg  line_39_valid_reg;
  wire [2:0] aFrag = repeater_io_deq_bits_size > 3'h3 ? 3'h3 : repeater_io_deq_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 287:24]
  wire [11:0] _aOrigOH1_T_1 = 12'h1f << repeater_io_deq_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] aOrigOH1 = ~_aOrigOH1_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[src/main/scala/util/package.scala 235:71]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[src/main/scala/util/package.scala 235:46]
  reg [1:0] gennum; // @[src/main/scala/tilelink/Fragmenter.scala 293:29]
  wire  aFirst = gennum == 2'h0; // @[src/main/scala/tilelink/Fragmenter.scala 294:29]
  wire [1:0] _old_gennum1_T_2 = gennum - 2'h1; // @[src/main/scala/tilelink/Fragmenter.scala 295:79]
  wire [1:0] old_gennum1 = aFirst ? aOrigOH1[4:3] : _old_gennum1_T_2; // @[src/main/scala/tilelink/Fragmenter.scala 295:30]
  wire [1:0] _new_gennum_T = ~old_gennum1; // @[src/main/scala/tilelink/Fragmenter.scala 296:28]
  wire [1:0] new_gennum = ~_new_gennum_T; // @[src/main/scala/tilelink/Fragmenter.scala 296:26]
  reg  aToggle_r; // @[src/main/scala/tilelink/Fragmenter.scala 299:54]
  wire  line_40_clock;
  wire  line_40_reset;
  wire  line_40_valid;
  reg  line_40_valid_reg;
  wire  _GEN_15 = aFirst ? dToggle : aToggle_r; // @[src/main/scala/tilelink/Fragmenter.scala 299:{54,54,54}]
  wire  aToggle = ~_GEN_15; // @[src/main/scala/tilelink/Fragmenter.scala 299:23]
  wire  nodeOut_a_valid = repeater_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Fragmenter.scala 305:15]
  wire  _T_8 = auto_out_a_ready & nodeOut_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_41_clock;
  wire  line_41_reset;
  wire  line_41_valid;
  reg  line_41_valid_reg;
  wire [4:0] _nodeOut_a_bits_address_T = {old_gennum1, 3'h0}; // @[src/main/scala/tilelink/Fragmenter.scala 306:65]
  wire [4:0] _nodeOut_a_bits_address_T_1 = ~aOrigOH1; // @[src/main/scala/tilelink/Fragmenter.scala 306:90]
  wire [4:0] _nodeOut_a_bits_address_T_2 = _nodeOut_a_bits_address_T | _nodeOut_a_bits_address_T_1; // @[src/main/scala/tilelink/Fragmenter.scala 306:88]
  wire [4:0] _GEN_19 = {{2'd0}, aFragOH1}; // @[src/main/scala/tilelink/Fragmenter.scala 306:100]
  wire [4:0] _nodeOut_a_bits_address_T_3 = _nodeOut_a_bits_address_T_2 | _GEN_19; // @[src/main/scala/tilelink/Fragmenter.scala 306:100]
  wire [4:0] _nodeOut_a_bits_address_T_4 = _nodeOut_a_bits_address_T_3 | 5'h7; // @[src/main/scala/tilelink/Fragmenter.scala 306:111]
  wire [4:0] _nodeOut_a_bits_address_T_5 = ~_nodeOut_a_bits_address_T_4; // @[src/main/scala/tilelink/Fragmenter.scala 306:51]
  wire [28:0] _GEN_20 = {{24'd0}, _nodeOut_a_bits_address_T_5}; // @[src/main/scala/tilelink/Fragmenter.scala 306:49]
  wire [2:0] nodeOut_a_bits_source_hi = {repeater_io_deq_bits_source,aToggle}; // @[src/main/scala/tilelink/Fragmenter.scala 307:33]
  wire  _T_9 = ~repeater_io_full; // @[src/main/scala/tilelink/Fragmenter.scala 311:17]
  wire  line_42_clock;
  wire  line_42_reset;
  wire  line_42_valid;
  reg  line_42_valid_reg;
  wire  line_43_clock;
  wire  line_43_reset;
  wire  line_43_valid;
  reg  line_43_valid_reg;
  wire  _T_20 = ~(_T_9 | repeater_io_deq_bits_mask == 8'hff); // @[src/main/scala/tilelink/Fragmenter.scala 314:16]
  wire  line_44_clock;
  wire  line_44_reset;
  wire  line_44_valid;
  reg  line_44_valid_reg;
  Repeater repeater ( // @[src/main/scala/tilelink/Fragmenter.scala 264:30]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask)
  );
  GEN_w1_line #(.COVER_INDEX(37)) line_37 (
    .clock(line_37_clock),
    .reset(line_37_reset),
    .valid(line_37_valid)
  );
  GEN_w1_line #(.COVER_INDEX(38)) line_38 (
    .clock(line_38_clock),
    .reset(line_38_reset),
    .valid(line_38_valid)
  );
  GEN_w1_line #(.COVER_INDEX(39)) line_39 (
    .clock(line_39_clock),
    .reset(line_39_reset),
    .valid(line_39_valid)
  );
  GEN_w1_line #(.COVER_INDEX(40)) line_40 (
    .clock(line_40_clock),
    .reset(line_40_reset),
    .valid(line_40_valid)
  );
  GEN_w1_line #(.COVER_INDEX(41)) line_41 (
    .clock(line_41_clock),
    .reset(line_41_reset),
    .valid(line_41_valid)
  );
  GEN_w1_line #(.COVER_INDEX(42)) line_42 (
    .clock(line_42_clock),
    .reset(line_42_reset),
    .valid(line_42_valid)
  );
  GEN_w1_line #(.COVER_INDEX(43)) line_43 (
    .clock(line_43_clock),
    .reset(line_43_reset),
    .valid(line_43_valid)
  );
  GEN_w1_line #(.COVER_INDEX(44)) line_44 (
    .clock(line_44_clock),
    .reset(line_44_reset),
    .valid(line_44_valid)
  );
  assign line_37_clock = clock;
  assign line_37_reset = reset;
  assign line_37_valid = _T_5 ^ line_37_valid_reg;
  assign line_38_clock = clock;
  assign line_38_reset = reset;
  assign line_38_valid = _T_7 ^ line_38_valid_reg;
  assign line_39_clock = clock;
  assign line_39_reset = reset;
  assign line_39_valid = dFirst ^ line_39_valid_reg;
  assign line_40_clock = clock;
  assign line_40_reset = reset;
  assign line_40_valid = aFirst ^ line_40_valid_reg;
  assign line_41_clock = clock;
  assign line_41_reset = reset;
  assign line_41_valid = _T_8 ^ line_41_valid_reg;
  assign line_42_clock = clock;
  assign line_42_reset = reset;
  assign line_42_valid = _T_5 ^ line_42_valid_reg;
  assign line_43_clock = clock;
  assign line_43_reset = reset;
  assign line_43_valid = _T_5 ^ line_43_valid_reg;
  assign line_44_clock = clock;
  assign line_44_reset = reset;
  assign line_44_valid = _T_20 ^ line_44_valid_reg;
  assign auto_in_a_ready = repeater_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Fragmenter.scala 265:25]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Fragmenter.scala 226:36]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[src/main/scala/tilelink/Fragmenter.scala 229:32]
  assign auto_in_d_bits_source = auto_out_d_bits_source[4:3]; // @[src/main/scala/tilelink/Fragmenter.scala 228:47]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Fragmenter.scala 305:15]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Fragmenter.scala 308:25]
  assign auto_out_a_bits_source = {nodeOut_a_bits_source_hi,new_gennum}; // @[src/main/scala/tilelink/Fragmenter.scala 307:33]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_20; // @[src/main/scala/tilelink/Fragmenter.scala 306:49]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/tilelink/Fragmenter.scala 225:35]
  assign repeater_clock = clock;
  assign repeater_reset = reset;
  assign repeater_io_repeat = new_gennum != 2'h0; // @[src/main/scala/tilelink/Fragmenter.scala 304:53]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Fragmenter.scala 191:29]
      acknum <= 2'h0; // @[src/main/scala/tilelink/Fragmenter.scala 191:29]
    end else if (_T_7) begin // @[src/main/scala/tilelink/Fragmenter.scala 210:27]
      if (dFirst) begin // @[src/main/scala/tilelink/Fragmenter.scala 211:24]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[src/main/scala/tilelink/Fragmenter.scala 210:27]
      if (dFirst) begin // @[src/main/scala/tilelink/Fragmenter.scala 212:25]
        dOrig <= dFirst_size; // @[src/main/scala/tilelink/Fragmenter.scala 213:19]
      end
    end
    if (reset) begin // @[src/main/scala/tilelink/Fragmenter.scala 193:30]
      dToggle <= 1'h0; // @[src/main/scala/tilelink/Fragmenter.scala 193:30]
    end else if (_T_7) begin // @[src/main/scala/tilelink/Fragmenter.scala 210:27]
      if (dFirst) begin // @[src/main/scala/tilelink/Fragmenter.scala 212:25]
        dToggle <= auto_out_d_bits_source[2]; // @[src/main/scala/tilelink/Fragmenter.scala 214:21]
      end
    end
    line_37_valid_reg <= _T_5;
    line_38_valid_reg <= _T_7;
    line_39_valid_reg <= dFirst;
    if (reset) begin // @[src/main/scala/tilelink/Fragmenter.scala 293:29]
      gennum <= 2'h0; // @[src/main/scala/tilelink/Fragmenter.scala 293:29]
    end else if (_T_8) begin // @[src/main/scala/tilelink/Fragmenter.scala 302:27]
      gennum <= new_gennum; // @[src/main/scala/tilelink/Fragmenter.scala 302:36]
    end
    if (aFirst) begin // @[src/main/scala/tilelink/Fragmenter.scala 299:54]
      aToggle_r <= dToggle; // @[src/main/scala/tilelink/Fragmenter.scala 299:54]
    end
    line_40_valid_reg <= aFirst;
    line_41_valid_reg <= _T_8;
    line_42_valid_reg <= _T_5;
    line_43_valid_reg <= _T_5;
    line_44_valid_reg <= _T_20;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & ~(_T_9 | repeater_io_deq_bits_mask == 8'hff)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[src/main/scala/tilelink/Fragmenter.scala 314:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_37_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_38_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_39_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  gennum = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  aToggle_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_40_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_41_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_42_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_43_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_44_valid_reg = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/tilelink/Fragmenter.scala 204:16]
    end
    //
    if (_T_5) begin
      assert(1'h1); // @[src/main/scala/tilelink/Fragmenter.scala 311:16]
    end
    //
    if (_T_5) begin
      assert(_T_9 | repeater_io_deq_bits_mask == 8'hff); // @[src/main/scala/tilelink/Fragmenter.scala 314:16]
    end
  end
endmodule
module TLInterconnectCoupler_6(
  input         clock,
  input         reset,
  input         auto_fragmenter_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fragmenter_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_fragmenter_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [4:0]  auto_fragmenter_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_fragmenter_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fragmenter_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_fragmenter_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_fragmenter_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [4:0]  auto_fragmenter_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_fragmenter_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_tl_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_tl_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_in_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  fragmenter_clock; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_reset; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_in_a_ready; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_in_a_valid; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [1:0] fragmenter_auto_in_a_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_in_d_ready; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_in_d_valid; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [1:0] fragmenter_auto_in_d_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_out_a_ready; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_out_a_valid; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [4:0] fragmenter_auto_out_a_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_out_d_ready; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_auto_out_d_valid; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [4:0] fragmenter_auto_out_d_bits_source; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  TLFragmenter fragmenter ( // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data)
  );
  assign auto_fragmenter_out_a_valid = fragmenter_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fragmenter_out_a_bits_size = fragmenter_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fragmenter_out_a_bits_source = fragmenter_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fragmenter_out_a_bits_address = fragmenter_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fragmenter_out_d_ready = fragmenter_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_a_ready = fragmenter_auto_in_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_tl_in_d_valid = fragmenter_auto_in_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_tl_in_d_bits_size = fragmenter_auto_in_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_tl_in_d_bits_source = fragmenter_auto_in_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_tl_in_d_bits_data = fragmenter_auto_in_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign fragmenter_auto_in_a_valid = auto_tl_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_in_a_bits_size = auto_tl_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_in_a_bits_source = auto_tl_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_in_a_bits_address = auto_tl_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_in_a_bits_mask = auto_tl_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_in_d_ready = auto_tl_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign fragmenter_auto_out_a_ready = auto_fragmenter_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign fragmenter_auto_out_d_valid = auto_fragmenter_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign fragmenter_auto_out_d_bits_size = auto_fragmenter_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign fragmenter_auto_out_d_bits_source = auto_fragmenter_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign fragmenter_auto_out_d_bits_data = auto_fragmenter_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
endmodule
module PeripheryBus_1(
  input         auto_coupler_to_bootrom_fragmenter_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bootrom_fragmenter_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_bootrom_fragmenter_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [4:0]  auto_coupler_to_bootrom_fragmenter_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [28:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bootrom_fragmenter_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bootrom_fragmenter_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_bootrom_fragmenter_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [4:0]  auto_coupler_to_bootrom_fragmenter_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_fixedClockNode_out_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_bus_xing_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_bus_xing_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_bus_xing_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_bus_xing_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_bus_xing_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_bus_xing_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_cbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_cbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_1_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_1_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_0_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_0_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  fixer_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_in_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_in_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [1:0] fixer_auto_in_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [28:0] fixer_auto_in_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_in_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_in_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [1:0] fixer_auto_in_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_in_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_out_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [1:0] fixer_auto_out_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [28:0] fixer_auto_out_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  fixer_auto_out_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [2:0] fixer_auto_out_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [1:0] fixer_auto_out_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire [63:0] fixer_auto_out_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
  wire  in_xbar_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_in_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_in_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [28:0] in_xbar_auto_in_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [7:0] in_xbar_auto_in_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_in_d_bits_opcode; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_in_d_bits_param; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_in_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_in_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_d_bits_sink; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_d_bits_denied; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [63:0] in_xbar_auto_in_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_out_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_out_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [28:0] in_xbar_auto_out_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [7:0] in_xbar_auto_out_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_out_d_bits_opcode; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_out_d_bits_param; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [2:0] in_xbar_auto_out_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [1:0] in_xbar_auto_out_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_d_bits_sink; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_d_bits_denied; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire [63:0] in_xbar_auto_out_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  in_xbar_auto_out_d_bits_corrupt; // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
  wire  out_xbar_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_in_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [1:0] out_xbar_auto_in_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [28:0] out_xbar_auto_in_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_in_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_in_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_in_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [1:0] out_xbar_auto_in_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_in_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [1:0] out_xbar_auto_out_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [28:0] out_xbar_auto_out_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [7:0] out_xbar_auto_out_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  out_xbar_auto_out_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [2:0] out_xbar_auto_out_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [1:0] out_xbar_auto_out_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire [63:0] out_xbar_auto_out_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [28:0] buffer_auto_in_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [28:0] buffer_auto_out_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  atomics_clock; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_reset; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_a_ready; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_a_valid; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_in_a_bits_size; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_in_a_bits_source; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [28:0] atomics_auto_in_a_bits_address; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [7:0] atomics_auto_in_a_bits_mask; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_d_ready; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_d_valid; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_in_d_bits_param; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_in_d_bits_size; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_in_d_bits_source; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_d_bits_sink; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_d_bits_denied; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [63:0] atomics_auto_in_d_bits_data; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_a_ready; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_a_valid; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_out_a_bits_size; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_out_a_bits_source; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [28:0] atomics_auto_out_a_bits_address; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [7:0] atomics_auto_out_a_bits_mask; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_d_ready; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_d_valid; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_out_d_bits_param; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [2:0] atomics_auto_out_d_bits_size; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [1:0] atomics_auto_out_d_bits_source; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_d_bits_sink; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_d_bits_denied; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire [63:0] atomics_auto_out_d_bits_data; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  atomics_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
  wire  buffer_1_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_in_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_in_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [28:0] buffer_1_auto_in_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_in_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_in_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_in_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_out_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_out_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [28:0] buffer_1_auto_out_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_1_auto_out_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_1_auto_out_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  coupler_to_bus_named_subsystem_pbus_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_pbus_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_tile_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_tile_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [4:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [28:0] coupler_to_bootrom_auto_fragmenter_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_fragmenter_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [4:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bootrom_auto_fragmenter_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_tl_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_tl_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bootrom_auto_tl_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bootrom_auto_tl_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [28:0] coupler_to_bootrom_auto_tl_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bootrom_auto_tl_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_tl_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bootrom_auto_tl_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bootrom_auto_tl_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_bootrom_auto_tl_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bootrom_auto_tl_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  ClockGroupAggregator_3 subsystem_cbus_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_cbus_1_clock(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock),
    .auto_in_member_subsystem_cbus_1_reset(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset),
    .auto_in_member_subsystem_cbus_0_clock(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock),
    .auto_in_member_subsystem_cbus_0_reset(subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset),
    .auto_out_1_member_subsystem_pbus_0_clock(subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock),
    .auto_out_1_member_subsystem_pbus_0_reset(subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset),
    .auto_out_0_member_subsystem_cbus_0_clock(subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock),
    .auto_out_0_member_subsystem_cbus_0_reset(subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset)
  );
  ClockGroup_3 clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_cbus_0_clock(clockGroup_auto_in_member_subsystem_cbus_0_clock),
    .auto_in_member_subsystem_cbus_0_reset(clockGroup_auto_in_member_subsystem_cbus_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast_3 fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_1_clock(fixedClockNode_auto_out_1_clock),
    .auto_out_1_reset(fixedClockNode_auto_out_1_reset),
    .auto_out_0_clock(fixedClockNode_auto_out_0_clock),
    .auto_out_0_reset(fixedClockNode_auto_out_0_reset)
  );
  BundleBridgeNexus_3 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLFIFOFixer_2 fixer ( // @[src/main/scala/subsystem/PeripheryBus.scala 47:33]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data)
  );
  TLXbar_4 in_xbar ( // @[src/main/scala/subsystem/PeripheryBus.scala 49:29]
    .clock(in_xbar_clock),
    .reset(in_xbar_reset),
    .auto_in_a_ready(in_xbar_auto_in_a_ready),
    .auto_in_a_valid(in_xbar_auto_in_a_valid),
    .auto_in_a_bits_size(in_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(in_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(in_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(in_xbar_auto_in_a_bits_mask),
    .auto_in_d_ready(in_xbar_auto_in_d_ready),
    .auto_in_d_valid(in_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(in_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(in_xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(in_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(in_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(in_xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(in_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(in_xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(in_xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(in_xbar_auto_out_a_ready),
    .auto_out_a_valid(in_xbar_auto_out_a_valid),
    .auto_out_a_bits_size(in_xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(in_xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(in_xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(in_xbar_auto_out_a_bits_mask),
    .auto_out_d_ready(in_xbar_auto_out_d_ready),
    .auto_out_d_valid(in_xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(in_xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(in_xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(in_xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(in_xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(in_xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(in_xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(in_xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(in_xbar_auto_out_d_bits_corrupt)
  );
  TLXbar_5 out_xbar ( // @[src/main/scala/subsystem/PeripheryBus.scala 50:30]
    .clock(out_xbar_clock),
    .reset(out_xbar_reset),
    .auto_in_a_ready(out_xbar_auto_in_a_ready),
    .auto_in_a_valid(out_xbar_auto_in_a_valid),
    .auto_in_a_bits_size(out_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(out_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(out_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(out_xbar_auto_in_a_bits_mask),
    .auto_in_d_ready(out_xbar_auto_in_d_ready),
    .auto_in_d_valid(out_xbar_auto_in_d_valid),
    .auto_in_d_bits_size(out_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(out_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_data(out_xbar_auto_in_d_bits_data),
    .auto_out_a_ready(out_xbar_auto_out_a_ready),
    .auto_out_a_valid(out_xbar_auto_out_a_valid),
    .auto_out_a_bits_size(out_xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(out_xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(out_xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(out_xbar_auto_out_a_bits_mask),
    .auto_out_d_ready(out_xbar_auto_out_d_ready),
    .auto_out_d_valid(out_xbar_auto_out_d_valid),
    .auto_out_d_bits_size(out_xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(out_xbar_auto_out_d_bits_source),
    .auto_out_d_bits_data(out_xbar_auto_out_d_bits_data)
  );
  TLBuffer_3 buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLAtomicAutomata_1 atomics ( // @[src/main/scala/tilelink/AtomicAutomata.scala 285:29]
    .clock(atomics_clock),
    .reset(atomics_reset),
    .auto_in_a_ready(atomics_auto_in_a_ready),
    .auto_in_a_valid(atomics_auto_in_a_valid),
    .auto_in_a_bits_size(atomics_auto_in_a_bits_size),
    .auto_in_a_bits_source(atomics_auto_in_a_bits_source),
    .auto_in_a_bits_address(atomics_auto_in_a_bits_address),
    .auto_in_a_bits_mask(atomics_auto_in_a_bits_mask),
    .auto_in_d_ready(atomics_auto_in_d_ready),
    .auto_in_d_valid(atomics_auto_in_d_valid),
    .auto_in_d_bits_opcode(atomics_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(atomics_auto_in_d_bits_param),
    .auto_in_d_bits_size(atomics_auto_in_d_bits_size),
    .auto_in_d_bits_source(atomics_auto_in_d_bits_source),
    .auto_in_d_bits_sink(atomics_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(atomics_auto_in_d_bits_denied),
    .auto_in_d_bits_data(atomics_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(atomics_auto_in_d_bits_corrupt),
    .auto_out_a_ready(atomics_auto_out_a_ready),
    .auto_out_a_valid(atomics_auto_out_a_valid),
    .auto_out_a_bits_size(atomics_auto_out_a_bits_size),
    .auto_out_a_bits_source(atomics_auto_out_a_bits_source),
    .auto_out_a_bits_address(atomics_auto_out_a_bits_address),
    .auto_out_a_bits_mask(atomics_auto_out_a_bits_mask),
    .auto_out_d_ready(atomics_auto_out_d_ready),
    .auto_out_d_valid(atomics_auto_out_d_valid),
    .auto_out_d_bits_opcode(atomics_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(atomics_auto_out_d_bits_param),
    .auto_out_d_bits_size(atomics_auto_out_d_bits_size),
    .auto_out_d_bits_source(atomics_auto_out_d_bits_source),
    .auto_out_d_bits_sink(atomics_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(atomics_auto_out_d_bits_denied),
    .auto_out_d_bits_data(atomics_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(atomics_auto_out_d_bits_corrupt)
  );
  TLBuffer_4 buffer_1 ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_1_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  TLInterconnectCoupler_4 coupler_to_bus_named_subsystem_pbus ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_bus_named_subsystem_pbus_clock),
    .reset(coupler_to_bus_named_subsystem_pbus_reset)
  );
  TLInterconnectCoupler_5 coupler_to_tile ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_tile_clock),
    .reset(coupler_to_tile_reset)
  );
  TLInterconnectCoupler_6 coupler_to_bootrom ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_bootrom_clock),
    .reset(coupler_to_bootrom_reset),
    .auto_fragmenter_out_a_ready(coupler_to_bootrom_auto_fragmenter_out_a_ready),
    .auto_fragmenter_out_a_valid(coupler_to_bootrom_auto_fragmenter_out_a_valid),
    .auto_fragmenter_out_a_bits_size(coupler_to_bootrom_auto_fragmenter_out_a_bits_size),
    .auto_fragmenter_out_a_bits_source(coupler_to_bootrom_auto_fragmenter_out_a_bits_source),
    .auto_fragmenter_out_a_bits_address(coupler_to_bootrom_auto_fragmenter_out_a_bits_address),
    .auto_fragmenter_out_d_ready(coupler_to_bootrom_auto_fragmenter_out_d_ready),
    .auto_fragmenter_out_d_valid(coupler_to_bootrom_auto_fragmenter_out_d_valid),
    .auto_fragmenter_out_d_bits_size(coupler_to_bootrom_auto_fragmenter_out_d_bits_size),
    .auto_fragmenter_out_d_bits_source(coupler_to_bootrom_auto_fragmenter_out_d_bits_source),
    .auto_fragmenter_out_d_bits_data(coupler_to_bootrom_auto_fragmenter_out_d_bits_data),
    .auto_tl_in_a_ready(coupler_to_bootrom_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_bootrom_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_size(coupler_to_bootrom_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_bootrom_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_bootrom_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_bootrom_auto_tl_in_a_bits_mask),
    .auto_tl_in_d_ready(coupler_to_bootrom_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_bootrom_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_size(coupler_to_bootrom_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_bootrom_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_data(coupler_to_bootrom_auto_tl_in_d_bits_data)
  );
  assign auto_coupler_to_bootrom_fragmenter_out_a_valid = coupler_to_bootrom_auto_fragmenter_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_size = coupler_to_bootrom_auto_fragmenter_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_source = coupler_to_bootrom_auto_fragmenter_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bootrom_fragmenter_out_a_bits_address = coupler_to_bootrom_auto_fragmenter_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bootrom_fragmenter_out_d_ready = coupler_to_bootrom_auto_fragmenter_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_clock = fixedClockNode_auto_out_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_fixedClockNode_out_reset = fixedClockNode_auto_out_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock =
    subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset =
    subsystem_cbus_clock_groups_auto_out_1_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_bus_xing_in_a_ready = buffer_1_auto_in_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_valid = buffer_1_auto_in_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_opcode = buffer_1_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_param = buffer_1_auto_in_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_size = buffer_1_auto_in_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_source = buffer_1_auto_in_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_sink = buffer_1_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_denied = buffer_1_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_data = buffer_1_auto_in_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_corrupt = buffer_1_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_clock =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_1_reset =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_clock =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_cbus_clock_groups_auto_in_member_subsystem_cbus_0_reset =
    auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_cbus_0_clock =
    subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_cbus_0_reset =
    subsystem_cbus_clock_groups_auto_out_0_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_valid = buffer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_d_ready = buffer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_a_ready = out_xbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_auto_out_d_valid = out_xbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_auto_out_d_bits_size = out_xbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_auto_out_d_bits_source = out_xbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_auto_out_d_bits_data = out_xbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_a_valid = buffer_1_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_in_d_ready = buffer_1_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign in_xbar_auto_out_a_ready = atomics_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_valid = atomics_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_opcode = atomics_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_param = atomics_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_size = atomics_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_source = atomics_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_sink = atomics_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_denied = atomics_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_data = atomics_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign in_xbar_auto_out_d_bits_corrupt = atomics_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign out_xbar_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign out_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_out_a_ready = coupler_to_bootrom_auto_tl_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_out_d_valid = coupler_to_bootrom_auto_tl_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_out_d_bits_size = coupler_to_bootrom_auto_tl_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_out_d_bits_source = coupler_to_bootrom_auto_tl_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign out_xbar_auto_out_d_bits_data = coupler_to_bootrom_auto_tl_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_valid = atomics_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_size = atomics_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_source = atomics_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_address = atomics_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_mask = atomics_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_d_ready = atomics_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_a_ready = fixer_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_valid = fixer_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_in_a_valid = in_xbar_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_in_a_bits_size = in_xbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_in_a_bits_source = in_xbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_in_a_bits_address = in_xbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_in_a_bits_mask = in_xbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_in_d_ready = in_xbar_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign atomics_auto_out_a_ready = buffer_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_valid = buffer_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign atomics_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_in_a_valid = auto_bus_xing_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_in_d_ready = auto_bus_xing_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_auto_out_a_ready = in_xbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_valid = in_xbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_opcode = in_xbar_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_param = in_xbar_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_size = in_xbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_source = in_xbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_sink = in_xbar_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_denied = in_xbar_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_data = in_xbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_1_auto_out_d_bits_corrupt = in_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_pbus_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_pbus_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_tile_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_tile_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bootrom_clock = fixedClockNode_auto_out_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bootrom_reset = fixedClockNode_auto_out_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bootrom_auto_fragmenter_out_a_ready = auto_coupler_to_bootrom_fragmenter_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_valid = auto_coupler_to_bootrom_fragmenter_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_size = auto_coupler_to_bootrom_fragmenter_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_source = auto_coupler_to_bootrom_fragmenter_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bootrom_auto_fragmenter_out_d_bits_data = auto_coupler_to_bootrom_fragmenter_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bootrom_auto_tl_in_a_valid = out_xbar_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bootrom_auto_tl_in_a_bits_size = out_xbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bootrom_auto_tl_in_a_bits_source = out_xbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bootrom_auto_tl_in_a_bits_address = out_xbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bootrom_auto_tl_in_a_bits_mask = out_xbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bootrom_auto_tl_in_d_ready = out_xbar_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
endmodule
module ClockGroupAggregator_4(
  input   auto_in_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_mbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_member_subsystem_mbus_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_member_subsystem_mbus_0_clock = auto_in_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_member_subsystem_mbus_0_reset = auto_in_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup_4(
  input   auto_in_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_mbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_4(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_4(
  input   clock,
  input   reset
);
endmodule
module TLXbar_6(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLFIFOFixer_3(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  wire  _a_first_T = auto_out_a_ready & auto_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _a_first_beats1_decode_T_1 = 12'h1f << auto_in_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  reg [1:0] a_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] a_first_counter1 = a_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_45_clock;
  wire  line_45_reset;
  wire  line_45_valid;
  reg  line_45_valid_reg;
  wire  _d_first_T = auto_in_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _d_first_beats1_decode_T_1 = 12'h1f << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  d_first_beats1_opdata = auto_out_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  reg [1:0] d_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] d_first_counter1 = d_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  d_first_first = d_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_46_clock;
  wire  line_46_reset;
  wire  line_46_valid;
  reg  line_46_valid_reg;
  wire  d_first = d_first_first & auto_out_d_bits_opcode != 3'h6; // @[src/main/scala/tilelink/FIFOFixer.scala 69:42]
  wire  _T_1 = a_first & _a_first_T; // @[src/main/scala/tilelink/FIFOFixer.scala 74:21]
  wire  line_47_clock;
  wire  line_47_reset;
  wire  line_47_valid;
  reg  line_47_valid_reg;
  wire  line_48_clock;
  wire  line_48_reset;
  wire  line_48_valid;
  reg  line_48_valid_reg;
  wire  line_49_clock;
  wire  line_49_reset;
  wire  line_49_valid;
  reg  line_49_valid_reg;
  wire  line_50_clock;
  wire  line_50_reset;
  wire  line_50_valid;
  reg  line_50_valid_reg;
  wire  line_51_clock;
  wire  line_51_reset;
  wire  line_51_valid;
  reg  line_51_valid_reg;
  wire  line_52_clock;
  wire  line_52_reset;
  wire  line_52_valid;
  reg  line_52_valid_reg;
  wire  line_53_clock;
  wire  line_53_reset;
  wire  line_53_valid;
  reg  line_53_valid_reg;
  wire  line_54_clock;
  wire  line_54_reset;
  wire  line_54_valid;
  reg  line_54_valid_reg;
  wire  line_55_clock;
  wire  line_55_reset;
  wire  line_55_valid;
  reg  line_55_valid_reg;
  wire  line_56_clock;
  wire  line_56_reset;
  wire  line_56_valid;
  reg  line_56_valid_reg;
  wire  line_57_clock;
  wire  line_57_reset;
  wire  line_57_valid;
  reg  line_57_valid_reg;
  wire  line_58_clock;
  wire  line_58_reset;
  wire  line_58_valid;
  reg  line_58_valid_reg;
  wire  line_59_clock;
  wire  line_59_reset;
  wire  line_59_valid;
  reg  line_59_valid_reg;
  wire  line_60_clock;
  wire  line_60_reset;
  wire  line_60_valid;
  reg  line_60_valid_reg;
  wire  line_61_clock;
  wire  line_61_reset;
  wire  line_61_valid;
  reg  line_61_valid_reg;
  wire  line_62_clock;
  wire  line_62_reset;
  wire  line_62_valid;
  reg  line_62_valid_reg;
  wire  line_63_clock;
  wire  line_63_reset;
  wire  line_63_valid;
  reg  line_63_valid_reg;
  wire  _T_3 = d_first & _d_first_T; // @[src/main/scala/tilelink/FIFOFixer.scala 75:21]
  wire  line_64_clock;
  wire  line_64_reset;
  wire  line_64_valid;
  reg  line_64_valid_reg;
  wire  line_65_clock;
  wire  line_65_reset;
  wire  line_65_valid;
  reg  line_65_valid_reg;
  wire  line_66_clock;
  wire  line_66_reset;
  wire  line_66_valid;
  reg  line_66_valid_reg;
  wire  line_67_clock;
  wire  line_67_reset;
  wire  line_67_valid;
  reg  line_67_valid_reg;
  wire  line_68_clock;
  wire  line_68_reset;
  wire  line_68_valid;
  reg  line_68_valid_reg;
  wire  line_69_clock;
  wire  line_69_reset;
  wire  line_69_valid;
  reg  line_69_valid_reg;
  wire  line_70_clock;
  wire  line_70_reset;
  wire  line_70_valid;
  reg  line_70_valid_reg;
  wire  line_71_clock;
  wire  line_71_reset;
  wire  line_71_valid;
  reg  line_71_valid_reg;
  wire  line_72_clock;
  wire  line_72_reset;
  wire  line_72_valid;
  reg  line_72_valid_reg;
  wire  line_73_clock;
  wire  line_73_reset;
  wire  line_73_valid;
  reg  line_73_valid_reg;
  wire  line_74_clock;
  wire  line_74_reset;
  wire  line_74_valid;
  reg  line_74_valid_reg;
  wire  line_75_clock;
  wire  line_75_reset;
  wire  line_75_valid;
  reg  line_75_valid_reg;
  wire  line_76_clock;
  wire  line_76_reset;
  wire  line_76_valid;
  reg  line_76_valid_reg;
  wire  line_77_clock;
  wire  line_77_reset;
  wire  line_77_valid;
  reg  line_77_valid_reg;
  wire  line_78_clock;
  wire  line_78_reset;
  wire  line_78_valid;
  reg  line_78_valid_reg;
  wire  line_79_clock;
  wire  line_79_reset;
  wire  line_79_valid;
  reg  line_79_valid_reg;
  wire  line_80_clock;
  wire  line_80_reset;
  wire  line_80_valid;
  reg  line_80_valid_reg;
  wire  line_81_clock;
  wire  line_81_reset;
  wire  line_81_valid;
  reg  line_81_valid_reg;
  wire  line_82_clock;
  wire  line_82_reset;
  wire  line_82_valid;
  reg  line_82_valid_reg;
  GEN_w1_line #(.COVER_INDEX(45)) line_45 (
    .clock(line_45_clock),
    .reset(line_45_reset),
    .valid(line_45_valid)
  );
  GEN_w1_line #(.COVER_INDEX(46)) line_46 (
    .clock(line_46_clock),
    .reset(line_46_reset),
    .valid(line_46_valid)
  );
  GEN_w1_line #(.COVER_INDEX(47)) line_47 (
    .clock(line_47_clock),
    .reset(line_47_reset),
    .valid(line_47_valid)
  );
  GEN_w1_line #(.COVER_INDEX(48)) line_48 (
    .clock(line_48_clock),
    .reset(line_48_reset),
    .valid(line_48_valid)
  );
  GEN_w1_line #(.COVER_INDEX(49)) line_49 (
    .clock(line_49_clock),
    .reset(line_49_reset),
    .valid(line_49_valid)
  );
  GEN_w1_line #(.COVER_INDEX(50)) line_50 (
    .clock(line_50_clock),
    .reset(line_50_reset),
    .valid(line_50_valid)
  );
  GEN_w1_line #(.COVER_INDEX(51)) line_51 (
    .clock(line_51_clock),
    .reset(line_51_reset),
    .valid(line_51_valid)
  );
  GEN_w1_line #(.COVER_INDEX(52)) line_52 (
    .clock(line_52_clock),
    .reset(line_52_reset),
    .valid(line_52_valid)
  );
  GEN_w1_line #(.COVER_INDEX(53)) line_53 (
    .clock(line_53_clock),
    .reset(line_53_reset),
    .valid(line_53_valid)
  );
  GEN_w1_line #(.COVER_INDEX(54)) line_54 (
    .clock(line_54_clock),
    .reset(line_54_reset),
    .valid(line_54_valid)
  );
  GEN_w1_line #(.COVER_INDEX(55)) line_55 (
    .clock(line_55_clock),
    .reset(line_55_reset),
    .valid(line_55_valid)
  );
  GEN_w1_line #(.COVER_INDEX(56)) line_56 (
    .clock(line_56_clock),
    .reset(line_56_reset),
    .valid(line_56_valid)
  );
  GEN_w1_line #(.COVER_INDEX(57)) line_57 (
    .clock(line_57_clock),
    .reset(line_57_reset),
    .valid(line_57_valid)
  );
  GEN_w1_line #(.COVER_INDEX(58)) line_58 (
    .clock(line_58_clock),
    .reset(line_58_reset),
    .valid(line_58_valid)
  );
  GEN_w1_line #(.COVER_INDEX(59)) line_59 (
    .clock(line_59_clock),
    .reset(line_59_reset),
    .valid(line_59_valid)
  );
  GEN_w1_line #(.COVER_INDEX(60)) line_60 (
    .clock(line_60_clock),
    .reset(line_60_reset),
    .valid(line_60_valid)
  );
  GEN_w1_line #(.COVER_INDEX(61)) line_61 (
    .clock(line_61_clock),
    .reset(line_61_reset),
    .valid(line_61_valid)
  );
  GEN_w1_line #(.COVER_INDEX(62)) line_62 (
    .clock(line_62_clock),
    .reset(line_62_reset),
    .valid(line_62_valid)
  );
  GEN_w1_line #(.COVER_INDEX(63)) line_63 (
    .clock(line_63_clock),
    .reset(line_63_reset),
    .valid(line_63_valid)
  );
  GEN_w1_line #(.COVER_INDEX(64)) line_64 (
    .clock(line_64_clock),
    .reset(line_64_reset),
    .valid(line_64_valid)
  );
  GEN_w1_line #(.COVER_INDEX(65)) line_65 (
    .clock(line_65_clock),
    .reset(line_65_reset),
    .valid(line_65_valid)
  );
  GEN_w1_line #(.COVER_INDEX(66)) line_66 (
    .clock(line_66_clock),
    .reset(line_66_reset),
    .valid(line_66_valid)
  );
  GEN_w1_line #(.COVER_INDEX(67)) line_67 (
    .clock(line_67_clock),
    .reset(line_67_reset),
    .valid(line_67_valid)
  );
  GEN_w1_line #(.COVER_INDEX(68)) line_68 (
    .clock(line_68_clock),
    .reset(line_68_reset),
    .valid(line_68_valid)
  );
  GEN_w1_line #(.COVER_INDEX(69)) line_69 (
    .clock(line_69_clock),
    .reset(line_69_reset),
    .valid(line_69_valid)
  );
  GEN_w1_line #(.COVER_INDEX(70)) line_70 (
    .clock(line_70_clock),
    .reset(line_70_reset),
    .valid(line_70_valid)
  );
  GEN_w1_line #(.COVER_INDEX(71)) line_71 (
    .clock(line_71_clock),
    .reset(line_71_reset),
    .valid(line_71_valid)
  );
  GEN_w1_line #(.COVER_INDEX(72)) line_72 (
    .clock(line_72_clock),
    .reset(line_72_reset),
    .valid(line_72_valid)
  );
  GEN_w1_line #(.COVER_INDEX(73)) line_73 (
    .clock(line_73_clock),
    .reset(line_73_reset),
    .valid(line_73_valid)
  );
  GEN_w1_line #(.COVER_INDEX(74)) line_74 (
    .clock(line_74_clock),
    .reset(line_74_reset),
    .valid(line_74_valid)
  );
  GEN_w1_line #(.COVER_INDEX(75)) line_75 (
    .clock(line_75_clock),
    .reset(line_75_reset),
    .valid(line_75_valid)
  );
  GEN_w1_line #(.COVER_INDEX(76)) line_76 (
    .clock(line_76_clock),
    .reset(line_76_reset),
    .valid(line_76_valid)
  );
  GEN_w1_line #(.COVER_INDEX(77)) line_77 (
    .clock(line_77_clock),
    .reset(line_77_reset),
    .valid(line_77_valid)
  );
  GEN_w1_line #(.COVER_INDEX(78)) line_78 (
    .clock(line_78_clock),
    .reset(line_78_reset),
    .valid(line_78_valid)
  );
  GEN_w1_line #(.COVER_INDEX(79)) line_79 (
    .clock(line_79_clock),
    .reset(line_79_reset),
    .valid(line_79_valid)
  );
  GEN_w1_line #(.COVER_INDEX(80)) line_80 (
    .clock(line_80_clock),
    .reset(line_80_reset),
    .valid(line_80_valid)
  );
  GEN_w1_line #(.COVER_INDEX(81)) line_81 (
    .clock(line_81_clock),
    .reset(line_81_reset),
    .valid(line_81_valid)
  );
  GEN_w1_line #(.COVER_INDEX(82)) line_82 (
    .clock(line_82_clock),
    .reset(line_82_reset),
    .valid(line_82_valid)
  );
  assign line_45_clock = clock;
  assign line_45_reset = reset;
  assign line_45_valid = _a_first_T ^ line_45_valid_reg;
  assign line_46_clock = clock;
  assign line_46_reset = reset;
  assign line_46_valid = _d_first_T ^ line_46_valid_reg;
  assign line_47_clock = clock;
  assign line_47_reset = reset;
  assign line_47_valid = _T_1 ^ line_47_valid_reg;
  assign line_48_clock = clock;
  assign line_48_reset = reset;
  assign line_48_valid = 4'h0 == auto_in_a_bits_source ^ line_48_valid_reg;
  assign line_49_clock = clock;
  assign line_49_reset = reset;
  assign line_49_valid = 4'h1 == auto_in_a_bits_source ^ line_49_valid_reg;
  assign line_50_clock = clock;
  assign line_50_reset = reset;
  assign line_50_valid = 4'h2 == auto_in_a_bits_source ^ line_50_valid_reg;
  assign line_51_clock = clock;
  assign line_51_reset = reset;
  assign line_51_valid = 4'h3 == auto_in_a_bits_source ^ line_51_valid_reg;
  assign line_52_clock = clock;
  assign line_52_reset = reset;
  assign line_52_valid = 4'h4 == auto_in_a_bits_source ^ line_52_valid_reg;
  assign line_53_clock = clock;
  assign line_53_reset = reset;
  assign line_53_valid = 4'h5 == auto_in_a_bits_source ^ line_53_valid_reg;
  assign line_54_clock = clock;
  assign line_54_reset = reset;
  assign line_54_valid = 4'h6 == auto_in_a_bits_source ^ line_54_valid_reg;
  assign line_55_clock = clock;
  assign line_55_reset = reset;
  assign line_55_valid = 4'h7 == auto_in_a_bits_source ^ line_55_valid_reg;
  assign line_56_clock = clock;
  assign line_56_reset = reset;
  assign line_56_valid = 4'h8 == auto_in_a_bits_source ^ line_56_valid_reg;
  assign line_57_clock = clock;
  assign line_57_reset = reset;
  assign line_57_valid = 4'h9 == auto_in_a_bits_source ^ line_57_valid_reg;
  assign line_58_clock = clock;
  assign line_58_reset = reset;
  assign line_58_valid = 4'ha == auto_in_a_bits_source ^ line_58_valid_reg;
  assign line_59_clock = clock;
  assign line_59_reset = reset;
  assign line_59_valid = 4'hb == auto_in_a_bits_source ^ line_59_valid_reg;
  assign line_60_clock = clock;
  assign line_60_reset = reset;
  assign line_60_valid = 4'hc == auto_in_a_bits_source ^ line_60_valid_reg;
  assign line_61_clock = clock;
  assign line_61_reset = reset;
  assign line_61_valid = 4'hd == auto_in_a_bits_source ^ line_61_valid_reg;
  assign line_62_clock = clock;
  assign line_62_reset = reset;
  assign line_62_valid = 4'he == auto_in_a_bits_source ^ line_62_valid_reg;
  assign line_63_clock = clock;
  assign line_63_reset = reset;
  assign line_63_valid = 4'hf == auto_in_a_bits_source ^ line_63_valid_reg;
  assign line_64_clock = clock;
  assign line_64_reset = reset;
  assign line_64_valid = _T_3 ^ line_64_valid_reg;
  assign line_65_clock = clock;
  assign line_65_reset = reset;
  assign line_65_valid = 4'h0 == auto_out_d_bits_source ^ line_65_valid_reg;
  assign line_66_clock = clock;
  assign line_66_reset = reset;
  assign line_66_valid = 4'h1 == auto_out_d_bits_source ^ line_66_valid_reg;
  assign line_67_clock = clock;
  assign line_67_reset = reset;
  assign line_67_valid = 4'h2 == auto_out_d_bits_source ^ line_67_valid_reg;
  assign line_68_clock = clock;
  assign line_68_reset = reset;
  assign line_68_valid = 4'h3 == auto_out_d_bits_source ^ line_68_valid_reg;
  assign line_69_clock = clock;
  assign line_69_reset = reset;
  assign line_69_valid = 4'h4 == auto_out_d_bits_source ^ line_69_valid_reg;
  assign line_70_clock = clock;
  assign line_70_reset = reset;
  assign line_70_valid = 4'h5 == auto_out_d_bits_source ^ line_70_valid_reg;
  assign line_71_clock = clock;
  assign line_71_reset = reset;
  assign line_71_valid = 4'h6 == auto_out_d_bits_source ^ line_71_valid_reg;
  assign line_72_clock = clock;
  assign line_72_reset = reset;
  assign line_72_valid = 4'h7 == auto_out_d_bits_source ^ line_72_valid_reg;
  assign line_73_clock = clock;
  assign line_73_reset = reset;
  assign line_73_valid = 4'h8 == auto_out_d_bits_source ^ line_73_valid_reg;
  assign line_74_clock = clock;
  assign line_74_reset = reset;
  assign line_74_valid = 4'h9 == auto_out_d_bits_source ^ line_74_valid_reg;
  assign line_75_clock = clock;
  assign line_75_reset = reset;
  assign line_75_valid = 4'ha == auto_out_d_bits_source ^ line_75_valid_reg;
  assign line_76_clock = clock;
  assign line_76_reset = reset;
  assign line_76_valid = 4'hb == auto_out_d_bits_source ^ line_76_valid_reg;
  assign line_77_clock = clock;
  assign line_77_reset = reset;
  assign line_77_valid = 4'hc == auto_out_d_bits_source ^ line_77_valid_reg;
  assign line_78_clock = clock;
  assign line_78_reset = reset;
  assign line_78_valid = 4'hd == auto_out_d_bits_source ^ line_78_valid_reg;
  assign line_79_clock = clock;
  assign line_79_reset = reset;
  assign line_79_valid = 4'he == auto_out_d_bits_source ^ line_79_valid_reg;
  assign line_80_clock = clock;
  assign line_80_reset = reset;
  assign line_80_valid = 4'hf == auto_out_d_bits_source ^ line_80_valid_reg;
  assign line_81_clock = clock;
  assign line_81_reset = reset;
  assign line_81_valid = _T_1 ^ line_81_valid_reg;
  assign line_82_clock = clock;
  assign line_82_reset = reset;
  assign line_82_valid = _T_3 ^ line_82_valid_reg;
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 90:33]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 89:33]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      a_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_a_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (a_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (a_first_beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 2'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    line_45_valid_reg <= _a_first_T;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      d_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_d_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (d_first_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (d_first_beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 2'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    line_46_valid_reg <= _d_first_T;
    line_47_valid_reg <= _T_1;
    line_48_valid_reg <= 4'h0 == auto_in_a_bits_source;
    line_49_valid_reg <= 4'h1 == auto_in_a_bits_source;
    line_50_valid_reg <= 4'h2 == auto_in_a_bits_source;
    line_51_valid_reg <= 4'h3 == auto_in_a_bits_source;
    line_52_valid_reg <= 4'h4 == auto_in_a_bits_source;
    line_53_valid_reg <= 4'h5 == auto_in_a_bits_source;
    line_54_valid_reg <= 4'h6 == auto_in_a_bits_source;
    line_55_valid_reg <= 4'h7 == auto_in_a_bits_source;
    line_56_valid_reg <= 4'h8 == auto_in_a_bits_source;
    line_57_valid_reg <= 4'h9 == auto_in_a_bits_source;
    line_58_valid_reg <= 4'ha == auto_in_a_bits_source;
    line_59_valid_reg <= 4'hb == auto_in_a_bits_source;
    line_60_valid_reg <= 4'hc == auto_in_a_bits_source;
    line_61_valid_reg <= 4'hd == auto_in_a_bits_source;
    line_62_valid_reg <= 4'he == auto_in_a_bits_source;
    line_63_valid_reg <= 4'hf == auto_in_a_bits_source;
    line_64_valid_reg <= _T_3;
    line_65_valid_reg <= 4'h0 == auto_out_d_bits_source;
    line_66_valid_reg <= 4'h1 == auto_out_d_bits_source;
    line_67_valid_reg <= 4'h2 == auto_out_d_bits_source;
    line_68_valid_reg <= 4'h3 == auto_out_d_bits_source;
    line_69_valid_reg <= 4'h4 == auto_out_d_bits_source;
    line_70_valid_reg <= 4'h5 == auto_out_d_bits_source;
    line_71_valid_reg <= 4'h6 == auto_out_d_bits_source;
    line_72_valid_reg <= 4'h7 == auto_out_d_bits_source;
    line_73_valid_reg <= 4'h8 == auto_out_d_bits_source;
    line_74_valid_reg <= 4'h9 == auto_out_d_bits_source;
    line_75_valid_reg <= 4'ha == auto_out_d_bits_source;
    line_76_valid_reg <= 4'hb == auto_out_d_bits_source;
    line_77_valid_reg <= 4'hc == auto_out_d_bits_source;
    line_78_valid_reg <= 4'hd == auto_out_d_bits_source;
    line_79_valid_reg <= 4'he == auto_out_d_bits_source;
    line_80_valid_reg <= 4'hf == auto_out_d_bits_source;
    line_81_valid_reg <= _T_1;
    line_82_valid_reg <= _T_3;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_45_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  d_first_counter = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  line_46_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_47_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_48_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_49_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_50_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_51_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_52_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_53_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_54_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_55_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_56_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_57_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_58_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_59_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_60_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_61_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_62_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_63_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_64_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_65_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_66_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_67_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_68_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_69_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_70_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_71_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_72_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_73_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_74_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_75_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_76_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_77_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_78_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_79_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_80_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_81_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_82_valid_reg = _RAND_39[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ProbePicker(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLBuffer_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLXbar_7(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module Queue_2(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_83_clock;
  wire  line_83_reset;
  wire  line_83_valid;
  reg  line_83_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_84_clock;
  wire  line_84_reset;
  wire  line_84_valid;
  reg  line_84_valid_reg;
  GEN_w1_line #(.COVER_INDEX(83)) line_83 (
    .clock(line_83_clock),
    .reset(line_83_reset),
    .valid(line_83_valid)
  );
  GEN_w1_line #(.COVER_INDEX(84)) line_84 (
    .clock(line_84_clock),
    .reset(line_84_reset),
    .valid(line_84_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_83_clock = clock;
  assign line_83_reset = reset;
  assign line_83_valid = do_enq ^ line_83_valid_reg;
  assign line_84_clock = clock;
  assign line_84_reset = reset;
  assign line_84_valid = _T ^ line_84_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_83_valid_reg <= do_enq;
    line_84_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_83_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_84_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_85_clock;
  wire  line_85_reset;
  wire  line_85_valid;
  reg  line_85_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_86_clock;
  wire  line_86_reset;
  wire  line_86_valid;
  reg  line_86_valid_reg;
  GEN_w1_line #(.COVER_INDEX(85)) line_85 (
    .clock(line_85_clock),
    .reset(line_85_reset),
    .valid(line_85_valid)
  );
  GEN_w1_line #(.COVER_INDEX(86)) line_86 (
    .clock(line_86_clock),
    .reset(line_86_reset),
    .valid(line_86_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_85_clock = clock;
  assign line_85_reset = reset;
  assign line_85_valid = do_enq ^ line_85_valid_reg;
  assign line_86_clock = clock;
  assign line_86_reset = reset;
  assign line_86_valid = _T ^ line_86_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_85_valid_reg <= do_enq;
    line_86_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_85_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_86_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_87_clock;
  wire  line_87_reset;
  wire  line_87_valid;
  reg  line_87_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_88_clock;
  wire  line_88_reset;
  wire  line_88_valid;
  reg  line_88_valid_reg;
  GEN_w1_line #(.COVER_INDEX(87)) line_87 (
    .clock(line_87_clock),
    .reset(line_87_reset),
    .valid(line_87_valid)
  );
  GEN_w1_line #(.COVER_INDEX(88)) line_88 (
    .clock(line_88_clock),
    .reset(line_88_reset),
    .valid(line_88_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_87_clock = clock;
  assign line_87_reset = reset;
  assign line_87_valid = do_enq ^ line_87_valid_reg;
  assign line_88_clock = clock;
  assign line_88_reset = reset;
  assign line_88_valid = _T ^ line_88_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_87_valid_reg <= do_enq;
    line_88_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_87_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_88_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_5(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_89_clock;
  wire  line_89_reset;
  wire  line_89_valid;
  reg  line_89_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_90_clock;
  wire  line_90_reset;
  wire  line_90_valid;
  reg  line_90_valid_reg;
  GEN_w1_line #(.COVER_INDEX(89)) line_89 (
    .clock(line_89_clock),
    .reset(line_89_reset),
    .valid(line_89_valid)
  );
  GEN_w1_line #(.COVER_INDEX(90)) line_90 (
    .clock(line_90_clock),
    .reset(line_90_reset),
    .valid(line_90_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_89_clock = clock;
  assign line_89_reset = reset;
  assign line_89_valid = do_enq ^ line_89_valid_reg;
  assign line_90_clock = clock;
  assign line_90_reset = reset;
  assign line_90_valid = _T ^ line_90_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_89_valid_reg <= do_enq;
    line_90_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_89_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_90_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_91_clock;
  wire  line_91_reset;
  wire  line_91_valid;
  reg  line_91_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_92_clock;
  wire  line_92_reset;
  wire  line_92_valid;
  reg  line_92_valid_reg;
  GEN_w1_line #(.COVER_INDEX(91)) line_91 (
    .clock(line_91_clock),
    .reset(line_91_reset),
    .valid(line_91_valid)
  );
  GEN_w1_line #(.COVER_INDEX(92)) line_92 (
    .clock(line_92_clock),
    .reset(line_92_reset),
    .valid(line_92_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_91_clock = clock;
  assign line_91_reset = reset;
  assign line_91_valid = do_enq ^ line_91_valid_reg;
  assign line_92_clock = clock;
  assign line_92_reset = reset;
  assign line_92_valid = _T ^ line_92_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_91_valid_reg <= do_enq;
    line_92_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_91_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_92_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_93_clock;
  wire  line_93_reset;
  wire  line_93_valid;
  reg  line_93_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_94_clock;
  wire  line_94_reset;
  wire  line_94_valid;
  reg  line_94_valid_reg;
  GEN_w1_line #(.COVER_INDEX(93)) line_93 (
    .clock(line_93_clock),
    .reset(line_93_reset),
    .valid(line_93_valid)
  );
  GEN_w1_line #(.COVER_INDEX(94)) line_94 (
    .clock(line_94_clock),
    .reset(line_94_reset),
    .valid(line_94_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_93_clock = clock;
  assign line_93_reset = reset;
  assign line_93_valid = do_enq ^ line_93_valid_reg;
  assign line_94_clock = clock;
  assign line_94_reset = reset;
  assign line_94_valid = _T ^ line_94_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_93_valid_reg <= do_enq;
    line_94_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_93_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_94_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_8(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_95_clock;
  wire  line_95_reset;
  wire  line_95_valid;
  reg  line_95_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_96_clock;
  wire  line_96_reset;
  wire  line_96_valid;
  reg  line_96_valid_reg;
  GEN_w1_line #(.COVER_INDEX(95)) line_95 (
    .clock(line_95_clock),
    .reset(line_95_reset),
    .valid(line_95_valid)
  );
  GEN_w1_line #(.COVER_INDEX(96)) line_96 (
    .clock(line_96_clock),
    .reset(line_96_reset),
    .valid(line_96_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_95_clock = clock;
  assign line_95_reset = reset;
  assign line_95_valid = do_enq ^ line_95_valid_reg;
  assign line_96_clock = clock;
  assign line_96_reset = reset;
  assign line_96_valid = _T ^ line_96_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_95_valid_reg <= do_enq;
    line_96_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_95_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_96_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_9(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_97_clock;
  wire  line_97_reset;
  wire  line_97_valid;
  reg  line_97_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_98_clock;
  wire  line_98_reset;
  wire  line_98_valid;
  reg  line_98_valid_reg;
  GEN_w1_line #(.COVER_INDEX(97)) line_97 (
    .clock(line_97_clock),
    .reset(line_97_reset),
    .valid(line_97_valid)
  );
  GEN_w1_line #(.COVER_INDEX(98)) line_98 (
    .clock(line_98_clock),
    .reset(line_98_reset),
    .valid(line_98_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_97_clock = clock;
  assign line_97_reset = reset;
  assign line_97_valid = do_enq ^ line_97_valid_reg;
  assign line_98_clock = clock;
  assign line_98_reset = reset;
  assign line_98_valid = _T ^ line_98_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_97_valid_reg <= do_enq;
    line_98_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_97_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_98_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_10(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_99_clock;
  wire  line_99_reset;
  wire  line_99_valid;
  reg  line_99_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_100_clock;
  wire  line_100_reset;
  wire  line_100_valid;
  reg  line_100_valid_reg;
  GEN_w1_line #(.COVER_INDEX(99)) line_99 (
    .clock(line_99_clock),
    .reset(line_99_reset),
    .valid(line_99_valid)
  );
  GEN_w1_line #(.COVER_INDEX(100)) line_100 (
    .clock(line_100_clock),
    .reset(line_100_reset),
    .valid(line_100_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_99_clock = clock;
  assign line_99_reset = reset;
  assign line_99_valid = do_enq ^ line_99_valid_reg;
  assign line_100_clock = clock;
  assign line_100_reset = reset;
  assign line_100_valid = _T ^ line_100_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_99_valid_reg <= do_enq;
    line_100_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_99_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_100_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_11(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_101_clock;
  wire  line_101_reset;
  wire  line_101_valid;
  reg  line_101_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_102_clock;
  wire  line_102_reset;
  wire  line_102_valid;
  reg  line_102_valid_reg;
  GEN_w1_line #(.COVER_INDEX(101)) line_101 (
    .clock(line_101_clock),
    .reset(line_101_reset),
    .valid(line_101_valid)
  );
  GEN_w1_line #(.COVER_INDEX(102)) line_102 (
    .clock(line_102_clock),
    .reset(line_102_reset),
    .valid(line_102_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_101_clock = clock;
  assign line_101_reset = reset;
  assign line_101_valid = do_enq ^ line_101_valid_reg;
  assign line_102_clock = clock;
  assign line_102_reset = reset;
  assign line_102_valid = _T ^ line_102_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_101_valid_reg <= do_enq;
    line_102_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_101_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_102_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_12(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_103_clock;
  wire  line_103_reset;
  wire  line_103_valid;
  reg  line_103_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_104_clock;
  wire  line_104_reset;
  wire  line_104_valid;
  reg  line_104_valid_reg;
  GEN_w1_line #(.COVER_INDEX(103)) line_103 (
    .clock(line_103_clock),
    .reset(line_103_reset),
    .valid(line_103_valid)
  );
  GEN_w1_line #(.COVER_INDEX(104)) line_104 (
    .clock(line_104_clock),
    .reset(line_104_reset),
    .valid(line_104_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_103_clock = clock;
  assign line_103_reset = reset;
  assign line_103_valid = do_enq ^ line_103_valid_reg;
  assign line_104_clock = clock;
  assign line_104_reset = reset;
  assign line_104_valid = _T ^ line_104_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_103_valid_reg <= do_enq;
    line_104_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_103_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_104_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_13(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_105_clock;
  wire  line_105_reset;
  wire  line_105_valid;
  reg  line_105_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_106_clock;
  wire  line_106_reset;
  wire  line_106_valid;
  reg  line_106_valid_reg;
  GEN_w1_line #(.COVER_INDEX(105)) line_105 (
    .clock(line_105_clock),
    .reset(line_105_reset),
    .valid(line_105_valid)
  );
  GEN_w1_line #(.COVER_INDEX(106)) line_106 (
    .clock(line_106_clock),
    .reset(line_106_reset),
    .valid(line_106_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_105_clock = clock;
  assign line_105_reset = reset;
  assign line_105_valid = do_enq ^ line_105_valid_reg;
  assign line_106_clock = clock;
  assign line_106_reset = reset;
  assign line_106_valid = _T ^ line_106_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_105_valid_reg <= do_enq;
    line_106_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_105_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_106_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_14(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_107_clock;
  wire  line_107_reset;
  wire  line_107_valid;
  reg  line_107_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_108_clock;
  wire  line_108_reset;
  wire  line_108_valid;
  reg  line_108_valid_reg;
  GEN_w1_line #(.COVER_INDEX(107)) line_107 (
    .clock(line_107_clock),
    .reset(line_107_reset),
    .valid(line_107_valid)
  );
  GEN_w1_line #(.COVER_INDEX(108)) line_108 (
    .clock(line_108_clock),
    .reset(line_108_reset),
    .valid(line_108_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_107_clock = clock;
  assign line_107_reset = reset;
  assign line_107_valid = do_enq ^ line_107_valid_reg;
  assign line_108_clock = clock;
  assign line_108_reset = reset;
  assign line_108_valid = _T ^ line_108_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_107_valid_reg <= do_enq;
    line_108_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_107_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_108_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_15(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_109_clock;
  wire  line_109_reset;
  wire  line_109_valid;
  reg  line_109_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_110_clock;
  wire  line_110_reset;
  wire  line_110_valid;
  reg  line_110_valid_reg;
  GEN_w1_line #(.COVER_INDEX(109)) line_109 (
    .clock(line_109_clock),
    .reset(line_109_reset),
    .valid(line_109_valid)
  );
  GEN_w1_line #(.COVER_INDEX(110)) line_110 (
    .clock(line_110_clock),
    .reset(line_110_reset),
    .valid(line_110_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_109_clock = clock;
  assign line_109_reset = reset;
  assign line_109_valid = do_enq ^ line_109_valid_reg;
  assign line_110_clock = clock;
  assign line_110_reset = reset;
  assign line_110_valid = _T ^ line_110_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_109_valid_reg <= do_enq;
    line_110_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_109_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_110_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_16(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_111_clock;
  wire  line_111_reset;
  wire  line_111_valid;
  reg  line_111_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_112_clock;
  wire  line_112_reset;
  wire  line_112_valid;
  reg  line_112_valid_reg;
  GEN_w1_line #(.COVER_INDEX(111)) line_111 (
    .clock(line_111_clock),
    .reset(line_111_reset),
    .valid(line_111_valid)
  );
  GEN_w1_line #(.COVER_INDEX(112)) line_112 (
    .clock(line_112_clock),
    .reset(line_112_reset),
    .valid(line_112_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_111_clock = clock;
  assign line_111_reset = reset;
  assign line_111_valid = do_enq ^ line_111_valid_reg;
  assign line_112_clock = clock;
  assign line_112_reset = reset;
  assign line_112_valid = _T ^ line_112_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_111_valid_reg <= do_enq;
    line_112_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_111_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_112_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_17(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_113_clock;
  wire  line_113_reset;
  wire  line_113_valid;
  reg  line_113_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_114_clock;
  wire  line_114_reset;
  wire  line_114_valid;
  reg  line_114_valid_reg;
  GEN_w1_line #(.COVER_INDEX(113)) line_113 (
    .clock(line_113_clock),
    .reset(line_113_reset),
    .valid(line_113_valid)
  );
  GEN_w1_line #(.COVER_INDEX(114)) line_114 (
    .clock(line_114_clock),
    .reset(line_114_reset),
    .valid(line_114_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_113_clock = clock;
  assign line_113_reset = reset;
  assign line_113_valid = do_enq ^ line_113_valid_reg;
  assign line_114_clock = clock;
  assign line_114_reset = reset;
  assign line_114_valid = _T ^ line_114_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_113_valid_reg <= do_enq;
    line_114_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_113_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_114_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_18(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_115_clock;
  wire  line_115_reset;
  wire  line_115_valid;
  reg  line_115_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_116_clock;
  wire  line_116_reset;
  wire  line_116_valid;
  reg  line_116_valid_reg;
  GEN_w1_line #(.COVER_INDEX(115)) line_115 (
    .clock(line_115_clock),
    .reset(line_115_reset),
    .valid(line_115_valid)
  );
  GEN_w1_line #(.COVER_INDEX(116)) line_116 (
    .clock(line_116_clock),
    .reset(line_116_reset),
    .valid(line_116_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_115_clock = clock;
  assign line_115_reset = reset;
  assign line_115_valid = do_enq ^ line_115_valid_reg;
  assign line_116_clock = clock;
  assign line_116_reset = reset;
  assign line_116_valid = _T ^ line_116_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_115_valid_reg <= do_enq;
    line_116_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_115_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_116_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_19(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_117_clock;
  wire  line_117_reset;
  wire  line_117_valid;
  reg  line_117_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_118_clock;
  wire  line_118_reset;
  wire  line_118_valid;
  reg  line_118_valid_reg;
  GEN_w1_line #(.COVER_INDEX(117)) line_117 (
    .clock(line_117_clock),
    .reset(line_117_reset),
    .valid(line_117_valid)
  );
  GEN_w1_line #(.COVER_INDEX(118)) line_118 (
    .clock(line_118_clock),
    .reset(line_118_reset),
    .valid(line_118_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_117_clock = clock;
  assign line_117_reset = reset;
  assign line_117_valid = do_enq ^ line_117_valid_reg;
  assign line_118_clock = clock;
  assign line_118_reset = reset;
  assign line_118_valid = _T ^ line_118_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_117_valid_reg <= do_enq;
    line_118_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_117_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_118_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_20(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_119_clock;
  wire  line_119_reset;
  wire  line_119_valid;
  reg  line_119_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_120_clock;
  wire  line_120_reset;
  wire  line_120_valid;
  reg  line_120_valid_reg;
  GEN_w1_line #(.COVER_INDEX(119)) line_119 (
    .clock(line_119_clock),
    .reset(line_119_reset),
    .valid(line_119_valid)
  );
  GEN_w1_line #(.COVER_INDEX(120)) line_120 (
    .clock(line_120_clock),
    .reset(line_120_reset),
    .valid(line_120_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_119_clock = clock;
  assign line_119_reset = reset;
  assign line_119_valid = do_enq ^ line_119_valid_reg;
  assign line_120_clock = clock;
  assign line_120_reset = reset;
  assign line_120_valid = _T ^ line_120_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_119_valid_reg <= do_enq;
    line_120_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_119_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_120_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_21(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_121_clock;
  wire  line_121_reset;
  wire  line_121_valid;
  reg  line_121_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_122_clock;
  wire  line_122_reset;
  wire  line_122_valid;
  reg  line_122_valid_reg;
  GEN_w1_line #(.COVER_INDEX(121)) line_121 (
    .clock(line_121_clock),
    .reset(line_121_reset),
    .valid(line_121_valid)
  );
  GEN_w1_line #(.COVER_INDEX(122)) line_122 (
    .clock(line_122_clock),
    .reset(line_122_reset),
    .valid(line_122_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_121_clock = clock;
  assign line_121_reset = reset;
  assign line_121_valid = do_enq ^ line_121_valid_reg;
  assign line_122_clock = clock;
  assign line_122_reset = reset;
  assign line_122_valid = _T ^ line_122_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_121_valid_reg <= do_enq;
    line_122_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_121_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_122_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_22(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_123_clock;
  wire  line_123_reset;
  wire  line_123_valid;
  reg  line_123_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_124_clock;
  wire  line_124_reset;
  wire  line_124_valid;
  reg  line_124_valid_reg;
  GEN_w1_line #(.COVER_INDEX(123)) line_123 (
    .clock(line_123_clock),
    .reset(line_123_reset),
    .valid(line_123_valid)
  );
  GEN_w1_line #(.COVER_INDEX(124)) line_124 (
    .clock(line_124_clock),
    .reset(line_124_reset),
    .valid(line_124_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_123_clock = clock;
  assign line_123_reset = reset;
  assign line_123_valid = do_enq ^ line_123_valid_reg;
  assign line_124_clock = clock;
  assign line_124_reset = reset;
  assign line_124_valid = _T ^ line_124_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_123_valid_reg <= do_enq;
    line_124_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_123_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_124_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_23(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_125_clock;
  wire  line_125_reset;
  wire  line_125_valid;
  reg  line_125_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_126_clock;
  wire  line_126_reset;
  wire  line_126_valid;
  reg  line_126_valid_reg;
  GEN_w1_line #(.COVER_INDEX(125)) line_125 (
    .clock(line_125_clock),
    .reset(line_125_reset),
    .valid(line_125_valid)
  );
  GEN_w1_line #(.COVER_INDEX(126)) line_126 (
    .clock(line_126_clock),
    .reset(line_126_reset),
    .valid(line_126_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_125_clock = clock;
  assign line_125_reset = reset;
  assign line_125_valid = do_enq ^ line_125_valid_reg;
  assign line_126_clock = clock;
  assign line_126_reset = reset;
  assign line_126_valid = _T ^ line_126_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_125_valid_reg <= do_enq;
    line_126_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_125_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_126_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_24(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_127_clock;
  wire  line_127_reset;
  wire  line_127_valid;
  reg  line_127_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_128_clock;
  wire  line_128_reset;
  wire  line_128_valid;
  reg  line_128_valid_reg;
  GEN_w1_line #(.COVER_INDEX(127)) line_127 (
    .clock(line_127_clock),
    .reset(line_127_reset),
    .valid(line_127_valid)
  );
  GEN_w1_line #(.COVER_INDEX(128)) line_128 (
    .clock(line_128_clock),
    .reset(line_128_reset),
    .valid(line_128_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_127_clock = clock;
  assign line_127_reset = reset;
  assign line_127_valid = do_enq ^ line_127_valid_reg;
  assign line_128_clock = clock;
  assign line_128_reset = reset;
  assign line_128_valid = _T ^ line_128_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_127_valid_reg <= do_enq;
    line_128_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_127_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_128_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_25(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_129_clock;
  wire  line_129_reset;
  wire  line_129_valid;
  reg  line_129_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_130_clock;
  wire  line_130_reset;
  wire  line_130_valid;
  reg  line_130_valid_reg;
  GEN_w1_line #(.COVER_INDEX(129)) line_129 (
    .clock(line_129_clock),
    .reset(line_129_reset),
    .valid(line_129_valid)
  );
  GEN_w1_line #(.COVER_INDEX(130)) line_130 (
    .clock(line_130_clock),
    .reset(line_130_reset),
    .valid(line_130_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_129_clock = clock;
  assign line_129_reset = reset;
  assign line_129_valid = do_enq ^ line_129_valid_reg;
  assign line_130_clock = clock;
  assign line_130_reset = reset;
  assign line_130_valid = _T ^ line_130_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_129_valid_reg <= do_enq;
    line_130_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_129_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_130_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_26(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_131_clock;
  wire  line_131_reset;
  wire  line_131_valid;
  reg  line_131_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_132_clock;
  wire  line_132_reset;
  wire  line_132_valid;
  reg  line_132_valid_reg;
  GEN_w1_line #(.COVER_INDEX(131)) line_131 (
    .clock(line_131_clock),
    .reset(line_131_reset),
    .valid(line_131_valid)
  );
  GEN_w1_line #(.COVER_INDEX(132)) line_132 (
    .clock(line_132_clock),
    .reset(line_132_reset),
    .valid(line_132_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_131_clock = clock;
  assign line_131_reset = reset;
  assign line_131_valid = do_enq ^ line_131_valid_reg;
  assign line_132_clock = clock;
  assign line_132_reset = reset;
  assign line_132_valid = _T ^ line_132_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_131_valid_reg <= do_enq;
    line_132_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_131_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_132_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_27(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_133_clock;
  wire  line_133_reset;
  wire  line_133_valid;
  reg  line_133_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_134_clock;
  wire  line_134_reset;
  wire  line_134_valid;
  reg  line_134_valid_reg;
  GEN_w1_line #(.COVER_INDEX(133)) line_133 (
    .clock(line_133_clock),
    .reset(line_133_reset),
    .valid(line_133_valid)
  );
  GEN_w1_line #(.COVER_INDEX(134)) line_134 (
    .clock(line_134_clock),
    .reset(line_134_reset),
    .valid(line_134_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_133_clock = clock;
  assign line_133_reset = reset;
  assign line_133_valid = do_enq ^ line_133_valid_reg;
  assign line_134_clock = clock;
  assign line_134_reset = reset;
  assign line_134_valid = _T ^ line_134_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_133_valid_reg <= do_enq;
    line_134_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_133_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_134_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_28(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_135_clock;
  wire  line_135_reset;
  wire  line_135_valid;
  reg  line_135_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_136_clock;
  wire  line_136_reset;
  wire  line_136_valid;
  reg  line_136_valid_reg;
  GEN_w1_line #(.COVER_INDEX(135)) line_135 (
    .clock(line_135_clock),
    .reset(line_135_reset),
    .valid(line_135_valid)
  );
  GEN_w1_line #(.COVER_INDEX(136)) line_136 (
    .clock(line_136_clock),
    .reset(line_136_reset),
    .valid(line_136_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_135_clock = clock;
  assign line_135_reset = reset;
  assign line_135_valid = do_enq ^ line_135_valid_reg;
  assign line_136_clock = clock;
  assign line_136_reset = reset;
  assign line_136_valid = _T ^ line_136_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_135_valid_reg <= do_enq;
    line_136_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_135_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_136_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_29(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_137_clock;
  wire  line_137_reset;
  wire  line_137_valid;
  reg  line_137_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_138_clock;
  wire  line_138_reset;
  wire  line_138_valid;
  reg  line_138_valid_reg;
  GEN_w1_line #(.COVER_INDEX(137)) line_137 (
    .clock(line_137_clock),
    .reset(line_137_reset),
    .valid(line_137_valid)
  );
  GEN_w1_line #(.COVER_INDEX(138)) line_138 (
    .clock(line_138_clock),
    .reset(line_138_reset),
    .valid(line_138_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_137_clock = clock;
  assign line_137_reset = reset;
  assign line_137_valid = do_enq ^ line_137_valid_reg;
  assign line_138_clock = clock;
  assign line_138_reset = reset;
  assign line_138_valid = _T ^ line_138_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_137_valid_reg <= do_enq;
    line_138_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_137_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_138_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_30(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_139_clock;
  wire  line_139_reset;
  wire  line_139_valid;
  reg  line_139_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_140_clock;
  wire  line_140_reset;
  wire  line_140_valid;
  reg  line_140_valid_reg;
  GEN_w1_line #(.COVER_INDEX(139)) line_139 (
    .clock(line_139_clock),
    .reset(line_139_reset),
    .valid(line_139_valid)
  );
  GEN_w1_line #(.COVER_INDEX(140)) line_140 (
    .clock(line_140_clock),
    .reset(line_140_reset),
    .valid(line_140_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_139_clock = clock;
  assign line_139_reset = reset;
  assign line_139_valid = do_enq ^ line_139_valid_reg;
  assign line_140_clock = clock;
  assign line_140_reset = reset;
  assign line_140_valid = _T ^ line_140_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_139_valid_reg <= do_enq;
    line_140_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_139_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_140_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_31(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_141_clock;
  wire  line_141_reset;
  wire  line_141_valid;
  reg  line_141_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_142_clock;
  wire  line_142_reset;
  wire  line_142_valid;
  reg  line_142_valid_reg;
  GEN_w1_line #(.COVER_INDEX(141)) line_141 (
    .clock(line_141_clock),
    .reset(line_141_reset),
    .valid(line_141_valid)
  );
  GEN_w1_line #(.COVER_INDEX(142)) line_142 (
    .clock(line_142_clock),
    .reset(line_142_reset),
    .valid(line_142_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_141_clock = clock;
  assign line_141_reset = reset;
  assign line_141_valid = do_enq ^ line_141_valid_reg;
  assign line_142_clock = clock;
  assign line_142_reset = reset;
  assign line_142_valid = _T ^ line_142_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_141_valid_reg <= do_enq;
    line_142_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_141_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_142_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_32(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_143_clock;
  wire  line_143_reset;
  wire  line_143_valid;
  reg  line_143_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_144_clock;
  wire  line_144_reset;
  wire  line_144_valid;
  reg  line_144_valid_reg;
  GEN_w1_line #(.COVER_INDEX(143)) line_143 (
    .clock(line_143_clock),
    .reset(line_143_reset),
    .valid(line_143_valid)
  );
  GEN_w1_line #(.COVER_INDEX(144)) line_144 (
    .clock(line_144_clock),
    .reset(line_144_reset),
    .valid(line_144_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_143_clock = clock;
  assign line_143_reset = reset;
  assign line_143_valid = do_enq ^ line_143_valid_reg;
  assign line_144_clock = clock;
  assign line_144_reset = reset;
  assign line_144_valid = _T ^ line_144_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_143_valid_reg <= do_enq;
    line_144_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_143_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_144_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_33(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_tl_state_source // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_145_clock;
  wire  line_145_reset;
  wire  line_145_valid;
  reg  line_145_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_146_clock;
  wire  line_146_reset;
  wire  line_146_valid;
  reg  line_146_valid_reg;
  GEN_w1_line #(.COVER_INDEX(145)) line_145 (
    .clock(line_145_clock),
    .reset(line_145_reset),
    .valid(line_145_valid)
  );
  GEN_w1_line #(.COVER_INDEX(146)) line_146 (
    .clock(line_146_clock),
    .reset(line_146_reset),
    .valid(line_146_valid)
  );
  assign ram_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_size_io_deq_bits_MPORT_data = ram_tl_state_size[ram_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_size_MPORT_data = io_enq_bits_tl_state_size;
  assign ram_tl_state_size_MPORT_addr = 1'h0;
  assign ram_tl_state_size_MPORT_mask = 1'h1;
  assign ram_tl_state_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tl_state_source_io_deq_bits_MPORT_data = ram_tl_state_source[ram_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_tl_state_source_MPORT_data = io_enq_bits_tl_state_source;
  assign ram_tl_state_source_MPORT_addr = 1'h0;
  assign ram_tl_state_source_MPORT_mask = 1'h1;
  assign ram_tl_state_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_145_clock = clock;
  assign line_145_reset = reset;
  assign line_145_valid = do_enq ^ line_145_valid_reg;
  assign line_146_clock = clock;
  assign line_146_reset = reset;
  assign line_146_valid = _T ^ line_146_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_tl_state_size = ram_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_tl_state_source = ram_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_tl_state_size_MPORT_en & ram_tl_state_size_MPORT_mask) begin
      ram_tl_state_size[ram_tl_state_size_MPORT_addr] <= ram_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_tl_state_source_MPORT_en & ram_tl_state_source_MPORT_mask) begin
      ram_tl_state_source[ram_tl_state_source_MPORT_addr] <= ram_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_145_valid_reg <= do_enq;
    line_146_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_size[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tl_state_source[initvar] = _RAND_1[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_145_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_146_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4UserYanker(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
`endif // RANDOMIZE_REG_INIT
  wire  Queue_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_1_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_1_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_1_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_1_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_1_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_2_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_2_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_2_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_2_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_2_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_3_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_3_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_3_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_3_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_3_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_4_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_4_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_4_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_4_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_4_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_5_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_5_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_5_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_5_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_5_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_6_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_6_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_6_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_6_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_6_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_7_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_7_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_7_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_7_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_7_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_8_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_8_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_8_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_8_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_8_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_9_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_9_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_9_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_9_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_9_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_10_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_10_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_10_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_10_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_10_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_11_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_11_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_11_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_11_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_11_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_12_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_12_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_12_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_12_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_12_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_13_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_13_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_13_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_13_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_13_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_14_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_14_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_14_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_14_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_14_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_15_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_15_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_15_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_15_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_15_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_16_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_16_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_16_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_16_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_16_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_17_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_17_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_17_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_17_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_17_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_18_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_18_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_18_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_18_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_18_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_19_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_19_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_19_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_19_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_19_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_20_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_20_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_20_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_20_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_20_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_21_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_21_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_21_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_21_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_21_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_22_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_22_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_22_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_22_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_22_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_23_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_23_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_23_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_23_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_23_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_24_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_24_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_24_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_24_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_24_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_25_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_25_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_25_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_25_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_25_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_26_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_26_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_26_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_26_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_26_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_27_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_27_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_27_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_27_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_27_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_28_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_28_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_28_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_28_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_28_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_29_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_29_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_29_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_29_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_29_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_30_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_30_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_30_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_30_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_30_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_io_enq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_31_io_enq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_31_io_enq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_io_deq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  Queue_31_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_31_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire [3:0] Queue_31_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
  wire  line_147_clock;
  wire  line_147_reset;
  wire  line_147_valid;
  reg  line_147_valid_reg;
  wire  _ar_ready_WIRE_0 = Queue_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  line_148_clock;
  wire  line_148_reset;
  wire  line_148_valid;
  reg  line_148_valid_reg;
  wire  _ar_ready_WIRE_1 = Queue_1_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_165 = 4'h1 == auto_in_ar_bits_id ? _ar_ready_WIRE_1 : _ar_ready_WIRE_0; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_149_clock;
  wire  line_149_reset;
  wire  line_149_valid;
  reg  line_149_valid_reg;
  wire  _ar_ready_WIRE_2 = Queue_2_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_166 = 4'h2 == auto_in_ar_bits_id ? _ar_ready_WIRE_2 : _GEN_165; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_150_clock;
  wire  line_150_reset;
  wire  line_150_valid;
  reg  line_150_valid_reg;
  wire  _ar_ready_WIRE_3 = Queue_3_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_167 = 4'h3 == auto_in_ar_bits_id ? _ar_ready_WIRE_3 : _GEN_166; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_151_clock;
  wire  line_151_reset;
  wire  line_151_valid;
  reg  line_151_valid_reg;
  wire  _ar_ready_WIRE_4 = Queue_4_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_168 = 4'h4 == auto_in_ar_bits_id ? _ar_ready_WIRE_4 : _GEN_167; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_152_clock;
  wire  line_152_reset;
  wire  line_152_valid;
  reg  line_152_valid_reg;
  wire  _ar_ready_WIRE_5 = Queue_5_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_169 = 4'h5 == auto_in_ar_bits_id ? _ar_ready_WIRE_5 : _GEN_168; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_153_clock;
  wire  line_153_reset;
  wire  line_153_valid;
  reg  line_153_valid_reg;
  wire  _ar_ready_WIRE_6 = Queue_6_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_170 = 4'h6 == auto_in_ar_bits_id ? _ar_ready_WIRE_6 : _GEN_169; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_154_clock;
  wire  line_154_reset;
  wire  line_154_valid;
  reg  line_154_valid_reg;
  wire  _ar_ready_WIRE_7 = Queue_7_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_171 = 4'h7 == auto_in_ar_bits_id ? _ar_ready_WIRE_7 : _GEN_170; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_155_clock;
  wire  line_155_reset;
  wire  line_155_valid;
  reg  line_155_valid_reg;
  wire  _ar_ready_WIRE_8 = Queue_8_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_172 = 4'h8 == auto_in_ar_bits_id ? _ar_ready_WIRE_8 : _GEN_171; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_156_clock;
  wire  line_156_reset;
  wire  line_156_valid;
  reg  line_156_valid_reg;
  wire  _ar_ready_WIRE_9 = Queue_9_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_173 = 4'h9 == auto_in_ar_bits_id ? _ar_ready_WIRE_9 : _GEN_172; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_157_clock;
  wire  line_157_reset;
  wire  line_157_valid;
  reg  line_157_valid_reg;
  wire  _ar_ready_WIRE_10 = Queue_10_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_174 = 4'ha == auto_in_ar_bits_id ? _ar_ready_WIRE_10 : _GEN_173; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_158_clock;
  wire  line_158_reset;
  wire  line_158_valid;
  reg  line_158_valid_reg;
  wire  _ar_ready_WIRE_11 = Queue_11_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_175 = 4'hb == auto_in_ar_bits_id ? _ar_ready_WIRE_11 : _GEN_174; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_159_clock;
  wire  line_159_reset;
  wire  line_159_valid;
  reg  line_159_valid_reg;
  wire  _ar_ready_WIRE_12 = Queue_12_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_176 = 4'hc == auto_in_ar_bits_id ? _ar_ready_WIRE_12 : _GEN_175; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_160_clock;
  wire  line_160_reset;
  wire  line_160_valid;
  reg  line_160_valid_reg;
  wire  _ar_ready_WIRE_13 = Queue_13_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_177 = 4'hd == auto_in_ar_bits_id ? _ar_ready_WIRE_13 : _GEN_176; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_161_clock;
  wire  line_161_reset;
  wire  line_161_valid;
  reg  line_161_valid_reg;
  wire  _ar_ready_WIRE_14 = Queue_14_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_178 = 4'he == auto_in_ar_bits_id ? _ar_ready_WIRE_14 : _GEN_177; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_162_clock;
  wire  line_162_reset;
  wire  line_162_valid;
  reg  line_162_valid_reg;
  wire  _ar_ready_WIRE_15 = Queue_15_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 56:{29,29}]
  wire  _GEN_179 = 4'hf == auto_in_ar_bits_id ? _ar_ready_WIRE_15 : _GEN_178; // @[src/main/scala/amba/axi4/UserYanker.scala 57:{36,36}]
  wire  line_163_clock;
  wire  line_163_reset;
  wire  line_163_valid;
  reg  line_163_valid_reg;
  wire  line_164_clock;
  wire  line_164_reset;
  wire  line_164_valid;
  reg  line_164_valid_reg;
  wire  line_165_clock;
  wire  line_165_reset;
  wire  line_165_valid;
  reg  line_165_valid_reg;
  wire  line_166_clock;
  wire  line_166_reset;
  wire  line_166_valid;
  reg  line_166_valid_reg;
  wire  line_167_clock;
  wire  line_167_reset;
  wire  line_167_valid;
  reg  line_167_valid_reg;
  wire  line_168_clock;
  wire  line_168_reset;
  wire  line_168_valid;
  reg  line_168_valid_reg;
  wire  line_169_clock;
  wire  line_169_reset;
  wire  line_169_valid;
  reg  line_169_valid_reg;
  wire  line_170_clock;
  wire  line_170_reset;
  wire  line_170_valid;
  reg  line_170_valid_reg;
  wire  line_171_clock;
  wire  line_171_reset;
  wire  line_171_valid;
  reg  line_171_valid_reg;
  wire  line_172_clock;
  wire  line_172_reset;
  wire  line_172_valid;
  reg  line_172_valid_reg;
  wire  line_173_clock;
  wire  line_173_reset;
  wire  line_173_valid;
  reg  line_173_valid_reg;
  wire  line_174_clock;
  wire  line_174_reset;
  wire  line_174_valid;
  reg  line_174_valid_reg;
  wire  line_175_clock;
  wire  line_175_reset;
  wire  line_175_valid;
  reg  line_175_valid_reg;
  wire  line_176_clock;
  wire  line_176_reset;
  wire  line_176_valid;
  reg  line_176_valid_reg;
  wire  line_177_clock;
  wire  line_177_reset;
  wire  line_177_valid;
  reg  line_177_valid_reg;
  wire  line_178_clock;
  wire  line_178_reset;
  wire  line_178_valid;
  reg  line_178_valid_reg;
  wire  line_179_clock;
  wire  line_179_reset;
  wire  line_179_valid;
  reg  line_179_valid_reg;
  wire  _r_valid_WIRE_0 = Queue_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  line_180_clock;
  wire  line_180_reset;
  wire  line_180_valid;
  reg  line_180_valid_reg;
  wire  _r_valid_WIRE_1 = Queue_1_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_181 = 4'h1 == auto_out_r_bits_id ? _r_valid_WIRE_1 : _r_valid_WIRE_0; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_181_clock;
  wire  line_181_reset;
  wire  line_181_valid;
  reg  line_181_valid_reg;
  wire  _r_valid_WIRE_2 = Queue_2_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_182 = 4'h2 == auto_out_r_bits_id ? _r_valid_WIRE_2 : _GEN_181; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_182_clock;
  wire  line_182_reset;
  wire  line_182_valid;
  reg  line_182_valid_reg;
  wire  _r_valid_WIRE_3 = Queue_3_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_183 = 4'h3 == auto_out_r_bits_id ? _r_valid_WIRE_3 : _GEN_182; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_183_clock;
  wire  line_183_reset;
  wire  line_183_valid;
  reg  line_183_valid_reg;
  wire  _r_valid_WIRE_4 = Queue_4_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_184 = 4'h4 == auto_out_r_bits_id ? _r_valid_WIRE_4 : _GEN_183; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_184_clock;
  wire  line_184_reset;
  wire  line_184_valid;
  reg  line_184_valid_reg;
  wire  _r_valid_WIRE_5 = Queue_5_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_185 = 4'h5 == auto_out_r_bits_id ? _r_valid_WIRE_5 : _GEN_184; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_185_clock;
  wire  line_185_reset;
  wire  line_185_valid;
  reg  line_185_valid_reg;
  wire  _r_valid_WIRE_6 = Queue_6_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_186 = 4'h6 == auto_out_r_bits_id ? _r_valid_WIRE_6 : _GEN_185; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_186_clock;
  wire  line_186_reset;
  wire  line_186_valid;
  reg  line_186_valid_reg;
  wire  _r_valid_WIRE_7 = Queue_7_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_187 = 4'h7 == auto_out_r_bits_id ? _r_valid_WIRE_7 : _GEN_186; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_187_clock;
  wire  line_187_reset;
  wire  line_187_valid;
  reg  line_187_valid_reg;
  wire  _r_valid_WIRE_8 = Queue_8_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_188 = 4'h8 == auto_out_r_bits_id ? _r_valid_WIRE_8 : _GEN_187; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_188_clock;
  wire  line_188_reset;
  wire  line_188_valid;
  reg  line_188_valid_reg;
  wire  _r_valid_WIRE_9 = Queue_9_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_189 = 4'h9 == auto_out_r_bits_id ? _r_valid_WIRE_9 : _GEN_188; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_189_clock;
  wire  line_189_reset;
  wire  line_189_valid;
  reg  line_189_valid_reg;
  wire  _r_valid_WIRE_10 = Queue_10_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_190 = 4'ha == auto_out_r_bits_id ? _r_valid_WIRE_10 : _GEN_189; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_190_clock;
  wire  line_190_reset;
  wire  line_190_valid;
  reg  line_190_valid_reg;
  wire  _r_valid_WIRE_11 = Queue_11_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_191 = 4'hb == auto_out_r_bits_id ? _r_valid_WIRE_11 : _GEN_190; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_191_clock;
  wire  line_191_reset;
  wire  line_191_valid;
  reg  line_191_valid_reg;
  wire  _r_valid_WIRE_12 = Queue_12_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_192 = 4'hc == auto_out_r_bits_id ? _r_valid_WIRE_12 : _GEN_191; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_192_clock;
  wire  line_192_reset;
  wire  line_192_valid;
  reg  line_192_valid_reg;
  wire  _r_valid_WIRE_13 = Queue_13_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_193 = 4'hd == auto_out_r_bits_id ? _r_valid_WIRE_13 : _GEN_192; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_193_clock;
  wire  line_193_reset;
  wire  line_193_valid;
  reg  line_193_valid_reg;
  wire  _r_valid_WIRE_14 = Queue_14_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_194 = 4'he == auto_out_r_bits_id ? _r_valid_WIRE_14 : _GEN_193; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  line_194_clock;
  wire  line_194_reset;
  wire  line_194_valid;
  reg  line_194_valid_reg;
  wire  _r_valid_WIRE_15 = Queue_15_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 64:{28,28}]
  wire  _GEN_195 = 4'hf == auto_out_r_bits_id ? _r_valid_WIRE_15 : _GEN_194; // @[src/main/scala/amba/axi4/UserYanker.scala 66:{28,28}]
  wire  _T_3 = ~reset; // @[src/main/scala/amba/axi4/UserYanker.scala 66:14]
  wire  line_195_clock;
  wire  line_195_reset;
  wire  line_195_valid;
  reg  line_195_valid_reg;
  wire  _T_4 = ~(~auto_out_r_valid | _GEN_195); // @[src/main/scala/amba/axi4/UserYanker.scala 66:14]
  wire  line_196_clock;
  wire  line_196_reset;
  wire  line_196_valid;
  reg  line_196_valid_reg;
  wire  line_197_clock;
  wire  line_197_reset;
  wire  line_197_valid;
  reg  line_197_valid_reg;
  wire [3:0] _r_bits_WIRE_0_tl_state_source = Queue_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire  line_198_clock;
  wire  line_198_reset;
  wire  line_198_valid;
  reg  line_198_valid_reg;
  wire [3:0] _r_bits_WIRE_1_tl_state_source = Queue_1_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_197 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_tl_state_source : _r_bits_WIRE_0_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_199_clock;
  wire  line_199_reset;
  wire  line_199_valid;
  reg  line_199_valid_reg;
  wire [3:0] _r_bits_WIRE_2_tl_state_source = Queue_2_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_198 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_tl_state_source : _GEN_197; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_200_clock;
  wire  line_200_reset;
  wire  line_200_valid;
  reg  line_200_valid_reg;
  wire [3:0] _r_bits_WIRE_3_tl_state_source = Queue_3_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_199 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_tl_state_source : _GEN_198; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_201_clock;
  wire  line_201_reset;
  wire  line_201_valid;
  reg  line_201_valid_reg;
  wire [3:0] _r_bits_WIRE_4_tl_state_source = Queue_4_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_200 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_tl_state_source : _GEN_199; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_202_clock;
  wire  line_202_reset;
  wire  line_202_valid;
  reg  line_202_valid_reg;
  wire [3:0] _r_bits_WIRE_5_tl_state_source = Queue_5_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_201 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_tl_state_source : _GEN_200; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_203_clock;
  wire  line_203_reset;
  wire  line_203_valid;
  reg  line_203_valid_reg;
  wire [3:0] _r_bits_WIRE_6_tl_state_source = Queue_6_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_202 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_tl_state_source : _GEN_201; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_204_clock;
  wire  line_204_reset;
  wire  line_204_valid;
  reg  line_204_valid_reg;
  wire [3:0] _r_bits_WIRE_7_tl_state_source = Queue_7_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_203 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_tl_state_source : _GEN_202; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_205_clock;
  wire  line_205_reset;
  wire  line_205_valid;
  reg  line_205_valid_reg;
  wire [3:0] _r_bits_WIRE_8_tl_state_source = Queue_8_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_204 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_tl_state_source : _GEN_203; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_206_clock;
  wire  line_206_reset;
  wire  line_206_valid;
  reg  line_206_valid_reg;
  wire [3:0] _r_bits_WIRE_9_tl_state_source = Queue_9_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_205 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_tl_state_source : _GEN_204; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_207_clock;
  wire  line_207_reset;
  wire  line_207_valid;
  reg  line_207_valid_reg;
  wire [3:0] _r_bits_WIRE_10_tl_state_source = Queue_10_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_206 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_tl_state_source : _GEN_205; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_208_clock;
  wire  line_208_reset;
  wire  line_208_valid;
  reg  line_208_valid_reg;
  wire [3:0] _r_bits_WIRE_11_tl_state_source = Queue_11_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_207 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_tl_state_source : _GEN_206; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_209_clock;
  wire  line_209_reset;
  wire  line_209_valid;
  reg  line_209_valid_reg;
  wire [3:0] _r_bits_WIRE_12_tl_state_source = Queue_12_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_208 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_tl_state_source : _GEN_207; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_210_clock;
  wire  line_210_reset;
  wire  line_210_valid;
  reg  line_210_valid_reg;
  wire [3:0] _r_bits_WIRE_13_tl_state_source = Queue_13_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_209 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_tl_state_source : _GEN_208; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_211_clock;
  wire  line_211_reset;
  wire  line_211_valid;
  reg  line_211_valid_reg;
  wire [3:0] _r_bits_WIRE_14_tl_state_source = Queue_14_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_210 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_tl_state_source : _GEN_209; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_212_clock;
  wire  line_212_reset;
  wire  line_212_valid;
  reg  line_212_valid_reg;
  wire [3:0] _r_bits_WIRE_15_tl_state_source = Queue_15_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire  line_213_clock;
  wire  line_213_reset;
  wire  line_213_valid;
  reg  line_213_valid_reg;
  wire [3:0] _r_bits_WIRE_0_tl_state_size = Queue_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire  line_214_clock;
  wire  line_214_reset;
  wire  line_214_valid;
  reg  line_214_valid_reg;
  wire [3:0] _r_bits_WIRE_1_tl_state_size = Queue_1_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_213 = 4'h1 == auto_out_r_bits_id ? _r_bits_WIRE_1_tl_state_size : _r_bits_WIRE_0_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_215_clock;
  wire  line_215_reset;
  wire  line_215_valid;
  reg  line_215_valid_reg;
  wire [3:0] _r_bits_WIRE_2_tl_state_size = Queue_2_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_214 = 4'h2 == auto_out_r_bits_id ? _r_bits_WIRE_2_tl_state_size : _GEN_213; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_216_clock;
  wire  line_216_reset;
  wire  line_216_valid;
  reg  line_216_valid_reg;
  wire [3:0] _r_bits_WIRE_3_tl_state_size = Queue_3_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_215 = 4'h3 == auto_out_r_bits_id ? _r_bits_WIRE_3_tl_state_size : _GEN_214; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_217_clock;
  wire  line_217_reset;
  wire  line_217_valid;
  reg  line_217_valid_reg;
  wire [3:0] _r_bits_WIRE_4_tl_state_size = Queue_4_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_216 = 4'h4 == auto_out_r_bits_id ? _r_bits_WIRE_4_tl_state_size : _GEN_215; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_218_clock;
  wire  line_218_reset;
  wire  line_218_valid;
  reg  line_218_valid_reg;
  wire [3:0] _r_bits_WIRE_5_tl_state_size = Queue_5_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_217 = 4'h5 == auto_out_r_bits_id ? _r_bits_WIRE_5_tl_state_size : _GEN_216; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_219_clock;
  wire  line_219_reset;
  wire  line_219_valid;
  reg  line_219_valid_reg;
  wire [3:0] _r_bits_WIRE_6_tl_state_size = Queue_6_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_218 = 4'h6 == auto_out_r_bits_id ? _r_bits_WIRE_6_tl_state_size : _GEN_217; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_220_clock;
  wire  line_220_reset;
  wire  line_220_valid;
  reg  line_220_valid_reg;
  wire [3:0] _r_bits_WIRE_7_tl_state_size = Queue_7_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_219 = 4'h7 == auto_out_r_bits_id ? _r_bits_WIRE_7_tl_state_size : _GEN_218; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_221_clock;
  wire  line_221_reset;
  wire  line_221_valid;
  reg  line_221_valid_reg;
  wire [3:0] _r_bits_WIRE_8_tl_state_size = Queue_8_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_220 = 4'h8 == auto_out_r_bits_id ? _r_bits_WIRE_8_tl_state_size : _GEN_219; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_222_clock;
  wire  line_222_reset;
  wire  line_222_valid;
  reg  line_222_valid_reg;
  wire [3:0] _r_bits_WIRE_9_tl_state_size = Queue_9_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_221 = 4'h9 == auto_out_r_bits_id ? _r_bits_WIRE_9_tl_state_size : _GEN_220; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_223_clock;
  wire  line_223_reset;
  wire  line_223_valid;
  reg  line_223_valid_reg;
  wire [3:0] _r_bits_WIRE_10_tl_state_size = Queue_10_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_222 = 4'ha == auto_out_r_bits_id ? _r_bits_WIRE_10_tl_state_size : _GEN_221; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_224_clock;
  wire  line_224_reset;
  wire  line_224_valid;
  reg  line_224_valid_reg;
  wire [3:0] _r_bits_WIRE_11_tl_state_size = Queue_11_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_223 = 4'hb == auto_out_r_bits_id ? _r_bits_WIRE_11_tl_state_size : _GEN_222; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_225_clock;
  wire  line_225_reset;
  wire  line_225_valid;
  reg  line_225_valid_reg;
  wire [3:0] _r_bits_WIRE_12_tl_state_size = Queue_12_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_224 = 4'hc == auto_out_r_bits_id ? _r_bits_WIRE_12_tl_state_size : _GEN_223; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_226_clock;
  wire  line_226_reset;
  wire  line_226_valid;
  reg  line_226_valid_reg;
  wire [3:0] _r_bits_WIRE_13_tl_state_size = Queue_13_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_225 = 4'hd == auto_out_r_bits_id ? _r_bits_WIRE_13_tl_state_size : _GEN_224; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_227_clock;
  wire  line_227_reset;
  wire  line_227_valid;
  reg  line_227_valid_reg;
  wire [3:0] _r_bits_WIRE_14_tl_state_size = Queue_14_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [3:0] _GEN_226 = 4'he == auto_out_r_bits_id ? _r_bits_WIRE_14_tl_state_size : _GEN_225; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  wire  line_228_clock;
  wire  line_228_reset;
  wire  line_228_valid;
  reg  line_228_valid_reg;
  wire [3:0] _r_bits_WIRE_15_tl_state_size = Queue_15_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 65:{27,27}]
  wire [15:0] _arsel_T = 16'h1 << auto_in_ar_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  arsel_0 = _arsel_T[0]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_1 = _arsel_T[1]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_2 = _arsel_T[2]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_3 = _arsel_T[3]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_4 = _arsel_T[4]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_5 = _arsel_T[5]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_6 = _arsel_T[6]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_7 = _arsel_T[7]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_8 = _arsel_T[8]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_9 = _arsel_T[9]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_10 = _arsel_T[10]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_11 = _arsel_T[11]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_12 = _arsel_T[12]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_13 = _arsel_T[13]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_14 = _arsel_T[14]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire  arsel_15 = _arsel_T[15]; // @[src/main/scala/amba/axi4/UserYanker.scala 72:55]
  wire [15:0] _rsel_T = 16'h1 << auto_out_r_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  rsel_0 = _rsel_T[0]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_1 = _rsel_T[1]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_2 = _rsel_T[2]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_3 = _rsel_T[3]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_4 = _rsel_T[4]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_5 = _rsel_T[5]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_6 = _rsel_T[6]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_7 = _rsel_T[7]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_8 = _rsel_T[8]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_9 = _rsel_T[9]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_10 = _rsel_T[10]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_11 = _rsel_T[11]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_12 = _rsel_T[12]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_13 = _rsel_T[13]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_14 = _rsel_T[14]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  rsel_15 = _rsel_T[15]; // @[src/main/scala/amba/axi4/UserYanker.scala 73:55]
  wire  line_229_clock;
  wire  line_229_reset;
  wire  line_229_valid;
  reg  line_229_valid_reg;
  wire  _aw_ready_WIRE_0 = Queue_16_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  line_230_clock;
  wire  line_230_reset;
  wire  line_230_valid;
  reg  line_230_valid_reg;
  wire  _aw_ready_WIRE_1 = Queue_17_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_229 = 4'h1 == auto_in_aw_bits_id ? _aw_ready_WIRE_1 : _aw_ready_WIRE_0; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_231_clock;
  wire  line_231_reset;
  wire  line_231_valid;
  reg  line_231_valid_reg;
  wire  _aw_ready_WIRE_2 = Queue_18_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_230 = 4'h2 == auto_in_aw_bits_id ? _aw_ready_WIRE_2 : _GEN_229; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_232_clock;
  wire  line_232_reset;
  wire  line_232_valid;
  reg  line_232_valid_reg;
  wire  _aw_ready_WIRE_3 = Queue_19_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_231 = 4'h3 == auto_in_aw_bits_id ? _aw_ready_WIRE_3 : _GEN_230; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_233_clock;
  wire  line_233_reset;
  wire  line_233_valid;
  reg  line_233_valid_reg;
  wire  _aw_ready_WIRE_4 = Queue_20_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_232 = 4'h4 == auto_in_aw_bits_id ? _aw_ready_WIRE_4 : _GEN_231; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_234_clock;
  wire  line_234_reset;
  wire  line_234_valid;
  reg  line_234_valid_reg;
  wire  _aw_ready_WIRE_5 = Queue_21_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_233 = 4'h5 == auto_in_aw_bits_id ? _aw_ready_WIRE_5 : _GEN_232; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_235_clock;
  wire  line_235_reset;
  wire  line_235_valid;
  reg  line_235_valid_reg;
  wire  _aw_ready_WIRE_6 = Queue_22_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_234 = 4'h6 == auto_in_aw_bits_id ? _aw_ready_WIRE_6 : _GEN_233; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_236_clock;
  wire  line_236_reset;
  wire  line_236_valid;
  reg  line_236_valid_reg;
  wire  _aw_ready_WIRE_7 = Queue_23_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_235 = 4'h7 == auto_in_aw_bits_id ? _aw_ready_WIRE_7 : _GEN_234; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_237_clock;
  wire  line_237_reset;
  wire  line_237_valid;
  reg  line_237_valid_reg;
  wire  _aw_ready_WIRE_8 = Queue_24_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_236 = 4'h8 == auto_in_aw_bits_id ? _aw_ready_WIRE_8 : _GEN_235; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_238_clock;
  wire  line_238_reset;
  wire  line_238_valid;
  reg  line_238_valid_reg;
  wire  _aw_ready_WIRE_9 = Queue_25_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_237 = 4'h9 == auto_in_aw_bits_id ? _aw_ready_WIRE_9 : _GEN_236; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_239_clock;
  wire  line_239_reset;
  wire  line_239_valid;
  reg  line_239_valid_reg;
  wire  _aw_ready_WIRE_10 = Queue_26_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_238 = 4'ha == auto_in_aw_bits_id ? _aw_ready_WIRE_10 : _GEN_237; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_240_clock;
  wire  line_240_reset;
  wire  line_240_valid;
  reg  line_240_valid_reg;
  wire  _aw_ready_WIRE_11 = Queue_27_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_239 = 4'hb == auto_in_aw_bits_id ? _aw_ready_WIRE_11 : _GEN_238; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_241_clock;
  wire  line_241_reset;
  wire  line_241_valid;
  reg  line_241_valid_reg;
  wire  _aw_ready_WIRE_12 = Queue_28_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_240 = 4'hc == auto_in_aw_bits_id ? _aw_ready_WIRE_12 : _GEN_239; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_242_clock;
  wire  line_242_reset;
  wire  line_242_valid;
  reg  line_242_valid_reg;
  wire  _aw_ready_WIRE_13 = Queue_29_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_241 = 4'hd == auto_in_aw_bits_id ? _aw_ready_WIRE_13 : _GEN_240; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_243_clock;
  wire  line_243_reset;
  wire  line_243_valid;
  reg  line_243_valid_reg;
  wire  _aw_ready_WIRE_14 = Queue_30_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_242 = 4'he == auto_in_aw_bits_id ? _aw_ready_WIRE_14 : _GEN_241; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_244_clock;
  wire  line_244_reset;
  wire  line_244_valid;
  reg  line_244_valid_reg;
  wire  _aw_ready_WIRE_15 = Queue_31_io_enq_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 85:{29,29}]
  wire  _GEN_243 = 4'hf == auto_in_aw_bits_id ? _aw_ready_WIRE_15 : _GEN_242; // @[src/main/scala/amba/axi4/UserYanker.scala 86:{36,36}]
  wire  line_245_clock;
  wire  line_245_reset;
  wire  line_245_valid;
  reg  line_245_valid_reg;
  wire  line_246_clock;
  wire  line_246_reset;
  wire  line_246_valid;
  reg  line_246_valid_reg;
  wire  line_247_clock;
  wire  line_247_reset;
  wire  line_247_valid;
  reg  line_247_valid_reg;
  wire  line_248_clock;
  wire  line_248_reset;
  wire  line_248_valid;
  reg  line_248_valid_reg;
  wire  line_249_clock;
  wire  line_249_reset;
  wire  line_249_valid;
  reg  line_249_valid_reg;
  wire  line_250_clock;
  wire  line_250_reset;
  wire  line_250_valid;
  reg  line_250_valid_reg;
  wire  line_251_clock;
  wire  line_251_reset;
  wire  line_251_valid;
  reg  line_251_valid_reg;
  wire  line_252_clock;
  wire  line_252_reset;
  wire  line_252_valid;
  reg  line_252_valid_reg;
  wire  line_253_clock;
  wire  line_253_reset;
  wire  line_253_valid;
  reg  line_253_valid_reg;
  wire  line_254_clock;
  wire  line_254_reset;
  wire  line_254_valid;
  reg  line_254_valid_reg;
  wire  line_255_clock;
  wire  line_255_reset;
  wire  line_255_valid;
  reg  line_255_valid_reg;
  wire  line_256_clock;
  wire  line_256_reset;
  wire  line_256_valid;
  reg  line_256_valid_reg;
  wire  line_257_clock;
  wire  line_257_reset;
  wire  line_257_valid;
  reg  line_257_valid_reg;
  wire  line_258_clock;
  wire  line_258_reset;
  wire  line_258_valid;
  reg  line_258_valid_reg;
  wire  line_259_clock;
  wire  line_259_reset;
  wire  line_259_valid;
  reg  line_259_valid_reg;
  wire  line_260_clock;
  wire  line_260_reset;
  wire  line_260_valid;
  reg  line_260_valid_reg;
  wire  line_261_clock;
  wire  line_261_reset;
  wire  line_261_valid;
  reg  line_261_valid_reg;
  wire  _b_valid_WIRE_0 = Queue_16_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  line_262_clock;
  wire  line_262_reset;
  wire  line_262_valid;
  reg  line_262_valid_reg;
  wire  _b_valid_WIRE_1 = Queue_17_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_245 = 4'h1 == auto_out_b_bits_id ? _b_valid_WIRE_1 : _b_valid_WIRE_0; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_263_clock;
  wire  line_263_reset;
  wire  line_263_valid;
  reg  line_263_valid_reg;
  wire  _b_valid_WIRE_2 = Queue_18_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_246 = 4'h2 == auto_out_b_bits_id ? _b_valid_WIRE_2 : _GEN_245; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_264_clock;
  wire  line_264_reset;
  wire  line_264_valid;
  reg  line_264_valid_reg;
  wire  _b_valid_WIRE_3 = Queue_19_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_247 = 4'h3 == auto_out_b_bits_id ? _b_valid_WIRE_3 : _GEN_246; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_265_clock;
  wire  line_265_reset;
  wire  line_265_valid;
  reg  line_265_valid_reg;
  wire  _b_valid_WIRE_4 = Queue_20_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_248 = 4'h4 == auto_out_b_bits_id ? _b_valid_WIRE_4 : _GEN_247; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_266_clock;
  wire  line_266_reset;
  wire  line_266_valid;
  reg  line_266_valid_reg;
  wire  _b_valid_WIRE_5 = Queue_21_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_249 = 4'h5 == auto_out_b_bits_id ? _b_valid_WIRE_5 : _GEN_248; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_267_clock;
  wire  line_267_reset;
  wire  line_267_valid;
  reg  line_267_valid_reg;
  wire  _b_valid_WIRE_6 = Queue_22_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_250 = 4'h6 == auto_out_b_bits_id ? _b_valid_WIRE_6 : _GEN_249; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_268_clock;
  wire  line_268_reset;
  wire  line_268_valid;
  reg  line_268_valid_reg;
  wire  _b_valid_WIRE_7 = Queue_23_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_251 = 4'h7 == auto_out_b_bits_id ? _b_valid_WIRE_7 : _GEN_250; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_269_clock;
  wire  line_269_reset;
  wire  line_269_valid;
  reg  line_269_valid_reg;
  wire  _b_valid_WIRE_8 = Queue_24_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_252 = 4'h8 == auto_out_b_bits_id ? _b_valid_WIRE_8 : _GEN_251; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_270_clock;
  wire  line_270_reset;
  wire  line_270_valid;
  reg  line_270_valid_reg;
  wire  _b_valid_WIRE_9 = Queue_25_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_253 = 4'h9 == auto_out_b_bits_id ? _b_valid_WIRE_9 : _GEN_252; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_271_clock;
  wire  line_271_reset;
  wire  line_271_valid;
  reg  line_271_valid_reg;
  wire  _b_valid_WIRE_10 = Queue_26_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_254 = 4'ha == auto_out_b_bits_id ? _b_valid_WIRE_10 : _GEN_253; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_272_clock;
  wire  line_272_reset;
  wire  line_272_valid;
  reg  line_272_valid_reg;
  wire  _b_valid_WIRE_11 = Queue_27_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_255 = 4'hb == auto_out_b_bits_id ? _b_valid_WIRE_11 : _GEN_254; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_273_clock;
  wire  line_273_reset;
  wire  line_273_valid;
  reg  line_273_valid_reg;
  wire  _b_valid_WIRE_12 = Queue_28_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_256 = 4'hc == auto_out_b_bits_id ? _b_valid_WIRE_12 : _GEN_255; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_274_clock;
  wire  line_274_reset;
  wire  line_274_valid;
  reg  line_274_valid_reg;
  wire  _b_valid_WIRE_13 = Queue_29_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_257 = 4'hd == auto_out_b_bits_id ? _b_valid_WIRE_13 : _GEN_256; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_275_clock;
  wire  line_275_reset;
  wire  line_275_valid;
  reg  line_275_valid_reg;
  wire  _b_valid_WIRE_14 = Queue_30_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_258 = 4'he == auto_out_b_bits_id ? _b_valid_WIRE_14 : _GEN_257; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_276_clock;
  wire  line_276_reset;
  wire  line_276_valid;
  reg  line_276_valid_reg;
  wire  _b_valid_WIRE_15 = Queue_31_io_deq_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 93:{28,28}]
  wire  _GEN_259 = 4'hf == auto_out_b_bits_id ? _b_valid_WIRE_15 : _GEN_258; // @[src/main/scala/amba/axi4/UserYanker.scala 95:{28,28}]
  wire  line_277_clock;
  wire  line_277_reset;
  wire  line_277_valid;
  reg  line_277_valid_reg;
  wire  _T_89 = ~(~auto_out_b_valid | _GEN_259); // @[src/main/scala/amba/axi4/UserYanker.scala 95:14]
  wire  line_278_clock;
  wire  line_278_reset;
  wire  line_278_valid;
  reg  line_278_valid_reg;
  wire  line_279_clock;
  wire  line_279_reset;
  wire  line_279_valid;
  reg  line_279_valid_reg;
  wire [3:0] _b_bits_WIRE_0_tl_state_source = Queue_16_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire  line_280_clock;
  wire  line_280_reset;
  wire  line_280_valid;
  reg  line_280_valid_reg;
  wire [3:0] _b_bits_WIRE_1_tl_state_source = Queue_17_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_261 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_tl_state_source : _b_bits_WIRE_0_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_281_clock;
  wire  line_281_reset;
  wire  line_281_valid;
  reg  line_281_valid_reg;
  wire [3:0] _b_bits_WIRE_2_tl_state_source = Queue_18_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_262 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_tl_state_source : _GEN_261; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_282_clock;
  wire  line_282_reset;
  wire  line_282_valid;
  reg  line_282_valid_reg;
  wire [3:0] _b_bits_WIRE_3_tl_state_source = Queue_19_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_263 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_tl_state_source : _GEN_262; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_283_clock;
  wire  line_283_reset;
  wire  line_283_valid;
  reg  line_283_valid_reg;
  wire [3:0] _b_bits_WIRE_4_tl_state_source = Queue_20_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_264 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_tl_state_source : _GEN_263; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_284_clock;
  wire  line_284_reset;
  wire  line_284_valid;
  reg  line_284_valid_reg;
  wire [3:0] _b_bits_WIRE_5_tl_state_source = Queue_21_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_265 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_tl_state_source : _GEN_264; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_285_clock;
  wire  line_285_reset;
  wire  line_285_valid;
  reg  line_285_valid_reg;
  wire [3:0] _b_bits_WIRE_6_tl_state_source = Queue_22_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_266 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_tl_state_source : _GEN_265; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_286_clock;
  wire  line_286_reset;
  wire  line_286_valid;
  reg  line_286_valid_reg;
  wire [3:0] _b_bits_WIRE_7_tl_state_source = Queue_23_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_267 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_tl_state_source : _GEN_266; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_287_clock;
  wire  line_287_reset;
  wire  line_287_valid;
  reg  line_287_valid_reg;
  wire [3:0] _b_bits_WIRE_8_tl_state_source = Queue_24_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_268 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_tl_state_source : _GEN_267; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_288_clock;
  wire  line_288_reset;
  wire  line_288_valid;
  reg  line_288_valid_reg;
  wire [3:0] _b_bits_WIRE_9_tl_state_source = Queue_25_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_269 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_tl_state_source : _GEN_268; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_289_clock;
  wire  line_289_reset;
  wire  line_289_valid;
  reg  line_289_valid_reg;
  wire [3:0] _b_bits_WIRE_10_tl_state_source = Queue_26_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_270 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_tl_state_source : _GEN_269; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_290_clock;
  wire  line_290_reset;
  wire  line_290_valid;
  reg  line_290_valid_reg;
  wire [3:0] _b_bits_WIRE_11_tl_state_source = Queue_27_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_271 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_tl_state_source : _GEN_270; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_291_clock;
  wire  line_291_reset;
  wire  line_291_valid;
  reg  line_291_valid_reg;
  wire [3:0] _b_bits_WIRE_12_tl_state_source = Queue_28_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_272 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_tl_state_source : _GEN_271; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_292_clock;
  wire  line_292_reset;
  wire  line_292_valid;
  reg  line_292_valid_reg;
  wire [3:0] _b_bits_WIRE_13_tl_state_source = Queue_29_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_273 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_tl_state_source : _GEN_272; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_293_clock;
  wire  line_293_reset;
  wire  line_293_valid;
  reg  line_293_valid_reg;
  wire [3:0] _b_bits_WIRE_14_tl_state_source = Queue_30_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_274 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_tl_state_source : _GEN_273; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_294_clock;
  wire  line_294_reset;
  wire  line_294_valid;
  reg  line_294_valid_reg;
  wire [3:0] _b_bits_WIRE_15_tl_state_source = Queue_31_io_deq_bits_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire  line_295_clock;
  wire  line_295_reset;
  wire  line_295_valid;
  reg  line_295_valid_reg;
  wire [3:0] _b_bits_WIRE_0_tl_state_size = Queue_16_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire  line_296_clock;
  wire  line_296_reset;
  wire  line_296_valid;
  reg  line_296_valid_reg;
  wire [3:0] _b_bits_WIRE_1_tl_state_size = Queue_17_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_277 = 4'h1 == auto_out_b_bits_id ? _b_bits_WIRE_1_tl_state_size : _b_bits_WIRE_0_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_297_clock;
  wire  line_297_reset;
  wire  line_297_valid;
  reg  line_297_valid_reg;
  wire [3:0] _b_bits_WIRE_2_tl_state_size = Queue_18_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_278 = 4'h2 == auto_out_b_bits_id ? _b_bits_WIRE_2_tl_state_size : _GEN_277; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_298_clock;
  wire  line_298_reset;
  wire  line_298_valid;
  reg  line_298_valid_reg;
  wire [3:0] _b_bits_WIRE_3_tl_state_size = Queue_19_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_279 = 4'h3 == auto_out_b_bits_id ? _b_bits_WIRE_3_tl_state_size : _GEN_278; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_299_clock;
  wire  line_299_reset;
  wire  line_299_valid;
  reg  line_299_valid_reg;
  wire [3:0] _b_bits_WIRE_4_tl_state_size = Queue_20_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_280 = 4'h4 == auto_out_b_bits_id ? _b_bits_WIRE_4_tl_state_size : _GEN_279; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_300_clock;
  wire  line_300_reset;
  wire  line_300_valid;
  reg  line_300_valid_reg;
  wire [3:0] _b_bits_WIRE_5_tl_state_size = Queue_21_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_281 = 4'h5 == auto_out_b_bits_id ? _b_bits_WIRE_5_tl_state_size : _GEN_280; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_301_clock;
  wire  line_301_reset;
  wire  line_301_valid;
  reg  line_301_valid_reg;
  wire [3:0] _b_bits_WIRE_6_tl_state_size = Queue_22_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_282 = 4'h6 == auto_out_b_bits_id ? _b_bits_WIRE_6_tl_state_size : _GEN_281; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_302_clock;
  wire  line_302_reset;
  wire  line_302_valid;
  reg  line_302_valid_reg;
  wire [3:0] _b_bits_WIRE_7_tl_state_size = Queue_23_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_283 = 4'h7 == auto_out_b_bits_id ? _b_bits_WIRE_7_tl_state_size : _GEN_282; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_303_clock;
  wire  line_303_reset;
  wire  line_303_valid;
  reg  line_303_valid_reg;
  wire [3:0] _b_bits_WIRE_8_tl_state_size = Queue_24_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_284 = 4'h8 == auto_out_b_bits_id ? _b_bits_WIRE_8_tl_state_size : _GEN_283; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_304_clock;
  wire  line_304_reset;
  wire  line_304_valid;
  reg  line_304_valid_reg;
  wire [3:0] _b_bits_WIRE_9_tl_state_size = Queue_25_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_285 = 4'h9 == auto_out_b_bits_id ? _b_bits_WIRE_9_tl_state_size : _GEN_284; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_305_clock;
  wire  line_305_reset;
  wire  line_305_valid;
  reg  line_305_valid_reg;
  wire [3:0] _b_bits_WIRE_10_tl_state_size = Queue_26_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_286 = 4'ha == auto_out_b_bits_id ? _b_bits_WIRE_10_tl_state_size : _GEN_285; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_306_clock;
  wire  line_306_reset;
  wire  line_306_valid;
  reg  line_306_valid_reg;
  wire [3:0] _b_bits_WIRE_11_tl_state_size = Queue_27_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_287 = 4'hb == auto_out_b_bits_id ? _b_bits_WIRE_11_tl_state_size : _GEN_286; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_307_clock;
  wire  line_307_reset;
  wire  line_307_valid;
  reg  line_307_valid_reg;
  wire [3:0] _b_bits_WIRE_12_tl_state_size = Queue_28_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_288 = 4'hc == auto_out_b_bits_id ? _b_bits_WIRE_12_tl_state_size : _GEN_287; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_308_clock;
  wire  line_308_reset;
  wire  line_308_valid;
  reg  line_308_valid_reg;
  wire [3:0] _b_bits_WIRE_13_tl_state_size = Queue_29_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_289 = 4'hd == auto_out_b_bits_id ? _b_bits_WIRE_13_tl_state_size : _GEN_288; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_309_clock;
  wire  line_309_reset;
  wire  line_309_valid;
  reg  line_309_valid_reg;
  wire [3:0] _b_bits_WIRE_14_tl_state_size = Queue_30_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [3:0] _GEN_290 = 4'he == auto_out_b_bits_id ? _b_bits_WIRE_14_tl_state_size : _GEN_289; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  wire  line_310_clock;
  wire  line_310_reset;
  wire  line_310_valid;
  reg  line_310_valid_reg;
  wire [3:0] _b_bits_WIRE_15_tl_state_size = Queue_31_io_deq_bits_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 94:{27,27}]
  wire [15:0] _awsel_T = 16'h1 << auto_in_aw_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  awsel_0 = _awsel_T[0]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_1 = _awsel_T[1]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_2 = _awsel_T[2]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_3 = _awsel_T[3]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_4 = _awsel_T[4]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_5 = _awsel_T[5]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_6 = _awsel_T[6]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_7 = _awsel_T[7]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_8 = _awsel_T[8]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_9 = _awsel_T[9]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_10 = _awsel_T[10]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_11 = _awsel_T[11]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_12 = _awsel_T[12]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_13 = _awsel_T[13]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_14 = _awsel_T[14]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire  awsel_15 = _awsel_T[15]; // @[src/main/scala/amba/axi4/UserYanker.scala 101:55]
  wire [15:0] _bsel_T = 16'h1 << auto_out_b_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  bsel_0 = _bsel_T[0]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_1 = _bsel_T[1]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_2 = _bsel_T[2]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_3 = _bsel_T[3]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_4 = _bsel_T[4]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_5 = _bsel_T[5]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_6 = _bsel_T[6]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_7 = _bsel_T[7]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_8 = _bsel_T[8]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_9 = _bsel_T[9]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_10 = _bsel_T[10]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_11 = _bsel_T[11]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_12 = _bsel_T[12]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_13 = _bsel_T[13]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_14 = _bsel_T[14]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  wire  bsel_15 = _bsel_T[15]; // @[src/main/scala/amba/axi4/UserYanker.scala 102:55]
  Queue_2 Queue ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_io_deq_bits_tl_state_source)
  );
  Queue_3 Queue_1 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_1_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_1_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_1_io_deq_bits_tl_state_source)
  );
  Queue_4 Queue_2 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_2_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_2_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_2_io_deq_bits_tl_state_source)
  );
  Queue_5 Queue_3 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_3_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_3_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_3_io_deq_bits_tl_state_source)
  );
  Queue_6 Queue_4 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_4_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_4_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_4_io_deq_bits_tl_state_source)
  );
  Queue_7 Queue_5 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_5_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_5_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_5_io_deq_bits_tl_state_source)
  );
  Queue_8 Queue_6 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_6_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_6_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_6_io_deq_bits_tl_state_source)
  );
  Queue_9 Queue_7 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_7_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_7_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_7_io_deq_bits_tl_state_source)
  );
  Queue_10 Queue_8 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_8_clock),
    .reset(Queue_8_reset),
    .io_enq_ready(Queue_8_io_enq_ready),
    .io_enq_valid(Queue_8_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_8_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_8_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_8_io_deq_ready),
    .io_deq_valid(Queue_8_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_8_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_8_io_deq_bits_tl_state_source)
  );
  Queue_11 Queue_9 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_9_clock),
    .reset(Queue_9_reset),
    .io_enq_ready(Queue_9_io_enq_ready),
    .io_enq_valid(Queue_9_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_9_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_9_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_9_io_deq_ready),
    .io_deq_valid(Queue_9_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_9_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_9_io_deq_bits_tl_state_source)
  );
  Queue_12 Queue_10 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_10_clock),
    .reset(Queue_10_reset),
    .io_enq_ready(Queue_10_io_enq_ready),
    .io_enq_valid(Queue_10_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_10_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_10_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_10_io_deq_ready),
    .io_deq_valid(Queue_10_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_10_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_10_io_deq_bits_tl_state_source)
  );
  Queue_13 Queue_11 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_11_clock),
    .reset(Queue_11_reset),
    .io_enq_ready(Queue_11_io_enq_ready),
    .io_enq_valid(Queue_11_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_11_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_11_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_11_io_deq_ready),
    .io_deq_valid(Queue_11_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_11_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_11_io_deq_bits_tl_state_source)
  );
  Queue_14 Queue_12 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_12_clock),
    .reset(Queue_12_reset),
    .io_enq_ready(Queue_12_io_enq_ready),
    .io_enq_valid(Queue_12_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_12_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_12_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_12_io_deq_ready),
    .io_deq_valid(Queue_12_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_12_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_12_io_deq_bits_tl_state_source)
  );
  Queue_15 Queue_13 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_13_clock),
    .reset(Queue_13_reset),
    .io_enq_ready(Queue_13_io_enq_ready),
    .io_enq_valid(Queue_13_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_13_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_13_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_13_io_deq_ready),
    .io_deq_valid(Queue_13_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_13_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_13_io_deq_bits_tl_state_source)
  );
  Queue_16 Queue_14 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_14_clock),
    .reset(Queue_14_reset),
    .io_enq_ready(Queue_14_io_enq_ready),
    .io_enq_valid(Queue_14_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_14_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_14_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_14_io_deq_ready),
    .io_deq_valid(Queue_14_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_14_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_14_io_deq_bits_tl_state_source)
  );
  Queue_17 Queue_15 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_15_clock),
    .reset(Queue_15_reset),
    .io_enq_ready(Queue_15_io_enq_ready),
    .io_enq_valid(Queue_15_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_15_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_15_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_15_io_deq_ready),
    .io_deq_valid(Queue_15_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_15_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_15_io_deq_bits_tl_state_source)
  );
  Queue_18 Queue_16 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_16_clock),
    .reset(Queue_16_reset),
    .io_enq_ready(Queue_16_io_enq_ready),
    .io_enq_valid(Queue_16_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_16_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_16_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_16_io_deq_ready),
    .io_deq_valid(Queue_16_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_16_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_16_io_deq_bits_tl_state_source)
  );
  Queue_19 Queue_17 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_17_clock),
    .reset(Queue_17_reset),
    .io_enq_ready(Queue_17_io_enq_ready),
    .io_enq_valid(Queue_17_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_17_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_17_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_17_io_deq_ready),
    .io_deq_valid(Queue_17_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_17_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_17_io_deq_bits_tl_state_source)
  );
  Queue_20 Queue_18 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_18_clock),
    .reset(Queue_18_reset),
    .io_enq_ready(Queue_18_io_enq_ready),
    .io_enq_valid(Queue_18_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_18_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_18_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_18_io_deq_ready),
    .io_deq_valid(Queue_18_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_18_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_18_io_deq_bits_tl_state_source)
  );
  Queue_21 Queue_19 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_19_clock),
    .reset(Queue_19_reset),
    .io_enq_ready(Queue_19_io_enq_ready),
    .io_enq_valid(Queue_19_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_19_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_19_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_19_io_deq_ready),
    .io_deq_valid(Queue_19_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_19_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_19_io_deq_bits_tl_state_source)
  );
  Queue_22 Queue_20 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_20_clock),
    .reset(Queue_20_reset),
    .io_enq_ready(Queue_20_io_enq_ready),
    .io_enq_valid(Queue_20_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_20_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_20_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_20_io_deq_ready),
    .io_deq_valid(Queue_20_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_20_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_20_io_deq_bits_tl_state_source)
  );
  Queue_23 Queue_21 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_21_clock),
    .reset(Queue_21_reset),
    .io_enq_ready(Queue_21_io_enq_ready),
    .io_enq_valid(Queue_21_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_21_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_21_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_21_io_deq_ready),
    .io_deq_valid(Queue_21_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_21_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_21_io_deq_bits_tl_state_source)
  );
  Queue_24 Queue_22 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_22_clock),
    .reset(Queue_22_reset),
    .io_enq_ready(Queue_22_io_enq_ready),
    .io_enq_valid(Queue_22_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_22_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_22_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_22_io_deq_ready),
    .io_deq_valid(Queue_22_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_22_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_22_io_deq_bits_tl_state_source)
  );
  Queue_25 Queue_23 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_23_clock),
    .reset(Queue_23_reset),
    .io_enq_ready(Queue_23_io_enq_ready),
    .io_enq_valid(Queue_23_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_23_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_23_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_23_io_deq_ready),
    .io_deq_valid(Queue_23_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_23_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_23_io_deq_bits_tl_state_source)
  );
  Queue_26 Queue_24 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_24_clock),
    .reset(Queue_24_reset),
    .io_enq_ready(Queue_24_io_enq_ready),
    .io_enq_valid(Queue_24_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_24_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_24_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_24_io_deq_ready),
    .io_deq_valid(Queue_24_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_24_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_24_io_deq_bits_tl_state_source)
  );
  Queue_27 Queue_25 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_25_clock),
    .reset(Queue_25_reset),
    .io_enq_ready(Queue_25_io_enq_ready),
    .io_enq_valid(Queue_25_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_25_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_25_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_25_io_deq_ready),
    .io_deq_valid(Queue_25_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_25_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_25_io_deq_bits_tl_state_source)
  );
  Queue_28 Queue_26 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_26_clock),
    .reset(Queue_26_reset),
    .io_enq_ready(Queue_26_io_enq_ready),
    .io_enq_valid(Queue_26_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_26_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_26_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_26_io_deq_ready),
    .io_deq_valid(Queue_26_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_26_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_26_io_deq_bits_tl_state_source)
  );
  Queue_29 Queue_27 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_27_clock),
    .reset(Queue_27_reset),
    .io_enq_ready(Queue_27_io_enq_ready),
    .io_enq_valid(Queue_27_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_27_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_27_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_27_io_deq_ready),
    .io_deq_valid(Queue_27_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_27_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_27_io_deq_bits_tl_state_source)
  );
  Queue_30 Queue_28 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_28_clock),
    .reset(Queue_28_reset),
    .io_enq_ready(Queue_28_io_enq_ready),
    .io_enq_valid(Queue_28_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_28_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_28_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_28_io_deq_ready),
    .io_deq_valid(Queue_28_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_28_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_28_io_deq_bits_tl_state_source)
  );
  Queue_31 Queue_29 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_29_clock),
    .reset(Queue_29_reset),
    .io_enq_ready(Queue_29_io_enq_ready),
    .io_enq_valid(Queue_29_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_29_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_29_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_29_io_deq_ready),
    .io_deq_valid(Queue_29_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_29_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_29_io_deq_bits_tl_state_source)
  );
  Queue_32 Queue_30 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_30_clock),
    .reset(Queue_30_reset),
    .io_enq_ready(Queue_30_io_enq_ready),
    .io_enq_valid(Queue_30_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_30_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_30_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_30_io_deq_ready),
    .io_deq_valid(Queue_30_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_30_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_30_io_deq_bits_tl_state_source)
  );
  Queue_33 Queue_31 ( // @[src/main/scala/amba/axi4/UserYanker.scala 48:17]
    .clock(Queue_31_clock),
    .reset(Queue_31_reset),
    .io_enq_ready(Queue_31_io_enq_ready),
    .io_enq_valid(Queue_31_io_enq_valid),
    .io_enq_bits_tl_state_size(Queue_31_io_enq_bits_tl_state_size),
    .io_enq_bits_tl_state_source(Queue_31_io_enq_bits_tl_state_source),
    .io_deq_ready(Queue_31_io_deq_ready),
    .io_deq_valid(Queue_31_io_deq_valid),
    .io_deq_bits_tl_state_size(Queue_31_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source(Queue_31_io_deq_bits_tl_state_source)
  );
  GEN_w1_line #(.COVER_INDEX(147)) line_147 (
    .clock(line_147_clock),
    .reset(line_147_reset),
    .valid(line_147_valid)
  );
  GEN_w1_line #(.COVER_INDEX(148)) line_148 (
    .clock(line_148_clock),
    .reset(line_148_reset),
    .valid(line_148_valid)
  );
  GEN_w1_line #(.COVER_INDEX(149)) line_149 (
    .clock(line_149_clock),
    .reset(line_149_reset),
    .valid(line_149_valid)
  );
  GEN_w1_line #(.COVER_INDEX(150)) line_150 (
    .clock(line_150_clock),
    .reset(line_150_reset),
    .valid(line_150_valid)
  );
  GEN_w1_line #(.COVER_INDEX(151)) line_151 (
    .clock(line_151_clock),
    .reset(line_151_reset),
    .valid(line_151_valid)
  );
  GEN_w1_line #(.COVER_INDEX(152)) line_152 (
    .clock(line_152_clock),
    .reset(line_152_reset),
    .valid(line_152_valid)
  );
  GEN_w1_line #(.COVER_INDEX(153)) line_153 (
    .clock(line_153_clock),
    .reset(line_153_reset),
    .valid(line_153_valid)
  );
  GEN_w1_line #(.COVER_INDEX(154)) line_154 (
    .clock(line_154_clock),
    .reset(line_154_reset),
    .valid(line_154_valid)
  );
  GEN_w1_line #(.COVER_INDEX(155)) line_155 (
    .clock(line_155_clock),
    .reset(line_155_reset),
    .valid(line_155_valid)
  );
  GEN_w1_line #(.COVER_INDEX(156)) line_156 (
    .clock(line_156_clock),
    .reset(line_156_reset),
    .valid(line_156_valid)
  );
  GEN_w1_line #(.COVER_INDEX(157)) line_157 (
    .clock(line_157_clock),
    .reset(line_157_reset),
    .valid(line_157_valid)
  );
  GEN_w1_line #(.COVER_INDEX(158)) line_158 (
    .clock(line_158_clock),
    .reset(line_158_reset),
    .valid(line_158_valid)
  );
  GEN_w1_line #(.COVER_INDEX(159)) line_159 (
    .clock(line_159_clock),
    .reset(line_159_reset),
    .valid(line_159_valid)
  );
  GEN_w1_line #(.COVER_INDEX(160)) line_160 (
    .clock(line_160_clock),
    .reset(line_160_reset),
    .valid(line_160_valid)
  );
  GEN_w1_line #(.COVER_INDEX(161)) line_161 (
    .clock(line_161_clock),
    .reset(line_161_reset),
    .valid(line_161_valid)
  );
  GEN_w1_line #(.COVER_INDEX(162)) line_162 (
    .clock(line_162_clock),
    .reset(line_162_reset),
    .valid(line_162_valid)
  );
  GEN_w1_line #(.COVER_INDEX(163)) line_163 (
    .clock(line_163_clock),
    .reset(line_163_reset),
    .valid(line_163_valid)
  );
  GEN_w1_line #(.COVER_INDEX(164)) line_164 (
    .clock(line_164_clock),
    .reset(line_164_reset),
    .valid(line_164_valid)
  );
  GEN_w1_line #(.COVER_INDEX(165)) line_165 (
    .clock(line_165_clock),
    .reset(line_165_reset),
    .valid(line_165_valid)
  );
  GEN_w1_line #(.COVER_INDEX(166)) line_166 (
    .clock(line_166_clock),
    .reset(line_166_reset),
    .valid(line_166_valid)
  );
  GEN_w1_line #(.COVER_INDEX(167)) line_167 (
    .clock(line_167_clock),
    .reset(line_167_reset),
    .valid(line_167_valid)
  );
  GEN_w1_line #(.COVER_INDEX(168)) line_168 (
    .clock(line_168_clock),
    .reset(line_168_reset),
    .valid(line_168_valid)
  );
  GEN_w1_line #(.COVER_INDEX(169)) line_169 (
    .clock(line_169_clock),
    .reset(line_169_reset),
    .valid(line_169_valid)
  );
  GEN_w1_line #(.COVER_INDEX(170)) line_170 (
    .clock(line_170_clock),
    .reset(line_170_reset),
    .valid(line_170_valid)
  );
  GEN_w1_line #(.COVER_INDEX(171)) line_171 (
    .clock(line_171_clock),
    .reset(line_171_reset),
    .valid(line_171_valid)
  );
  GEN_w1_line #(.COVER_INDEX(172)) line_172 (
    .clock(line_172_clock),
    .reset(line_172_reset),
    .valid(line_172_valid)
  );
  GEN_w1_line #(.COVER_INDEX(173)) line_173 (
    .clock(line_173_clock),
    .reset(line_173_reset),
    .valid(line_173_valid)
  );
  GEN_w1_line #(.COVER_INDEX(174)) line_174 (
    .clock(line_174_clock),
    .reset(line_174_reset),
    .valid(line_174_valid)
  );
  GEN_w1_line #(.COVER_INDEX(175)) line_175 (
    .clock(line_175_clock),
    .reset(line_175_reset),
    .valid(line_175_valid)
  );
  GEN_w1_line #(.COVER_INDEX(176)) line_176 (
    .clock(line_176_clock),
    .reset(line_176_reset),
    .valid(line_176_valid)
  );
  GEN_w1_line #(.COVER_INDEX(177)) line_177 (
    .clock(line_177_clock),
    .reset(line_177_reset),
    .valid(line_177_valid)
  );
  GEN_w1_line #(.COVER_INDEX(178)) line_178 (
    .clock(line_178_clock),
    .reset(line_178_reset),
    .valid(line_178_valid)
  );
  GEN_w1_line #(.COVER_INDEX(179)) line_179 (
    .clock(line_179_clock),
    .reset(line_179_reset),
    .valid(line_179_valid)
  );
  GEN_w1_line #(.COVER_INDEX(180)) line_180 (
    .clock(line_180_clock),
    .reset(line_180_reset),
    .valid(line_180_valid)
  );
  GEN_w1_line #(.COVER_INDEX(181)) line_181 (
    .clock(line_181_clock),
    .reset(line_181_reset),
    .valid(line_181_valid)
  );
  GEN_w1_line #(.COVER_INDEX(182)) line_182 (
    .clock(line_182_clock),
    .reset(line_182_reset),
    .valid(line_182_valid)
  );
  GEN_w1_line #(.COVER_INDEX(183)) line_183 (
    .clock(line_183_clock),
    .reset(line_183_reset),
    .valid(line_183_valid)
  );
  GEN_w1_line #(.COVER_INDEX(184)) line_184 (
    .clock(line_184_clock),
    .reset(line_184_reset),
    .valid(line_184_valid)
  );
  GEN_w1_line #(.COVER_INDEX(185)) line_185 (
    .clock(line_185_clock),
    .reset(line_185_reset),
    .valid(line_185_valid)
  );
  GEN_w1_line #(.COVER_INDEX(186)) line_186 (
    .clock(line_186_clock),
    .reset(line_186_reset),
    .valid(line_186_valid)
  );
  GEN_w1_line #(.COVER_INDEX(187)) line_187 (
    .clock(line_187_clock),
    .reset(line_187_reset),
    .valid(line_187_valid)
  );
  GEN_w1_line #(.COVER_INDEX(188)) line_188 (
    .clock(line_188_clock),
    .reset(line_188_reset),
    .valid(line_188_valid)
  );
  GEN_w1_line #(.COVER_INDEX(189)) line_189 (
    .clock(line_189_clock),
    .reset(line_189_reset),
    .valid(line_189_valid)
  );
  GEN_w1_line #(.COVER_INDEX(190)) line_190 (
    .clock(line_190_clock),
    .reset(line_190_reset),
    .valid(line_190_valid)
  );
  GEN_w1_line #(.COVER_INDEX(191)) line_191 (
    .clock(line_191_clock),
    .reset(line_191_reset),
    .valid(line_191_valid)
  );
  GEN_w1_line #(.COVER_INDEX(192)) line_192 (
    .clock(line_192_clock),
    .reset(line_192_reset),
    .valid(line_192_valid)
  );
  GEN_w1_line #(.COVER_INDEX(193)) line_193 (
    .clock(line_193_clock),
    .reset(line_193_reset),
    .valid(line_193_valid)
  );
  GEN_w1_line #(.COVER_INDEX(194)) line_194 (
    .clock(line_194_clock),
    .reset(line_194_reset),
    .valid(line_194_valid)
  );
  GEN_w1_line #(.COVER_INDEX(195)) line_195 (
    .clock(line_195_clock),
    .reset(line_195_reset),
    .valid(line_195_valid)
  );
  GEN_w1_line #(.COVER_INDEX(196)) line_196 (
    .clock(line_196_clock),
    .reset(line_196_reset),
    .valid(line_196_valid)
  );
  GEN_w1_line #(.COVER_INDEX(197)) line_197 (
    .clock(line_197_clock),
    .reset(line_197_reset),
    .valid(line_197_valid)
  );
  GEN_w1_line #(.COVER_INDEX(198)) line_198 (
    .clock(line_198_clock),
    .reset(line_198_reset),
    .valid(line_198_valid)
  );
  GEN_w1_line #(.COVER_INDEX(199)) line_199 (
    .clock(line_199_clock),
    .reset(line_199_reset),
    .valid(line_199_valid)
  );
  GEN_w1_line #(.COVER_INDEX(200)) line_200 (
    .clock(line_200_clock),
    .reset(line_200_reset),
    .valid(line_200_valid)
  );
  GEN_w1_line #(.COVER_INDEX(201)) line_201 (
    .clock(line_201_clock),
    .reset(line_201_reset),
    .valid(line_201_valid)
  );
  GEN_w1_line #(.COVER_INDEX(202)) line_202 (
    .clock(line_202_clock),
    .reset(line_202_reset),
    .valid(line_202_valid)
  );
  GEN_w1_line #(.COVER_INDEX(203)) line_203 (
    .clock(line_203_clock),
    .reset(line_203_reset),
    .valid(line_203_valid)
  );
  GEN_w1_line #(.COVER_INDEX(204)) line_204 (
    .clock(line_204_clock),
    .reset(line_204_reset),
    .valid(line_204_valid)
  );
  GEN_w1_line #(.COVER_INDEX(205)) line_205 (
    .clock(line_205_clock),
    .reset(line_205_reset),
    .valid(line_205_valid)
  );
  GEN_w1_line #(.COVER_INDEX(206)) line_206 (
    .clock(line_206_clock),
    .reset(line_206_reset),
    .valid(line_206_valid)
  );
  GEN_w1_line #(.COVER_INDEX(207)) line_207 (
    .clock(line_207_clock),
    .reset(line_207_reset),
    .valid(line_207_valid)
  );
  GEN_w1_line #(.COVER_INDEX(208)) line_208 (
    .clock(line_208_clock),
    .reset(line_208_reset),
    .valid(line_208_valid)
  );
  GEN_w1_line #(.COVER_INDEX(209)) line_209 (
    .clock(line_209_clock),
    .reset(line_209_reset),
    .valid(line_209_valid)
  );
  GEN_w1_line #(.COVER_INDEX(210)) line_210 (
    .clock(line_210_clock),
    .reset(line_210_reset),
    .valid(line_210_valid)
  );
  GEN_w1_line #(.COVER_INDEX(211)) line_211 (
    .clock(line_211_clock),
    .reset(line_211_reset),
    .valid(line_211_valid)
  );
  GEN_w1_line #(.COVER_INDEX(212)) line_212 (
    .clock(line_212_clock),
    .reset(line_212_reset),
    .valid(line_212_valid)
  );
  GEN_w1_line #(.COVER_INDEX(213)) line_213 (
    .clock(line_213_clock),
    .reset(line_213_reset),
    .valid(line_213_valid)
  );
  GEN_w1_line #(.COVER_INDEX(214)) line_214 (
    .clock(line_214_clock),
    .reset(line_214_reset),
    .valid(line_214_valid)
  );
  GEN_w1_line #(.COVER_INDEX(215)) line_215 (
    .clock(line_215_clock),
    .reset(line_215_reset),
    .valid(line_215_valid)
  );
  GEN_w1_line #(.COVER_INDEX(216)) line_216 (
    .clock(line_216_clock),
    .reset(line_216_reset),
    .valid(line_216_valid)
  );
  GEN_w1_line #(.COVER_INDEX(217)) line_217 (
    .clock(line_217_clock),
    .reset(line_217_reset),
    .valid(line_217_valid)
  );
  GEN_w1_line #(.COVER_INDEX(218)) line_218 (
    .clock(line_218_clock),
    .reset(line_218_reset),
    .valid(line_218_valid)
  );
  GEN_w1_line #(.COVER_INDEX(219)) line_219 (
    .clock(line_219_clock),
    .reset(line_219_reset),
    .valid(line_219_valid)
  );
  GEN_w1_line #(.COVER_INDEX(220)) line_220 (
    .clock(line_220_clock),
    .reset(line_220_reset),
    .valid(line_220_valid)
  );
  GEN_w1_line #(.COVER_INDEX(221)) line_221 (
    .clock(line_221_clock),
    .reset(line_221_reset),
    .valid(line_221_valid)
  );
  GEN_w1_line #(.COVER_INDEX(222)) line_222 (
    .clock(line_222_clock),
    .reset(line_222_reset),
    .valid(line_222_valid)
  );
  GEN_w1_line #(.COVER_INDEX(223)) line_223 (
    .clock(line_223_clock),
    .reset(line_223_reset),
    .valid(line_223_valid)
  );
  GEN_w1_line #(.COVER_INDEX(224)) line_224 (
    .clock(line_224_clock),
    .reset(line_224_reset),
    .valid(line_224_valid)
  );
  GEN_w1_line #(.COVER_INDEX(225)) line_225 (
    .clock(line_225_clock),
    .reset(line_225_reset),
    .valid(line_225_valid)
  );
  GEN_w1_line #(.COVER_INDEX(226)) line_226 (
    .clock(line_226_clock),
    .reset(line_226_reset),
    .valid(line_226_valid)
  );
  GEN_w1_line #(.COVER_INDEX(227)) line_227 (
    .clock(line_227_clock),
    .reset(line_227_reset),
    .valid(line_227_valid)
  );
  GEN_w1_line #(.COVER_INDEX(228)) line_228 (
    .clock(line_228_clock),
    .reset(line_228_reset),
    .valid(line_228_valid)
  );
  GEN_w1_line #(.COVER_INDEX(229)) line_229 (
    .clock(line_229_clock),
    .reset(line_229_reset),
    .valid(line_229_valid)
  );
  GEN_w1_line #(.COVER_INDEX(230)) line_230 (
    .clock(line_230_clock),
    .reset(line_230_reset),
    .valid(line_230_valid)
  );
  GEN_w1_line #(.COVER_INDEX(231)) line_231 (
    .clock(line_231_clock),
    .reset(line_231_reset),
    .valid(line_231_valid)
  );
  GEN_w1_line #(.COVER_INDEX(232)) line_232 (
    .clock(line_232_clock),
    .reset(line_232_reset),
    .valid(line_232_valid)
  );
  GEN_w1_line #(.COVER_INDEX(233)) line_233 (
    .clock(line_233_clock),
    .reset(line_233_reset),
    .valid(line_233_valid)
  );
  GEN_w1_line #(.COVER_INDEX(234)) line_234 (
    .clock(line_234_clock),
    .reset(line_234_reset),
    .valid(line_234_valid)
  );
  GEN_w1_line #(.COVER_INDEX(235)) line_235 (
    .clock(line_235_clock),
    .reset(line_235_reset),
    .valid(line_235_valid)
  );
  GEN_w1_line #(.COVER_INDEX(236)) line_236 (
    .clock(line_236_clock),
    .reset(line_236_reset),
    .valid(line_236_valid)
  );
  GEN_w1_line #(.COVER_INDEX(237)) line_237 (
    .clock(line_237_clock),
    .reset(line_237_reset),
    .valid(line_237_valid)
  );
  GEN_w1_line #(.COVER_INDEX(238)) line_238 (
    .clock(line_238_clock),
    .reset(line_238_reset),
    .valid(line_238_valid)
  );
  GEN_w1_line #(.COVER_INDEX(239)) line_239 (
    .clock(line_239_clock),
    .reset(line_239_reset),
    .valid(line_239_valid)
  );
  GEN_w1_line #(.COVER_INDEX(240)) line_240 (
    .clock(line_240_clock),
    .reset(line_240_reset),
    .valid(line_240_valid)
  );
  GEN_w1_line #(.COVER_INDEX(241)) line_241 (
    .clock(line_241_clock),
    .reset(line_241_reset),
    .valid(line_241_valid)
  );
  GEN_w1_line #(.COVER_INDEX(242)) line_242 (
    .clock(line_242_clock),
    .reset(line_242_reset),
    .valid(line_242_valid)
  );
  GEN_w1_line #(.COVER_INDEX(243)) line_243 (
    .clock(line_243_clock),
    .reset(line_243_reset),
    .valid(line_243_valid)
  );
  GEN_w1_line #(.COVER_INDEX(244)) line_244 (
    .clock(line_244_clock),
    .reset(line_244_reset),
    .valid(line_244_valid)
  );
  GEN_w1_line #(.COVER_INDEX(245)) line_245 (
    .clock(line_245_clock),
    .reset(line_245_reset),
    .valid(line_245_valid)
  );
  GEN_w1_line #(.COVER_INDEX(246)) line_246 (
    .clock(line_246_clock),
    .reset(line_246_reset),
    .valid(line_246_valid)
  );
  GEN_w1_line #(.COVER_INDEX(247)) line_247 (
    .clock(line_247_clock),
    .reset(line_247_reset),
    .valid(line_247_valid)
  );
  GEN_w1_line #(.COVER_INDEX(248)) line_248 (
    .clock(line_248_clock),
    .reset(line_248_reset),
    .valid(line_248_valid)
  );
  GEN_w1_line #(.COVER_INDEX(249)) line_249 (
    .clock(line_249_clock),
    .reset(line_249_reset),
    .valid(line_249_valid)
  );
  GEN_w1_line #(.COVER_INDEX(250)) line_250 (
    .clock(line_250_clock),
    .reset(line_250_reset),
    .valid(line_250_valid)
  );
  GEN_w1_line #(.COVER_INDEX(251)) line_251 (
    .clock(line_251_clock),
    .reset(line_251_reset),
    .valid(line_251_valid)
  );
  GEN_w1_line #(.COVER_INDEX(252)) line_252 (
    .clock(line_252_clock),
    .reset(line_252_reset),
    .valid(line_252_valid)
  );
  GEN_w1_line #(.COVER_INDEX(253)) line_253 (
    .clock(line_253_clock),
    .reset(line_253_reset),
    .valid(line_253_valid)
  );
  GEN_w1_line #(.COVER_INDEX(254)) line_254 (
    .clock(line_254_clock),
    .reset(line_254_reset),
    .valid(line_254_valid)
  );
  GEN_w1_line #(.COVER_INDEX(255)) line_255 (
    .clock(line_255_clock),
    .reset(line_255_reset),
    .valid(line_255_valid)
  );
  GEN_w1_line #(.COVER_INDEX(256)) line_256 (
    .clock(line_256_clock),
    .reset(line_256_reset),
    .valid(line_256_valid)
  );
  GEN_w1_line #(.COVER_INDEX(257)) line_257 (
    .clock(line_257_clock),
    .reset(line_257_reset),
    .valid(line_257_valid)
  );
  GEN_w1_line #(.COVER_INDEX(258)) line_258 (
    .clock(line_258_clock),
    .reset(line_258_reset),
    .valid(line_258_valid)
  );
  GEN_w1_line #(.COVER_INDEX(259)) line_259 (
    .clock(line_259_clock),
    .reset(line_259_reset),
    .valid(line_259_valid)
  );
  GEN_w1_line #(.COVER_INDEX(260)) line_260 (
    .clock(line_260_clock),
    .reset(line_260_reset),
    .valid(line_260_valid)
  );
  GEN_w1_line #(.COVER_INDEX(261)) line_261 (
    .clock(line_261_clock),
    .reset(line_261_reset),
    .valid(line_261_valid)
  );
  GEN_w1_line #(.COVER_INDEX(262)) line_262 (
    .clock(line_262_clock),
    .reset(line_262_reset),
    .valid(line_262_valid)
  );
  GEN_w1_line #(.COVER_INDEX(263)) line_263 (
    .clock(line_263_clock),
    .reset(line_263_reset),
    .valid(line_263_valid)
  );
  GEN_w1_line #(.COVER_INDEX(264)) line_264 (
    .clock(line_264_clock),
    .reset(line_264_reset),
    .valid(line_264_valid)
  );
  GEN_w1_line #(.COVER_INDEX(265)) line_265 (
    .clock(line_265_clock),
    .reset(line_265_reset),
    .valid(line_265_valid)
  );
  GEN_w1_line #(.COVER_INDEX(266)) line_266 (
    .clock(line_266_clock),
    .reset(line_266_reset),
    .valid(line_266_valid)
  );
  GEN_w1_line #(.COVER_INDEX(267)) line_267 (
    .clock(line_267_clock),
    .reset(line_267_reset),
    .valid(line_267_valid)
  );
  GEN_w1_line #(.COVER_INDEX(268)) line_268 (
    .clock(line_268_clock),
    .reset(line_268_reset),
    .valid(line_268_valid)
  );
  GEN_w1_line #(.COVER_INDEX(269)) line_269 (
    .clock(line_269_clock),
    .reset(line_269_reset),
    .valid(line_269_valid)
  );
  GEN_w1_line #(.COVER_INDEX(270)) line_270 (
    .clock(line_270_clock),
    .reset(line_270_reset),
    .valid(line_270_valid)
  );
  GEN_w1_line #(.COVER_INDEX(271)) line_271 (
    .clock(line_271_clock),
    .reset(line_271_reset),
    .valid(line_271_valid)
  );
  GEN_w1_line #(.COVER_INDEX(272)) line_272 (
    .clock(line_272_clock),
    .reset(line_272_reset),
    .valid(line_272_valid)
  );
  GEN_w1_line #(.COVER_INDEX(273)) line_273 (
    .clock(line_273_clock),
    .reset(line_273_reset),
    .valid(line_273_valid)
  );
  GEN_w1_line #(.COVER_INDEX(274)) line_274 (
    .clock(line_274_clock),
    .reset(line_274_reset),
    .valid(line_274_valid)
  );
  GEN_w1_line #(.COVER_INDEX(275)) line_275 (
    .clock(line_275_clock),
    .reset(line_275_reset),
    .valid(line_275_valid)
  );
  GEN_w1_line #(.COVER_INDEX(276)) line_276 (
    .clock(line_276_clock),
    .reset(line_276_reset),
    .valid(line_276_valid)
  );
  GEN_w1_line #(.COVER_INDEX(277)) line_277 (
    .clock(line_277_clock),
    .reset(line_277_reset),
    .valid(line_277_valid)
  );
  GEN_w1_line #(.COVER_INDEX(278)) line_278 (
    .clock(line_278_clock),
    .reset(line_278_reset),
    .valid(line_278_valid)
  );
  GEN_w1_line #(.COVER_INDEX(279)) line_279 (
    .clock(line_279_clock),
    .reset(line_279_reset),
    .valid(line_279_valid)
  );
  GEN_w1_line #(.COVER_INDEX(280)) line_280 (
    .clock(line_280_clock),
    .reset(line_280_reset),
    .valid(line_280_valid)
  );
  GEN_w1_line #(.COVER_INDEX(281)) line_281 (
    .clock(line_281_clock),
    .reset(line_281_reset),
    .valid(line_281_valid)
  );
  GEN_w1_line #(.COVER_INDEX(282)) line_282 (
    .clock(line_282_clock),
    .reset(line_282_reset),
    .valid(line_282_valid)
  );
  GEN_w1_line #(.COVER_INDEX(283)) line_283 (
    .clock(line_283_clock),
    .reset(line_283_reset),
    .valid(line_283_valid)
  );
  GEN_w1_line #(.COVER_INDEX(284)) line_284 (
    .clock(line_284_clock),
    .reset(line_284_reset),
    .valid(line_284_valid)
  );
  GEN_w1_line #(.COVER_INDEX(285)) line_285 (
    .clock(line_285_clock),
    .reset(line_285_reset),
    .valid(line_285_valid)
  );
  GEN_w1_line #(.COVER_INDEX(286)) line_286 (
    .clock(line_286_clock),
    .reset(line_286_reset),
    .valid(line_286_valid)
  );
  GEN_w1_line #(.COVER_INDEX(287)) line_287 (
    .clock(line_287_clock),
    .reset(line_287_reset),
    .valid(line_287_valid)
  );
  GEN_w1_line #(.COVER_INDEX(288)) line_288 (
    .clock(line_288_clock),
    .reset(line_288_reset),
    .valid(line_288_valid)
  );
  GEN_w1_line #(.COVER_INDEX(289)) line_289 (
    .clock(line_289_clock),
    .reset(line_289_reset),
    .valid(line_289_valid)
  );
  GEN_w1_line #(.COVER_INDEX(290)) line_290 (
    .clock(line_290_clock),
    .reset(line_290_reset),
    .valid(line_290_valid)
  );
  GEN_w1_line #(.COVER_INDEX(291)) line_291 (
    .clock(line_291_clock),
    .reset(line_291_reset),
    .valid(line_291_valid)
  );
  GEN_w1_line #(.COVER_INDEX(292)) line_292 (
    .clock(line_292_clock),
    .reset(line_292_reset),
    .valid(line_292_valid)
  );
  GEN_w1_line #(.COVER_INDEX(293)) line_293 (
    .clock(line_293_clock),
    .reset(line_293_reset),
    .valid(line_293_valid)
  );
  GEN_w1_line #(.COVER_INDEX(294)) line_294 (
    .clock(line_294_clock),
    .reset(line_294_reset),
    .valid(line_294_valid)
  );
  GEN_w1_line #(.COVER_INDEX(295)) line_295 (
    .clock(line_295_clock),
    .reset(line_295_reset),
    .valid(line_295_valid)
  );
  GEN_w1_line #(.COVER_INDEX(296)) line_296 (
    .clock(line_296_clock),
    .reset(line_296_reset),
    .valid(line_296_valid)
  );
  GEN_w1_line #(.COVER_INDEX(297)) line_297 (
    .clock(line_297_clock),
    .reset(line_297_reset),
    .valid(line_297_valid)
  );
  GEN_w1_line #(.COVER_INDEX(298)) line_298 (
    .clock(line_298_clock),
    .reset(line_298_reset),
    .valid(line_298_valid)
  );
  GEN_w1_line #(.COVER_INDEX(299)) line_299 (
    .clock(line_299_clock),
    .reset(line_299_reset),
    .valid(line_299_valid)
  );
  GEN_w1_line #(.COVER_INDEX(300)) line_300 (
    .clock(line_300_clock),
    .reset(line_300_reset),
    .valid(line_300_valid)
  );
  GEN_w1_line #(.COVER_INDEX(301)) line_301 (
    .clock(line_301_clock),
    .reset(line_301_reset),
    .valid(line_301_valid)
  );
  GEN_w1_line #(.COVER_INDEX(302)) line_302 (
    .clock(line_302_clock),
    .reset(line_302_reset),
    .valid(line_302_valid)
  );
  GEN_w1_line #(.COVER_INDEX(303)) line_303 (
    .clock(line_303_clock),
    .reset(line_303_reset),
    .valid(line_303_valid)
  );
  GEN_w1_line #(.COVER_INDEX(304)) line_304 (
    .clock(line_304_clock),
    .reset(line_304_reset),
    .valid(line_304_valid)
  );
  GEN_w1_line #(.COVER_INDEX(305)) line_305 (
    .clock(line_305_clock),
    .reset(line_305_reset),
    .valid(line_305_valid)
  );
  GEN_w1_line #(.COVER_INDEX(306)) line_306 (
    .clock(line_306_clock),
    .reset(line_306_reset),
    .valid(line_306_valid)
  );
  GEN_w1_line #(.COVER_INDEX(307)) line_307 (
    .clock(line_307_clock),
    .reset(line_307_reset),
    .valid(line_307_valid)
  );
  GEN_w1_line #(.COVER_INDEX(308)) line_308 (
    .clock(line_308_clock),
    .reset(line_308_reset),
    .valid(line_308_valid)
  );
  GEN_w1_line #(.COVER_INDEX(309)) line_309 (
    .clock(line_309_clock),
    .reset(line_309_reset),
    .valid(line_309_valid)
  );
  GEN_w1_line #(.COVER_INDEX(310)) line_310 (
    .clock(line_310_clock),
    .reset(line_310_reset),
    .valid(line_310_valid)
  );
  assign line_147_clock = clock;
  assign line_147_reset = reset;
  assign line_147_valid = 4'h0 == auto_in_ar_bits_id ^ line_147_valid_reg;
  assign line_148_clock = clock;
  assign line_148_reset = reset;
  assign line_148_valid = 4'h1 == auto_in_ar_bits_id ^ line_148_valid_reg;
  assign line_149_clock = clock;
  assign line_149_reset = reset;
  assign line_149_valid = 4'h2 == auto_in_ar_bits_id ^ line_149_valid_reg;
  assign line_150_clock = clock;
  assign line_150_reset = reset;
  assign line_150_valid = 4'h3 == auto_in_ar_bits_id ^ line_150_valid_reg;
  assign line_151_clock = clock;
  assign line_151_reset = reset;
  assign line_151_valid = 4'h4 == auto_in_ar_bits_id ^ line_151_valid_reg;
  assign line_152_clock = clock;
  assign line_152_reset = reset;
  assign line_152_valid = 4'h5 == auto_in_ar_bits_id ^ line_152_valid_reg;
  assign line_153_clock = clock;
  assign line_153_reset = reset;
  assign line_153_valid = 4'h6 == auto_in_ar_bits_id ^ line_153_valid_reg;
  assign line_154_clock = clock;
  assign line_154_reset = reset;
  assign line_154_valid = 4'h7 == auto_in_ar_bits_id ^ line_154_valid_reg;
  assign line_155_clock = clock;
  assign line_155_reset = reset;
  assign line_155_valid = 4'h8 == auto_in_ar_bits_id ^ line_155_valid_reg;
  assign line_156_clock = clock;
  assign line_156_reset = reset;
  assign line_156_valid = 4'h9 == auto_in_ar_bits_id ^ line_156_valid_reg;
  assign line_157_clock = clock;
  assign line_157_reset = reset;
  assign line_157_valid = 4'ha == auto_in_ar_bits_id ^ line_157_valid_reg;
  assign line_158_clock = clock;
  assign line_158_reset = reset;
  assign line_158_valid = 4'hb == auto_in_ar_bits_id ^ line_158_valid_reg;
  assign line_159_clock = clock;
  assign line_159_reset = reset;
  assign line_159_valid = 4'hc == auto_in_ar_bits_id ^ line_159_valid_reg;
  assign line_160_clock = clock;
  assign line_160_reset = reset;
  assign line_160_valid = 4'hd == auto_in_ar_bits_id ^ line_160_valid_reg;
  assign line_161_clock = clock;
  assign line_161_reset = reset;
  assign line_161_valid = 4'he == auto_in_ar_bits_id ^ line_161_valid_reg;
  assign line_162_clock = clock;
  assign line_162_reset = reset;
  assign line_162_valid = 4'hf == auto_in_ar_bits_id ^ line_162_valid_reg;
  assign line_163_clock = clock;
  assign line_163_reset = reset;
  assign line_163_valid = 4'h0 == auto_in_ar_bits_id ^ line_163_valid_reg;
  assign line_164_clock = clock;
  assign line_164_reset = reset;
  assign line_164_valid = 4'h1 == auto_in_ar_bits_id ^ line_164_valid_reg;
  assign line_165_clock = clock;
  assign line_165_reset = reset;
  assign line_165_valid = 4'h2 == auto_in_ar_bits_id ^ line_165_valid_reg;
  assign line_166_clock = clock;
  assign line_166_reset = reset;
  assign line_166_valid = 4'h3 == auto_in_ar_bits_id ^ line_166_valid_reg;
  assign line_167_clock = clock;
  assign line_167_reset = reset;
  assign line_167_valid = 4'h4 == auto_in_ar_bits_id ^ line_167_valid_reg;
  assign line_168_clock = clock;
  assign line_168_reset = reset;
  assign line_168_valid = 4'h5 == auto_in_ar_bits_id ^ line_168_valid_reg;
  assign line_169_clock = clock;
  assign line_169_reset = reset;
  assign line_169_valid = 4'h6 == auto_in_ar_bits_id ^ line_169_valid_reg;
  assign line_170_clock = clock;
  assign line_170_reset = reset;
  assign line_170_valid = 4'h7 == auto_in_ar_bits_id ^ line_170_valid_reg;
  assign line_171_clock = clock;
  assign line_171_reset = reset;
  assign line_171_valid = 4'h8 == auto_in_ar_bits_id ^ line_171_valid_reg;
  assign line_172_clock = clock;
  assign line_172_reset = reset;
  assign line_172_valid = 4'h9 == auto_in_ar_bits_id ^ line_172_valid_reg;
  assign line_173_clock = clock;
  assign line_173_reset = reset;
  assign line_173_valid = 4'ha == auto_in_ar_bits_id ^ line_173_valid_reg;
  assign line_174_clock = clock;
  assign line_174_reset = reset;
  assign line_174_valid = 4'hb == auto_in_ar_bits_id ^ line_174_valid_reg;
  assign line_175_clock = clock;
  assign line_175_reset = reset;
  assign line_175_valid = 4'hc == auto_in_ar_bits_id ^ line_175_valid_reg;
  assign line_176_clock = clock;
  assign line_176_reset = reset;
  assign line_176_valid = 4'hd == auto_in_ar_bits_id ^ line_176_valid_reg;
  assign line_177_clock = clock;
  assign line_177_reset = reset;
  assign line_177_valid = 4'he == auto_in_ar_bits_id ^ line_177_valid_reg;
  assign line_178_clock = clock;
  assign line_178_reset = reset;
  assign line_178_valid = 4'hf == auto_in_ar_bits_id ^ line_178_valid_reg;
  assign line_179_clock = clock;
  assign line_179_reset = reset;
  assign line_179_valid = 4'h0 == auto_out_r_bits_id ^ line_179_valid_reg;
  assign line_180_clock = clock;
  assign line_180_reset = reset;
  assign line_180_valid = 4'h1 == auto_out_r_bits_id ^ line_180_valid_reg;
  assign line_181_clock = clock;
  assign line_181_reset = reset;
  assign line_181_valid = 4'h2 == auto_out_r_bits_id ^ line_181_valid_reg;
  assign line_182_clock = clock;
  assign line_182_reset = reset;
  assign line_182_valid = 4'h3 == auto_out_r_bits_id ^ line_182_valid_reg;
  assign line_183_clock = clock;
  assign line_183_reset = reset;
  assign line_183_valid = 4'h4 == auto_out_r_bits_id ^ line_183_valid_reg;
  assign line_184_clock = clock;
  assign line_184_reset = reset;
  assign line_184_valid = 4'h5 == auto_out_r_bits_id ^ line_184_valid_reg;
  assign line_185_clock = clock;
  assign line_185_reset = reset;
  assign line_185_valid = 4'h6 == auto_out_r_bits_id ^ line_185_valid_reg;
  assign line_186_clock = clock;
  assign line_186_reset = reset;
  assign line_186_valid = 4'h7 == auto_out_r_bits_id ^ line_186_valid_reg;
  assign line_187_clock = clock;
  assign line_187_reset = reset;
  assign line_187_valid = 4'h8 == auto_out_r_bits_id ^ line_187_valid_reg;
  assign line_188_clock = clock;
  assign line_188_reset = reset;
  assign line_188_valid = 4'h9 == auto_out_r_bits_id ^ line_188_valid_reg;
  assign line_189_clock = clock;
  assign line_189_reset = reset;
  assign line_189_valid = 4'ha == auto_out_r_bits_id ^ line_189_valid_reg;
  assign line_190_clock = clock;
  assign line_190_reset = reset;
  assign line_190_valid = 4'hb == auto_out_r_bits_id ^ line_190_valid_reg;
  assign line_191_clock = clock;
  assign line_191_reset = reset;
  assign line_191_valid = 4'hc == auto_out_r_bits_id ^ line_191_valid_reg;
  assign line_192_clock = clock;
  assign line_192_reset = reset;
  assign line_192_valid = 4'hd == auto_out_r_bits_id ^ line_192_valid_reg;
  assign line_193_clock = clock;
  assign line_193_reset = reset;
  assign line_193_valid = 4'he == auto_out_r_bits_id ^ line_193_valid_reg;
  assign line_194_clock = clock;
  assign line_194_reset = reset;
  assign line_194_valid = 4'hf == auto_out_r_bits_id ^ line_194_valid_reg;
  assign line_195_clock = clock;
  assign line_195_reset = reset;
  assign line_195_valid = _T_3 ^ line_195_valid_reg;
  assign line_196_clock = clock;
  assign line_196_reset = reset;
  assign line_196_valid = _T_4 ^ line_196_valid_reg;
  assign line_197_clock = clock;
  assign line_197_reset = reset;
  assign line_197_valid = 4'h0 == auto_out_r_bits_id ^ line_197_valid_reg;
  assign line_198_clock = clock;
  assign line_198_reset = reset;
  assign line_198_valid = 4'h1 == auto_out_r_bits_id ^ line_198_valid_reg;
  assign line_199_clock = clock;
  assign line_199_reset = reset;
  assign line_199_valid = 4'h2 == auto_out_r_bits_id ^ line_199_valid_reg;
  assign line_200_clock = clock;
  assign line_200_reset = reset;
  assign line_200_valid = 4'h3 == auto_out_r_bits_id ^ line_200_valid_reg;
  assign line_201_clock = clock;
  assign line_201_reset = reset;
  assign line_201_valid = 4'h4 == auto_out_r_bits_id ^ line_201_valid_reg;
  assign line_202_clock = clock;
  assign line_202_reset = reset;
  assign line_202_valid = 4'h5 == auto_out_r_bits_id ^ line_202_valid_reg;
  assign line_203_clock = clock;
  assign line_203_reset = reset;
  assign line_203_valid = 4'h6 == auto_out_r_bits_id ^ line_203_valid_reg;
  assign line_204_clock = clock;
  assign line_204_reset = reset;
  assign line_204_valid = 4'h7 == auto_out_r_bits_id ^ line_204_valid_reg;
  assign line_205_clock = clock;
  assign line_205_reset = reset;
  assign line_205_valid = 4'h8 == auto_out_r_bits_id ^ line_205_valid_reg;
  assign line_206_clock = clock;
  assign line_206_reset = reset;
  assign line_206_valid = 4'h9 == auto_out_r_bits_id ^ line_206_valid_reg;
  assign line_207_clock = clock;
  assign line_207_reset = reset;
  assign line_207_valid = 4'ha == auto_out_r_bits_id ^ line_207_valid_reg;
  assign line_208_clock = clock;
  assign line_208_reset = reset;
  assign line_208_valid = 4'hb == auto_out_r_bits_id ^ line_208_valid_reg;
  assign line_209_clock = clock;
  assign line_209_reset = reset;
  assign line_209_valid = 4'hc == auto_out_r_bits_id ^ line_209_valid_reg;
  assign line_210_clock = clock;
  assign line_210_reset = reset;
  assign line_210_valid = 4'hd == auto_out_r_bits_id ^ line_210_valid_reg;
  assign line_211_clock = clock;
  assign line_211_reset = reset;
  assign line_211_valid = 4'he == auto_out_r_bits_id ^ line_211_valid_reg;
  assign line_212_clock = clock;
  assign line_212_reset = reset;
  assign line_212_valid = 4'hf == auto_out_r_bits_id ^ line_212_valid_reg;
  assign line_213_clock = clock;
  assign line_213_reset = reset;
  assign line_213_valid = 4'h0 == auto_out_r_bits_id ^ line_213_valid_reg;
  assign line_214_clock = clock;
  assign line_214_reset = reset;
  assign line_214_valid = 4'h1 == auto_out_r_bits_id ^ line_214_valid_reg;
  assign line_215_clock = clock;
  assign line_215_reset = reset;
  assign line_215_valid = 4'h2 == auto_out_r_bits_id ^ line_215_valid_reg;
  assign line_216_clock = clock;
  assign line_216_reset = reset;
  assign line_216_valid = 4'h3 == auto_out_r_bits_id ^ line_216_valid_reg;
  assign line_217_clock = clock;
  assign line_217_reset = reset;
  assign line_217_valid = 4'h4 == auto_out_r_bits_id ^ line_217_valid_reg;
  assign line_218_clock = clock;
  assign line_218_reset = reset;
  assign line_218_valid = 4'h5 == auto_out_r_bits_id ^ line_218_valid_reg;
  assign line_219_clock = clock;
  assign line_219_reset = reset;
  assign line_219_valid = 4'h6 == auto_out_r_bits_id ^ line_219_valid_reg;
  assign line_220_clock = clock;
  assign line_220_reset = reset;
  assign line_220_valid = 4'h7 == auto_out_r_bits_id ^ line_220_valid_reg;
  assign line_221_clock = clock;
  assign line_221_reset = reset;
  assign line_221_valid = 4'h8 == auto_out_r_bits_id ^ line_221_valid_reg;
  assign line_222_clock = clock;
  assign line_222_reset = reset;
  assign line_222_valid = 4'h9 == auto_out_r_bits_id ^ line_222_valid_reg;
  assign line_223_clock = clock;
  assign line_223_reset = reset;
  assign line_223_valid = 4'ha == auto_out_r_bits_id ^ line_223_valid_reg;
  assign line_224_clock = clock;
  assign line_224_reset = reset;
  assign line_224_valid = 4'hb == auto_out_r_bits_id ^ line_224_valid_reg;
  assign line_225_clock = clock;
  assign line_225_reset = reset;
  assign line_225_valid = 4'hc == auto_out_r_bits_id ^ line_225_valid_reg;
  assign line_226_clock = clock;
  assign line_226_reset = reset;
  assign line_226_valid = 4'hd == auto_out_r_bits_id ^ line_226_valid_reg;
  assign line_227_clock = clock;
  assign line_227_reset = reset;
  assign line_227_valid = 4'he == auto_out_r_bits_id ^ line_227_valid_reg;
  assign line_228_clock = clock;
  assign line_228_reset = reset;
  assign line_228_valid = 4'hf == auto_out_r_bits_id ^ line_228_valid_reg;
  assign line_229_clock = clock;
  assign line_229_reset = reset;
  assign line_229_valid = 4'h0 == auto_in_aw_bits_id ^ line_229_valid_reg;
  assign line_230_clock = clock;
  assign line_230_reset = reset;
  assign line_230_valid = 4'h1 == auto_in_aw_bits_id ^ line_230_valid_reg;
  assign line_231_clock = clock;
  assign line_231_reset = reset;
  assign line_231_valid = 4'h2 == auto_in_aw_bits_id ^ line_231_valid_reg;
  assign line_232_clock = clock;
  assign line_232_reset = reset;
  assign line_232_valid = 4'h3 == auto_in_aw_bits_id ^ line_232_valid_reg;
  assign line_233_clock = clock;
  assign line_233_reset = reset;
  assign line_233_valid = 4'h4 == auto_in_aw_bits_id ^ line_233_valid_reg;
  assign line_234_clock = clock;
  assign line_234_reset = reset;
  assign line_234_valid = 4'h5 == auto_in_aw_bits_id ^ line_234_valid_reg;
  assign line_235_clock = clock;
  assign line_235_reset = reset;
  assign line_235_valid = 4'h6 == auto_in_aw_bits_id ^ line_235_valid_reg;
  assign line_236_clock = clock;
  assign line_236_reset = reset;
  assign line_236_valid = 4'h7 == auto_in_aw_bits_id ^ line_236_valid_reg;
  assign line_237_clock = clock;
  assign line_237_reset = reset;
  assign line_237_valid = 4'h8 == auto_in_aw_bits_id ^ line_237_valid_reg;
  assign line_238_clock = clock;
  assign line_238_reset = reset;
  assign line_238_valid = 4'h9 == auto_in_aw_bits_id ^ line_238_valid_reg;
  assign line_239_clock = clock;
  assign line_239_reset = reset;
  assign line_239_valid = 4'ha == auto_in_aw_bits_id ^ line_239_valid_reg;
  assign line_240_clock = clock;
  assign line_240_reset = reset;
  assign line_240_valid = 4'hb == auto_in_aw_bits_id ^ line_240_valid_reg;
  assign line_241_clock = clock;
  assign line_241_reset = reset;
  assign line_241_valid = 4'hc == auto_in_aw_bits_id ^ line_241_valid_reg;
  assign line_242_clock = clock;
  assign line_242_reset = reset;
  assign line_242_valid = 4'hd == auto_in_aw_bits_id ^ line_242_valid_reg;
  assign line_243_clock = clock;
  assign line_243_reset = reset;
  assign line_243_valid = 4'he == auto_in_aw_bits_id ^ line_243_valid_reg;
  assign line_244_clock = clock;
  assign line_244_reset = reset;
  assign line_244_valid = 4'hf == auto_in_aw_bits_id ^ line_244_valid_reg;
  assign line_245_clock = clock;
  assign line_245_reset = reset;
  assign line_245_valid = 4'h0 == auto_in_aw_bits_id ^ line_245_valid_reg;
  assign line_246_clock = clock;
  assign line_246_reset = reset;
  assign line_246_valid = 4'h1 == auto_in_aw_bits_id ^ line_246_valid_reg;
  assign line_247_clock = clock;
  assign line_247_reset = reset;
  assign line_247_valid = 4'h2 == auto_in_aw_bits_id ^ line_247_valid_reg;
  assign line_248_clock = clock;
  assign line_248_reset = reset;
  assign line_248_valid = 4'h3 == auto_in_aw_bits_id ^ line_248_valid_reg;
  assign line_249_clock = clock;
  assign line_249_reset = reset;
  assign line_249_valid = 4'h4 == auto_in_aw_bits_id ^ line_249_valid_reg;
  assign line_250_clock = clock;
  assign line_250_reset = reset;
  assign line_250_valid = 4'h5 == auto_in_aw_bits_id ^ line_250_valid_reg;
  assign line_251_clock = clock;
  assign line_251_reset = reset;
  assign line_251_valid = 4'h6 == auto_in_aw_bits_id ^ line_251_valid_reg;
  assign line_252_clock = clock;
  assign line_252_reset = reset;
  assign line_252_valid = 4'h7 == auto_in_aw_bits_id ^ line_252_valid_reg;
  assign line_253_clock = clock;
  assign line_253_reset = reset;
  assign line_253_valid = 4'h8 == auto_in_aw_bits_id ^ line_253_valid_reg;
  assign line_254_clock = clock;
  assign line_254_reset = reset;
  assign line_254_valid = 4'h9 == auto_in_aw_bits_id ^ line_254_valid_reg;
  assign line_255_clock = clock;
  assign line_255_reset = reset;
  assign line_255_valid = 4'ha == auto_in_aw_bits_id ^ line_255_valid_reg;
  assign line_256_clock = clock;
  assign line_256_reset = reset;
  assign line_256_valid = 4'hb == auto_in_aw_bits_id ^ line_256_valid_reg;
  assign line_257_clock = clock;
  assign line_257_reset = reset;
  assign line_257_valid = 4'hc == auto_in_aw_bits_id ^ line_257_valid_reg;
  assign line_258_clock = clock;
  assign line_258_reset = reset;
  assign line_258_valid = 4'hd == auto_in_aw_bits_id ^ line_258_valid_reg;
  assign line_259_clock = clock;
  assign line_259_reset = reset;
  assign line_259_valid = 4'he == auto_in_aw_bits_id ^ line_259_valid_reg;
  assign line_260_clock = clock;
  assign line_260_reset = reset;
  assign line_260_valid = 4'hf == auto_in_aw_bits_id ^ line_260_valid_reg;
  assign line_261_clock = clock;
  assign line_261_reset = reset;
  assign line_261_valid = 4'h0 == auto_out_b_bits_id ^ line_261_valid_reg;
  assign line_262_clock = clock;
  assign line_262_reset = reset;
  assign line_262_valid = 4'h1 == auto_out_b_bits_id ^ line_262_valid_reg;
  assign line_263_clock = clock;
  assign line_263_reset = reset;
  assign line_263_valid = 4'h2 == auto_out_b_bits_id ^ line_263_valid_reg;
  assign line_264_clock = clock;
  assign line_264_reset = reset;
  assign line_264_valid = 4'h3 == auto_out_b_bits_id ^ line_264_valid_reg;
  assign line_265_clock = clock;
  assign line_265_reset = reset;
  assign line_265_valid = 4'h4 == auto_out_b_bits_id ^ line_265_valid_reg;
  assign line_266_clock = clock;
  assign line_266_reset = reset;
  assign line_266_valid = 4'h5 == auto_out_b_bits_id ^ line_266_valid_reg;
  assign line_267_clock = clock;
  assign line_267_reset = reset;
  assign line_267_valid = 4'h6 == auto_out_b_bits_id ^ line_267_valid_reg;
  assign line_268_clock = clock;
  assign line_268_reset = reset;
  assign line_268_valid = 4'h7 == auto_out_b_bits_id ^ line_268_valid_reg;
  assign line_269_clock = clock;
  assign line_269_reset = reset;
  assign line_269_valid = 4'h8 == auto_out_b_bits_id ^ line_269_valid_reg;
  assign line_270_clock = clock;
  assign line_270_reset = reset;
  assign line_270_valid = 4'h9 == auto_out_b_bits_id ^ line_270_valid_reg;
  assign line_271_clock = clock;
  assign line_271_reset = reset;
  assign line_271_valid = 4'ha == auto_out_b_bits_id ^ line_271_valid_reg;
  assign line_272_clock = clock;
  assign line_272_reset = reset;
  assign line_272_valid = 4'hb == auto_out_b_bits_id ^ line_272_valid_reg;
  assign line_273_clock = clock;
  assign line_273_reset = reset;
  assign line_273_valid = 4'hc == auto_out_b_bits_id ^ line_273_valid_reg;
  assign line_274_clock = clock;
  assign line_274_reset = reset;
  assign line_274_valid = 4'hd == auto_out_b_bits_id ^ line_274_valid_reg;
  assign line_275_clock = clock;
  assign line_275_reset = reset;
  assign line_275_valid = 4'he == auto_out_b_bits_id ^ line_275_valid_reg;
  assign line_276_clock = clock;
  assign line_276_reset = reset;
  assign line_276_valid = 4'hf == auto_out_b_bits_id ^ line_276_valid_reg;
  assign line_277_clock = clock;
  assign line_277_reset = reset;
  assign line_277_valid = _T_3 ^ line_277_valid_reg;
  assign line_278_clock = clock;
  assign line_278_reset = reset;
  assign line_278_valid = _T_89 ^ line_278_valid_reg;
  assign line_279_clock = clock;
  assign line_279_reset = reset;
  assign line_279_valid = 4'h0 == auto_out_b_bits_id ^ line_279_valid_reg;
  assign line_280_clock = clock;
  assign line_280_reset = reset;
  assign line_280_valid = 4'h1 == auto_out_b_bits_id ^ line_280_valid_reg;
  assign line_281_clock = clock;
  assign line_281_reset = reset;
  assign line_281_valid = 4'h2 == auto_out_b_bits_id ^ line_281_valid_reg;
  assign line_282_clock = clock;
  assign line_282_reset = reset;
  assign line_282_valid = 4'h3 == auto_out_b_bits_id ^ line_282_valid_reg;
  assign line_283_clock = clock;
  assign line_283_reset = reset;
  assign line_283_valid = 4'h4 == auto_out_b_bits_id ^ line_283_valid_reg;
  assign line_284_clock = clock;
  assign line_284_reset = reset;
  assign line_284_valid = 4'h5 == auto_out_b_bits_id ^ line_284_valid_reg;
  assign line_285_clock = clock;
  assign line_285_reset = reset;
  assign line_285_valid = 4'h6 == auto_out_b_bits_id ^ line_285_valid_reg;
  assign line_286_clock = clock;
  assign line_286_reset = reset;
  assign line_286_valid = 4'h7 == auto_out_b_bits_id ^ line_286_valid_reg;
  assign line_287_clock = clock;
  assign line_287_reset = reset;
  assign line_287_valid = 4'h8 == auto_out_b_bits_id ^ line_287_valid_reg;
  assign line_288_clock = clock;
  assign line_288_reset = reset;
  assign line_288_valid = 4'h9 == auto_out_b_bits_id ^ line_288_valid_reg;
  assign line_289_clock = clock;
  assign line_289_reset = reset;
  assign line_289_valid = 4'ha == auto_out_b_bits_id ^ line_289_valid_reg;
  assign line_290_clock = clock;
  assign line_290_reset = reset;
  assign line_290_valid = 4'hb == auto_out_b_bits_id ^ line_290_valid_reg;
  assign line_291_clock = clock;
  assign line_291_reset = reset;
  assign line_291_valid = 4'hc == auto_out_b_bits_id ^ line_291_valid_reg;
  assign line_292_clock = clock;
  assign line_292_reset = reset;
  assign line_292_valid = 4'hd == auto_out_b_bits_id ^ line_292_valid_reg;
  assign line_293_clock = clock;
  assign line_293_reset = reset;
  assign line_293_valid = 4'he == auto_out_b_bits_id ^ line_293_valid_reg;
  assign line_294_clock = clock;
  assign line_294_reset = reset;
  assign line_294_valid = 4'hf == auto_out_b_bits_id ^ line_294_valid_reg;
  assign line_295_clock = clock;
  assign line_295_reset = reset;
  assign line_295_valid = 4'h0 == auto_out_b_bits_id ^ line_295_valid_reg;
  assign line_296_clock = clock;
  assign line_296_reset = reset;
  assign line_296_valid = 4'h1 == auto_out_b_bits_id ^ line_296_valid_reg;
  assign line_297_clock = clock;
  assign line_297_reset = reset;
  assign line_297_valid = 4'h2 == auto_out_b_bits_id ^ line_297_valid_reg;
  assign line_298_clock = clock;
  assign line_298_reset = reset;
  assign line_298_valid = 4'h3 == auto_out_b_bits_id ^ line_298_valid_reg;
  assign line_299_clock = clock;
  assign line_299_reset = reset;
  assign line_299_valid = 4'h4 == auto_out_b_bits_id ^ line_299_valid_reg;
  assign line_300_clock = clock;
  assign line_300_reset = reset;
  assign line_300_valid = 4'h5 == auto_out_b_bits_id ^ line_300_valid_reg;
  assign line_301_clock = clock;
  assign line_301_reset = reset;
  assign line_301_valid = 4'h6 == auto_out_b_bits_id ^ line_301_valid_reg;
  assign line_302_clock = clock;
  assign line_302_reset = reset;
  assign line_302_valid = 4'h7 == auto_out_b_bits_id ^ line_302_valid_reg;
  assign line_303_clock = clock;
  assign line_303_reset = reset;
  assign line_303_valid = 4'h8 == auto_out_b_bits_id ^ line_303_valid_reg;
  assign line_304_clock = clock;
  assign line_304_reset = reset;
  assign line_304_valid = 4'h9 == auto_out_b_bits_id ^ line_304_valid_reg;
  assign line_305_clock = clock;
  assign line_305_reset = reset;
  assign line_305_valid = 4'ha == auto_out_b_bits_id ^ line_305_valid_reg;
  assign line_306_clock = clock;
  assign line_306_reset = reset;
  assign line_306_valid = 4'hb == auto_out_b_bits_id ^ line_306_valid_reg;
  assign line_307_clock = clock;
  assign line_307_reset = reset;
  assign line_307_valid = 4'hc == auto_out_b_bits_id ^ line_307_valid_reg;
  assign line_308_clock = clock;
  assign line_308_reset = reset;
  assign line_308_valid = 4'hd == auto_out_b_bits_id ^ line_308_valid_reg;
  assign line_309_clock = clock;
  assign line_309_reset = reset;
  assign line_309_valid = 4'he == auto_out_b_bits_id ^ line_309_valid_reg;
  assign line_310_clock = clock;
  assign line_310_reset = reset;
  assign line_310_valid = 4'hf == auto_out_b_bits_id ^ line_310_valid_reg;
  assign auto_in_aw_ready = auto_out_aw_ready & _GEN_243; // @[src/main/scala/amba/axi4/UserYanker.scala 86:36]
  assign auto_in_w_ready = auto_out_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_echo_tl_state_size = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_tl_state_size : _GEN_290; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  assign auto_in_b_bits_echo_tl_state_source = 4'hf == auto_out_b_bits_id ? _b_bits_WIRE_15_tl_state_source : _GEN_274; // @[src/main/scala/amba/axi4/UserYanker.scala 99:{22,22}]
  assign auto_in_ar_ready = auto_out_ar_ready & _GEN_179; // @[src/main/scala/amba/axi4/UserYanker.scala 57:36]
  assign auto_in_r_valid = auto_out_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_echo_tl_state_size = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_tl_state_size : _GEN_226; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  assign auto_in_r_bits_echo_tl_state_source = 4'hf == auto_out_r_bits_id ? _r_bits_WIRE_15_tl_state_source : _GEN_210; // @[src/main/scala/amba/axi4/UserYanker.scala 70:{22,22}]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_aw_valid = auto_in_aw_valid & _GEN_243; // @[src/main/scala/amba/axi4/UserYanker.scala 87:36]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_valid = auto_in_ar_valid & _GEN_179; // @[src/main/scala/amba/axi4/UserYanker.scala 58:36]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_0; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_0 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_1; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_1_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_1_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_1_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_1 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_2; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_2_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_2_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_2_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_2 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_3; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_3_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_3_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_3_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_3 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_4; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_4_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_4_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_4_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_4 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_5; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_5_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_5_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_5_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_5 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_6_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_6; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_6_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_6_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_6_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_6 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_7_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_7; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_7_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_7_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_7_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_7 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_8_clock = clock;
  assign Queue_8_reset = reset;
  assign Queue_8_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_8; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_8_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_8_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_8_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_8 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_9_clock = clock;
  assign Queue_9_reset = reset;
  assign Queue_9_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_9; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_9_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_9_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_9_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_9 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_10_clock = clock;
  assign Queue_10_reset = reset;
  assign Queue_10_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_10; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_10_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_10_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_10_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_10 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_11_clock = clock;
  assign Queue_11_reset = reset;
  assign Queue_11_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_11; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_11_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_11_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_11_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_11 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_12_clock = clock;
  assign Queue_12_reset = reset;
  assign Queue_12_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_12; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_12_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_12_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_12_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_12 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_13_clock = clock;
  assign Queue_13_reset = reset;
  assign Queue_13_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_13; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_13_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_13_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_13_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_13 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_14_clock = clock;
  assign Queue_14_reset = reset;
  assign Queue_14_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_14; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_14_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_14_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_14_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_14 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_15_clock = clock;
  assign Queue_15_reset = reset;
  assign Queue_15_io_enq_valid = auto_in_ar_valid & auto_out_ar_ready & arsel_15; // @[src/main/scala/amba/axi4/UserYanker.scala 78:53]
  assign Queue_15_io_enq_bits_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_15_io_enq_bits_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_15_io_deq_ready = auto_out_r_valid & auto_in_r_ready & rsel_15 & auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 75:58]
  assign Queue_16_clock = clock;
  assign Queue_16_reset = reset;
  assign Queue_16_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_0; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_16_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_16_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_16_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_0; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_17_clock = clock;
  assign Queue_17_reset = reset;
  assign Queue_17_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_1; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_17_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_17_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_17_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_1; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_18_clock = clock;
  assign Queue_18_reset = reset;
  assign Queue_18_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_2; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_18_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_18_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_18_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_2; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_19_clock = clock;
  assign Queue_19_reset = reset;
  assign Queue_19_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_3; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_19_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_19_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_19_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_3; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_20_clock = clock;
  assign Queue_20_reset = reset;
  assign Queue_20_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_4; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_20_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_20_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_20_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_4; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_21_clock = clock;
  assign Queue_21_reset = reset;
  assign Queue_21_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_5; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_21_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_21_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_21_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_5; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_22_clock = clock;
  assign Queue_22_reset = reset;
  assign Queue_22_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_6; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_22_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_22_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_22_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_6; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_23_clock = clock;
  assign Queue_23_reset = reset;
  assign Queue_23_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_7; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_23_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_23_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_23_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_7; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_24_clock = clock;
  assign Queue_24_reset = reset;
  assign Queue_24_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_8; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_24_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_24_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_24_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_8; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_25_clock = clock;
  assign Queue_25_reset = reset;
  assign Queue_25_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_9; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_25_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_25_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_25_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_9; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_26_clock = clock;
  assign Queue_26_reset = reset;
  assign Queue_26_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_10; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_26_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_26_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_26_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_10; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_27_clock = clock;
  assign Queue_27_reset = reset;
  assign Queue_27_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_11; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_27_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_27_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_27_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_11; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_28_clock = clock;
  assign Queue_28_reset = reset;
  assign Queue_28_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_12; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_28_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_28_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_28_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_12; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_29_clock = clock;
  assign Queue_29_reset = reset;
  assign Queue_29_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_13; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_29_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_29_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_29_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_13; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_30_clock = clock;
  assign Queue_30_reset = reset;
  assign Queue_30_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_14; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_30_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_30_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_30_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_14; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  assign Queue_31_clock = clock;
  assign Queue_31_reset = reset;
  assign Queue_31_io_enq_valid = auto_in_aw_valid & auto_out_aw_ready & awsel_15; // @[src/main/scala/amba/axi4/UserYanker.scala 107:53]
  assign Queue_31_io_enq_bits_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_31_io_enq_bits_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign Queue_31_io_deq_ready = auto_out_b_valid & auto_in_b_ready & bsel_15; // @[src/main/scala/amba/axi4/UserYanker.scala 104:53]
  always @(posedge clock) begin
    line_147_valid_reg <= 4'h0 == auto_in_ar_bits_id;
    line_148_valid_reg <= 4'h1 == auto_in_ar_bits_id;
    line_149_valid_reg <= 4'h2 == auto_in_ar_bits_id;
    line_150_valid_reg <= 4'h3 == auto_in_ar_bits_id;
    line_151_valid_reg <= 4'h4 == auto_in_ar_bits_id;
    line_152_valid_reg <= 4'h5 == auto_in_ar_bits_id;
    line_153_valid_reg <= 4'h6 == auto_in_ar_bits_id;
    line_154_valid_reg <= 4'h7 == auto_in_ar_bits_id;
    line_155_valid_reg <= 4'h8 == auto_in_ar_bits_id;
    line_156_valid_reg <= 4'h9 == auto_in_ar_bits_id;
    line_157_valid_reg <= 4'ha == auto_in_ar_bits_id;
    line_158_valid_reg <= 4'hb == auto_in_ar_bits_id;
    line_159_valid_reg <= 4'hc == auto_in_ar_bits_id;
    line_160_valid_reg <= 4'hd == auto_in_ar_bits_id;
    line_161_valid_reg <= 4'he == auto_in_ar_bits_id;
    line_162_valid_reg <= 4'hf == auto_in_ar_bits_id;
    line_163_valid_reg <= 4'h0 == auto_in_ar_bits_id;
    line_164_valid_reg <= 4'h1 == auto_in_ar_bits_id;
    line_165_valid_reg <= 4'h2 == auto_in_ar_bits_id;
    line_166_valid_reg <= 4'h3 == auto_in_ar_bits_id;
    line_167_valid_reg <= 4'h4 == auto_in_ar_bits_id;
    line_168_valid_reg <= 4'h5 == auto_in_ar_bits_id;
    line_169_valid_reg <= 4'h6 == auto_in_ar_bits_id;
    line_170_valid_reg <= 4'h7 == auto_in_ar_bits_id;
    line_171_valid_reg <= 4'h8 == auto_in_ar_bits_id;
    line_172_valid_reg <= 4'h9 == auto_in_ar_bits_id;
    line_173_valid_reg <= 4'ha == auto_in_ar_bits_id;
    line_174_valid_reg <= 4'hb == auto_in_ar_bits_id;
    line_175_valid_reg <= 4'hc == auto_in_ar_bits_id;
    line_176_valid_reg <= 4'hd == auto_in_ar_bits_id;
    line_177_valid_reg <= 4'he == auto_in_ar_bits_id;
    line_178_valid_reg <= 4'hf == auto_in_ar_bits_id;
    line_179_valid_reg <= 4'h0 == auto_out_r_bits_id;
    line_180_valid_reg <= 4'h1 == auto_out_r_bits_id;
    line_181_valid_reg <= 4'h2 == auto_out_r_bits_id;
    line_182_valid_reg <= 4'h3 == auto_out_r_bits_id;
    line_183_valid_reg <= 4'h4 == auto_out_r_bits_id;
    line_184_valid_reg <= 4'h5 == auto_out_r_bits_id;
    line_185_valid_reg <= 4'h6 == auto_out_r_bits_id;
    line_186_valid_reg <= 4'h7 == auto_out_r_bits_id;
    line_187_valid_reg <= 4'h8 == auto_out_r_bits_id;
    line_188_valid_reg <= 4'h9 == auto_out_r_bits_id;
    line_189_valid_reg <= 4'ha == auto_out_r_bits_id;
    line_190_valid_reg <= 4'hb == auto_out_r_bits_id;
    line_191_valid_reg <= 4'hc == auto_out_r_bits_id;
    line_192_valid_reg <= 4'hd == auto_out_r_bits_id;
    line_193_valid_reg <= 4'he == auto_out_r_bits_id;
    line_194_valid_reg <= 4'hf == auto_out_r_bits_id;
    line_195_valid_reg <= _T_3;
    line_196_valid_reg <= _T_4;
    line_197_valid_reg <= 4'h0 == auto_out_r_bits_id;
    line_198_valid_reg <= 4'h1 == auto_out_r_bits_id;
    line_199_valid_reg <= 4'h2 == auto_out_r_bits_id;
    line_200_valid_reg <= 4'h3 == auto_out_r_bits_id;
    line_201_valid_reg <= 4'h4 == auto_out_r_bits_id;
    line_202_valid_reg <= 4'h5 == auto_out_r_bits_id;
    line_203_valid_reg <= 4'h6 == auto_out_r_bits_id;
    line_204_valid_reg <= 4'h7 == auto_out_r_bits_id;
    line_205_valid_reg <= 4'h8 == auto_out_r_bits_id;
    line_206_valid_reg <= 4'h9 == auto_out_r_bits_id;
    line_207_valid_reg <= 4'ha == auto_out_r_bits_id;
    line_208_valid_reg <= 4'hb == auto_out_r_bits_id;
    line_209_valid_reg <= 4'hc == auto_out_r_bits_id;
    line_210_valid_reg <= 4'hd == auto_out_r_bits_id;
    line_211_valid_reg <= 4'he == auto_out_r_bits_id;
    line_212_valid_reg <= 4'hf == auto_out_r_bits_id;
    line_213_valid_reg <= 4'h0 == auto_out_r_bits_id;
    line_214_valid_reg <= 4'h1 == auto_out_r_bits_id;
    line_215_valid_reg <= 4'h2 == auto_out_r_bits_id;
    line_216_valid_reg <= 4'h3 == auto_out_r_bits_id;
    line_217_valid_reg <= 4'h4 == auto_out_r_bits_id;
    line_218_valid_reg <= 4'h5 == auto_out_r_bits_id;
    line_219_valid_reg <= 4'h6 == auto_out_r_bits_id;
    line_220_valid_reg <= 4'h7 == auto_out_r_bits_id;
    line_221_valid_reg <= 4'h8 == auto_out_r_bits_id;
    line_222_valid_reg <= 4'h9 == auto_out_r_bits_id;
    line_223_valid_reg <= 4'ha == auto_out_r_bits_id;
    line_224_valid_reg <= 4'hb == auto_out_r_bits_id;
    line_225_valid_reg <= 4'hc == auto_out_r_bits_id;
    line_226_valid_reg <= 4'hd == auto_out_r_bits_id;
    line_227_valid_reg <= 4'he == auto_out_r_bits_id;
    line_228_valid_reg <= 4'hf == auto_out_r_bits_id;
    line_229_valid_reg <= 4'h0 == auto_in_aw_bits_id;
    line_230_valid_reg <= 4'h1 == auto_in_aw_bits_id;
    line_231_valid_reg <= 4'h2 == auto_in_aw_bits_id;
    line_232_valid_reg <= 4'h3 == auto_in_aw_bits_id;
    line_233_valid_reg <= 4'h4 == auto_in_aw_bits_id;
    line_234_valid_reg <= 4'h5 == auto_in_aw_bits_id;
    line_235_valid_reg <= 4'h6 == auto_in_aw_bits_id;
    line_236_valid_reg <= 4'h7 == auto_in_aw_bits_id;
    line_237_valid_reg <= 4'h8 == auto_in_aw_bits_id;
    line_238_valid_reg <= 4'h9 == auto_in_aw_bits_id;
    line_239_valid_reg <= 4'ha == auto_in_aw_bits_id;
    line_240_valid_reg <= 4'hb == auto_in_aw_bits_id;
    line_241_valid_reg <= 4'hc == auto_in_aw_bits_id;
    line_242_valid_reg <= 4'hd == auto_in_aw_bits_id;
    line_243_valid_reg <= 4'he == auto_in_aw_bits_id;
    line_244_valid_reg <= 4'hf == auto_in_aw_bits_id;
    line_245_valid_reg <= 4'h0 == auto_in_aw_bits_id;
    line_246_valid_reg <= 4'h1 == auto_in_aw_bits_id;
    line_247_valid_reg <= 4'h2 == auto_in_aw_bits_id;
    line_248_valid_reg <= 4'h3 == auto_in_aw_bits_id;
    line_249_valid_reg <= 4'h4 == auto_in_aw_bits_id;
    line_250_valid_reg <= 4'h5 == auto_in_aw_bits_id;
    line_251_valid_reg <= 4'h6 == auto_in_aw_bits_id;
    line_252_valid_reg <= 4'h7 == auto_in_aw_bits_id;
    line_253_valid_reg <= 4'h8 == auto_in_aw_bits_id;
    line_254_valid_reg <= 4'h9 == auto_in_aw_bits_id;
    line_255_valid_reg <= 4'ha == auto_in_aw_bits_id;
    line_256_valid_reg <= 4'hb == auto_in_aw_bits_id;
    line_257_valid_reg <= 4'hc == auto_in_aw_bits_id;
    line_258_valid_reg <= 4'hd == auto_in_aw_bits_id;
    line_259_valid_reg <= 4'he == auto_in_aw_bits_id;
    line_260_valid_reg <= 4'hf == auto_in_aw_bits_id;
    line_261_valid_reg <= 4'h0 == auto_out_b_bits_id;
    line_262_valid_reg <= 4'h1 == auto_out_b_bits_id;
    line_263_valid_reg <= 4'h2 == auto_out_b_bits_id;
    line_264_valid_reg <= 4'h3 == auto_out_b_bits_id;
    line_265_valid_reg <= 4'h4 == auto_out_b_bits_id;
    line_266_valid_reg <= 4'h5 == auto_out_b_bits_id;
    line_267_valid_reg <= 4'h6 == auto_out_b_bits_id;
    line_268_valid_reg <= 4'h7 == auto_out_b_bits_id;
    line_269_valid_reg <= 4'h8 == auto_out_b_bits_id;
    line_270_valid_reg <= 4'h9 == auto_out_b_bits_id;
    line_271_valid_reg <= 4'ha == auto_out_b_bits_id;
    line_272_valid_reg <= 4'hb == auto_out_b_bits_id;
    line_273_valid_reg <= 4'hc == auto_out_b_bits_id;
    line_274_valid_reg <= 4'hd == auto_out_b_bits_id;
    line_275_valid_reg <= 4'he == auto_out_b_bits_id;
    line_276_valid_reg <= 4'hf == auto_out_b_bits_id;
    line_277_valid_reg <= _T_3;
    line_278_valid_reg <= _T_89;
    line_279_valid_reg <= 4'h0 == auto_out_b_bits_id;
    line_280_valid_reg <= 4'h1 == auto_out_b_bits_id;
    line_281_valid_reg <= 4'h2 == auto_out_b_bits_id;
    line_282_valid_reg <= 4'h3 == auto_out_b_bits_id;
    line_283_valid_reg <= 4'h4 == auto_out_b_bits_id;
    line_284_valid_reg <= 4'h5 == auto_out_b_bits_id;
    line_285_valid_reg <= 4'h6 == auto_out_b_bits_id;
    line_286_valid_reg <= 4'h7 == auto_out_b_bits_id;
    line_287_valid_reg <= 4'h8 == auto_out_b_bits_id;
    line_288_valid_reg <= 4'h9 == auto_out_b_bits_id;
    line_289_valid_reg <= 4'ha == auto_out_b_bits_id;
    line_290_valid_reg <= 4'hb == auto_out_b_bits_id;
    line_291_valid_reg <= 4'hc == auto_out_b_bits_id;
    line_292_valid_reg <= 4'hd == auto_out_b_bits_id;
    line_293_valid_reg <= 4'he == auto_out_b_bits_id;
    line_294_valid_reg <= 4'hf == auto_out_b_bits_id;
    line_295_valid_reg <= 4'h0 == auto_out_b_bits_id;
    line_296_valid_reg <= 4'h1 == auto_out_b_bits_id;
    line_297_valid_reg <= 4'h2 == auto_out_b_bits_id;
    line_298_valid_reg <= 4'h3 == auto_out_b_bits_id;
    line_299_valid_reg <= 4'h4 == auto_out_b_bits_id;
    line_300_valid_reg <= 4'h5 == auto_out_b_bits_id;
    line_301_valid_reg <= 4'h6 == auto_out_b_bits_id;
    line_302_valid_reg <= 4'h7 == auto_out_b_bits_id;
    line_303_valid_reg <= 4'h8 == auto_out_b_bits_id;
    line_304_valid_reg <= 4'h9 == auto_out_b_bits_id;
    line_305_valid_reg <= 4'ha == auto_out_b_bits_id;
    line_306_valid_reg <= 4'hb == auto_out_b_bits_id;
    line_307_valid_reg <= 4'hc == auto_out_b_bits_id;
    line_308_valid_reg <= 4'hd == auto_out_b_bits_id;
    line_309_valid_reg <= 4'he == auto_out_b_bits_id;
    line_310_valid_reg <= 4'hf == auto_out_b_bits_id;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_r_valid | _GEN_195)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n"
            ); // @[src/main/scala/amba/axi4/UserYanker.scala 66:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~auto_out_b_valid | _GEN_259)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UserYanker.scala:95 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n"
            ); // @[src/main/scala/amba/axi4/UserYanker.scala 95:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_147_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_148_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_149_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_150_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_151_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_152_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_153_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_154_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_155_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_156_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_157_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_158_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_159_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_160_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_161_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_162_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_163_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_164_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_165_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_166_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_167_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_168_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_169_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_170_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_171_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_172_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_173_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_174_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_175_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_176_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_177_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_178_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_179_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_180_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_181_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_182_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_183_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_184_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_185_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_186_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_187_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_188_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_189_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_190_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_191_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_192_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_193_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_194_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_195_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_196_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_197_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_198_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_199_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_200_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_201_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_202_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_203_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_204_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_205_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_206_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_207_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_208_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_209_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_210_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_211_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_212_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_213_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_214_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_215_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_216_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_217_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_218_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_219_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_220_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_221_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_222_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_223_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_224_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_225_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_226_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_227_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_228_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_229_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_230_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_231_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_232_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_233_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_234_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_235_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_236_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_237_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_238_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_239_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_240_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_241_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_242_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_243_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_244_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_245_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_246_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_247_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_248_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_249_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_250_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_251_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_252_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_253_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_254_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_255_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_256_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_257_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_258_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_259_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_260_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_261_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_262_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_263_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_264_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_265_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_266_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_267_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_268_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_269_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_270_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_271_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_272_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_273_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_274_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_275_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_276_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_277_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_278_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_279_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_280_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_281_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_282_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_283_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_284_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_285_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_286_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_287_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_288_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_289_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_290_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_291_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_292_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_293_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_294_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_295_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_296_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_297_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_298_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_299_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_300_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_301_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_302_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_303_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_304_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_305_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_306_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_307_valid_reg = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  line_308_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  line_309_valid_reg = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  line_310_valid_reg = _RAND_163[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~auto_out_r_valid | _GEN_195); // @[src/main/scala/amba/axi4/UserYanker.scala 66:14]
    end
    //
    if (_T_3) begin
      assert(~auto_out_b_valid | _GEN_259); // @[src/main/scala/amba/axi4/UserYanker.scala 95:14]
    end
  end
endmodule
module AXI4IdIndexer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_echo_tl_state_size = auto_out_b_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_echo_tl_state_source = auto_out_b_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_echo_tl_state_size = auto_out_r_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_echo_tl_state_source = auto_out_r_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_echo_tl_state_size = auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_echo_tl_state_source = auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_echo_tl_state_size = auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_echo_tl_state_source = auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module Queue_34(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_strb [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_last [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_17 = io_deq_ready ? 1'h0 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 324:26 286:27 324:35]
  wire  do_enq = empty ? _GEN_17 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 286:27]
  wire  line_311_clock;
  wire  line_311_reset;
  wire  line_311_valid;
  reg  line_311_valid_reg;
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 323:14 287:27]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_312_clock;
  wire  line_312_reset;
  wire  line_312_valid;
  reg  line_312_valid_reg;
  wire  line_313_clock;
  wire  line_313_reset;
  wire  line_313_valid;
  reg  line_313_valid_reg;
  wire  line_314_clock;
  wire  line_314_reset;
  wire  line_314_valid;
  reg  line_314_valid_reg;
  wire  line_315_clock;
  wire  line_315_reset;
  wire  line_315_valid;
  reg  line_315_valid_reg;
  GEN_w1_line #(.COVER_INDEX(311)) line_311 (
    .clock(line_311_clock),
    .reset(line_311_reset),
    .valid(line_311_valid)
  );
  GEN_w1_line #(.COVER_INDEX(312)) line_312 (
    .clock(line_312_clock),
    .reset(line_312_reset),
    .valid(line_312_valid)
  );
  GEN_w1_line #(.COVER_INDEX(313)) line_313 (
    .clock(line_313_clock),
    .reset(line_313_reset),
    .valid(line_313_valid)
  );
  GEN_w1_line #(.COVER_INDEX(314)) line_314 (
    .clock(line_314_clock),
    .reset(line_314_reset),
    .valid(line_314_valid)
  );
  GEN_w1_line #(.COVER_INDEX(315)) line_315 (
    .clock(line_315_clock),
    .reset(line_315_reset),
    .valid(line_315_valid)
  );
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = 1'h0;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign line_311_clock = clock;
  assign line_311_reset = reset;
  assign line_311_valid = do_enq ^ line_311_valid_reg;
  assign line_312_clock = clock;
  assign line_312_reset = reset;
  assign line_312_valid = _T ^ line_312_valid_reg;
  assign line_313_clock = clock;
  assign line_313_reset = reset;
  assign line_313_valid = io_enq_valid ^ line_313_valid_reg;
  assign line_314_clock = clock;
  assign line_314_reset = reset;
  assign line_314_valid = empty ^ line_314_valid_reg;
  assign line_315_clock = clock;
  assign line_315_reset = reset;
  assign line_315_valid = io_deq_ready ^ line_315_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:16 320:{24,39}]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_strb = empty ? io_enq_bits_strb : ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
        if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
          maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
        end else begin
          maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end
    if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
      if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
        line_311_valid_reg <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
      end else begin
        line_311_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end else begin
      line_311_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
    end
    line_312_valid_reg <= _T;
    line_313_valid_reg <= io_enq_valid;
    line_314_valid_reg <= empty;
    line_315_valid_reg <= io_deq_ready;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_311_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_312_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_313_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_314_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_315_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_35(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_echo_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_echo_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_wen, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_burst, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_echo_tl_state_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_echo_tl_state_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_wen // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_addr [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_len [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_burst [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_echo_tl_state_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_echo_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [3:0] ram_echo_tl_state_source [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_echo_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_tl_state_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_wen [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_wen_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_26 = io_deq_ready ? 1'h0 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 324:26 286:27 324:35]
  wire  do_enq = empty ? _GEN_26 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 286:27]
  wire  line_316_clock;
  wire  line_316_reset;
  wire  line_316_valid;
  reg  line_316_valid_reg;
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 323:14 287:27]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_317_clock;
  wire  line_317_reset;
  wire  line_317_valid;
  reg  line_317_valid_reg;
  wire  line_318_clock;
  wire  line_318_reset;
  wire  line_318_valid;
  reg  line_318_valid_reg;
  wire  line_319_clock;
  wire  line_319_reset;
  wire  line_319_valid;
  reg  line_319_valid_reg;
  wire  line_320_clock;
  wire  line_320_reset;
  wire  line_320_valid;
  reg  line_320_valid_reg;
  GEN_w1_line #(.COVER_INDEX(316)) line_316 (
    .clock(line_316_clock),
    .reset(line_316_reset),
    .valid(line_316_valid)
  );
  GEN_w1_line #(.COVER_INDEX(317)) line_317 (
    .clock(line_317_clock),
    .reset(line_317_reset),
    .valid(line_317_valid)
  );
  GEN_w1_line #(.COVER_INDEX(318)) line_318 (
    .clock(line_318_clock),
    .reset(line_318_reset),
    .valid(line_318_valid)
  );
  GEN_w1_line #(.COVER_INDEX(319)) line_319 (
    .clock(line_319_clock),
    .reset(line_319_reset),
    .valid(line_319_valid)
  );
  GEN_w1_line #(.COVER_INDEX(320)) line_320 (
    .clock(line_320_clock),
    .reset(line_320_reset),
    .valid(line_320_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_burst_MPORT_data = 2'h1;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_io_deq_bits_MPORT_data =
    ram_echo_tl_state_size[ram_echo_tl_state_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_tl_state_size_MPORT_data = io_enq_bits_echo_tl_state_size;
  assign ram_echo_tl_state_size_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_size_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_size_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_io_deq_bits_MPORT_data =
    ram_echo_tl_state_source[ram_echo_tl_state_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_tl_state_source_MPORT_data = io_enq_bits_echo_tl_state_source;
  assign ram_echo_tl_state_source_MPORT_addr = 1'h0;
  assign ram_echo_tl_state_source_MPORT_mask = 1'h1;
  assign ram_echo_tl_state_source_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign ram_wen_io_deq_bits_MPORT_en = 1'h1;
  assign ram_wen_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_wen_io_deq_bits_MPORT_data = ram_wen[ram_wen_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_wen_MPORT_data = io_enq_bits_wen;
  assign ram_wen_MPORT_addr = 1'h0;
  assign ram_wen_MPORT_mask = 1'h1;
  assign ram_wen_MPORT_en = empty ? _GEN_26 : _do_enq_T;
  assign line_316_clock = clock;
  assign line_316_reset = reset;
  assign line_316_valid = do_enq ^ line_316_valid_reg;
  assign line_317_clock = clock;
  assign line_317_reset = reset;
  assign line_317_valid = _T ^ line_317_valid_reg;
  assign line_318_clock = clock;
  assign line_318_reset = reset;
  assign line_318_valid = io_enq_valid ^ line_318_valid_reg;
  assign line_319_clock = clock;
  assign line_319_reset = reset;
  assign line_319_valid = empty ^ line_319_valid_reg;
  assign line_320_clock = clock;
  assign line_320_reset = reset;
  assign line_320_valid = io_deq_ready ^ line_320_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:16 320:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_burst = empty ? 2'h1 : ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_echo_tl_state_size = empty ? io_enq_bits_echo_tl_state_size :
    ram_echo_tl_state_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_echo_tl_state_source = empty ? io_enq_bits_echo_tl_state_source :
    ram_echo_tl_state_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_wen = empty ? io_enq_bits_wen : ram_wen_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_tl_state_size_MPORT_en & ram_echo_tl_state_size_MPORT_mask) begin
      ram_echo_tl_state_size[ram_echo_tl_state_size_MPORT_addr] <= ram_echo_tl_state_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_tl_state_source_MPORT_en & ram_echo_tl_state_source_MPORT_mask) begin
      ram_echo_tl_state_source[ram_echo_tl_state_source_MPORT_addr] <= ram_echo_tl_state_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_wen_MPORT_en & ram_wen_MPORT_mask) begin
      ram_wen[ram_wen_MPORT_addr] <= ram_wen_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
        if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
          maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
        end else begin
          maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end
    if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
      if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
        line_316_valid_reg <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
      end else begin
        line_316_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end else begin
      line_316_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
    end
    line_317_valid_reg <= _T;
    line_318_valid_reg <= io_enq_valid;
    line_319_valid_reg <= empty;
    line_320_valid_reg <= io_deq_ready;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_size[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_echo_tl_state_source[initvar] = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_316_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_317_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_318_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_319_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_320_valid_reg = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLToAXI4(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_echo_tl_state_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_echo_tl_state_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
`endif // RANDOMIZE_REG_INIT
  wire  nodeOut_w_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_w_deq_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_w_deq_q_io_enq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_enq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] queue_arw_deq_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] queue_arw_deq_q_io_enq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] queue_arw_deq_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_enq_bits_echo_tl_state_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_enq_bits_echo_tl_state_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_enq_bits_wen; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] queue_arw_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] queue_arw_deq_q_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] queue_arw_deq_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] queue_arw_deq_q_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_deq_bits_echo_tl_state_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] queue_arw_deq_q_io_deq_bits_echo_tl_state_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  queue_arw_deq_q_io_deq_bits_wen; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  a_isPut = ~auto_in_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  reg  count_16; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_15 = ~count_16; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_15; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_14 = ~count_15; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_14; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_13 = ~count_14; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_13; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_12 = ~count_13; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_12; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_11 = ~count_12; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_11; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_10 = ~count_11; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_10; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_9 = ~count_10; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_9; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_8 = ~count_9; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_8; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_7 = ~count_8; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_7; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_6 = ~count_7; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_6; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_5 = ~count_6; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_5; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_4 = ~count_5; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_4; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_3 = ~count_4; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_3; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_2 = ~count_3; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_2; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle_1 = ~count_2; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  reg  count_1; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
  wire  idle = ~count_1; // @[src/main/scala/tilelink/ToAXI4.scala 267:26]
  wire  _GEN_138 = 4'h1 == auto_in_a_bits_source ? count_2 : count_1; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_139 = 4'h2 == auto_in_a_bits_source ? count_3 : _GEN_138; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_140 = 4'h3 == auto_in_a_bits_source ? count_4 : _GEN_139; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_141 = 4'h4 == auto_in_a_bits_source ? count_5 : _GEN_140; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_142 = 4'h5 == auto_in_a_bits_source ? count_6 : _GEN_141; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_143 = 4'h6 == auto_in_a_bits_source ? count_7 : _GEN_142; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_144 = 4'h7 == auto_in_a_bits_source ? count_8 : _GEN_143; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_145 = 4'h8 == auto_in_a_bits_source ? count_9 : _GEN_144; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_146 = 4'h9 == auto_in_a_bits_source ? count_10 : _GEN_145; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_147 = 4'ha == auto_in_a_bits_source ? count_11 : _GEN_146; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_148 = 4'hb == auto_in_a_bits_source ? count_12 : _GEN_147; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_149 = 4'hc == auto_in_a_bits_source ? count_13 : _GEN_148; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_150 = 4'hd == auto_in_a_bits_source ? count_14 : _GEN_149; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_151 = 4'he == auto_in_a_bits_source ? count_15 : _GEN_150; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  wire  _GEN_152 = 4'hf == auto_in_a_bits_source ? count_16 : _GEN_151; // @[src/main/scala/tilelink/ToAXI4.scala 198:{49,49}]
  reg [1:0] counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire  a_first = counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  stall = _GEN_152 & a_first; // @[src/main/scala/tilelink/ToAXI4.scala 198:49]
  wire  _nodeIn_a_ready_T = ~stall; // @[src/main/scala/tilelink/ToAXI4.scala 199:21]
  reg  doneAW; // @[src/main/scala/tilelink/ToAXI4.scala 160:30]
  wire  out_arw_ready = queue_arw_deq_q_io_enq_ready; // @[src/main/scala/tilelink/ToAXI4.scala 146:25 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  wire  _nodeIn_a_ready_T_1 = doneAW | out_arw_ready; // @[src/main/scala/tilelink/ToAXI4.scala 199:52]
  wire  out_w_ready = nodeOut_w_deq_q_io_enq_ready; // @[src/main/scala/tilelink/ToAXI4.scala 147:23 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  wire  _nodeIn_a_ready_T_3 = a_isPut ? (doneAW | out_arw_ready) & out_w_ready : out_arw_ready; // @[src/main/scala/tilelink/ToAXI4.scala 199:34]
  wire  nodeIn_a_ready = ~stall & _nodeIn_a_ready_T_3; // @[src/main/scala/tilelink/ToAXI4.scala 199:28]
  wire  _T = nodeIn_a_ready & auto_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _beats1_decode_T_1 = 12'h1f << auto_in_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beats1_decode = _beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire [1:0] beats1 = a_isPut ? beats1_decode : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire [1:0] counter1 = counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  a_last = counter == 2'h1 | beats1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  line_321_clock;
  wire  line_321_reset;
  wire  line_321_valid;
  reg  line_321_valid_reg;
  wire  queue_arw_bits_wen = queue_arw_deq_q_io_deq_bits_wen; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire  queue_arw_valid = queue_arw_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  wire  line_322_clock;
  wire  line_322_reset;
  wire  line_322_valid;
  reg  line_322_valid_reg;
  wire  line_323_clock;
  wire  line_323_reset;
  wire  line_323_valid;
  reg  line_323_valid_reg;
  wire  line_324_clock;
  wire  line_324_reset;
  wire  line_324_valid;
  reg  line_324_valid_reg;
  wire [3:0] _GEN_122 = 4'h1 == auto_in_a_bits_source ? 4'h1 : 4'h0; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_325_clock;
  wire  line_325_reset;
  wire  line_325_valid;
  reg  line_325_valid_reg;
  wire [3:0] _GEN_123 = 4'h2 == auto_in_a_bits_source ? 4'h2 : _GEN_122; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_326_clock;
  wire  line_326_reset;
  wire  line_326_valid;
  reg  line_326_valid_reg;
  wire [3:0] _GEN_124 = 4'h3 == auto_in_a_bits_source ? 4'h3 : _GEN_123; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_327_clock;
  wire  line_327_reset;
  wire  line_327_valid;
  reg  line_327_valid_reg;
  wire [3:0] _GEN_125 = 4'h4 == auto_in_a_bits_source ? 4'h4 : _GEN_124; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_328_clock;
  wire  line_328_reset;
  wire  line_328_valid;
  reg  line_328_valid_reg;
  wire [3:0] _GEN_126 = 4'h5 == auto_in_a_bits_source ? 4'h5 : _GEN_125; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_329_clock;
  wire  line_329_reset;
  wire  line_329_valid;
  reg  line_329_valid_reg;
  wire [3:0] _GEN_127 = 4'h6 == auto_in_a_bits_source ? 4'h6 : _GEN_126; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_330_clock;
  wire  line_330_reset;
  wire  line_330_valid;
  reg  line_330_valid_reg;
  wire [3:0] _GEN_128 = 4'h7 == auto_in_a_bits_source ? 4'h7 : _GEN_127; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_331_clock;
  wire  line_331_reset;
  wire  line_331_valid;
  reg  line_331_valid_reg;
  wire [3:0] _GEN_129 = 4'h8 == auto_in_a_bits_source ? 4'h8 : _GEN_128; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_332_clock;
  wire  line_332_reset;
  wire  line_332_valid;
  reg  line_332_valid_reg;
  wire [3:0] _GEN_130 = 4'h9 == auto_in_a_bits_source ? 4'h9 : _GEN_129; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_333_clock;
  wire  line_333_reset;
  wire  line_333_valid;
  reg  line_333_valid_reg;
  wire [3:0] _GEN_131 = 4'ha == auto_in_a_bits_source ? 4'ha : _GEN_130; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_334_clock;
  wire  line_334_reset;
  wire  line_334_valid;
  reg  line_334_valid_reg;
  wire [3:0] _GEN_132 = 4'hb == auto_in_a_bits_source ? 4'hb : _GEN_131; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_335_clock;
  wire  line_335_reset;
  wire  line_335_valid;
  reg  line_335_valid_reg;
  wire [3:0] _GEN_133 = 4'hc == auto_in_a_bits_source ? 4'hc : _GEN_132; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_336_clock;
  wire  line_336_reset;
  wire  line_336_valid;
  reg  line_336_valid_reg;
  wire [3:0] _GEN_134 = 4'hd == auto_in_a_bits_source ? 4'hd : _GEN_133; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_337_clock;
  wire  line_337_reset;
  wire  line_337_valid;
  reg  line_337_valid_reg;
  wire [3:0] _GEN_135 = 4'he == auto_in_a_bits_source ? 4'he : _GEN_134; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire  line_338_clock;
  wire  line_338_reset;
  wire  line_338_valid;
  reg  line_338_valid_reg;
  wire [3:0] out_arw_bits_id = 4'hf == auto_in_a_bits_source ? 4'hf : _GEN_135; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  wire [17:0] _out_arw_bits_len_T_1 = 18'h7ff << auto_in_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [10:0] _out_arw_bits_len_T_3 = ~_out_arw_bits_len_T_1[10:0]; // @[src/main/scala/util/package.scala 235:46]
  wire  line_339_clock;
  wire  line_339_reset;
  wire  line_339_valid;
  reg  line_339_valid_reg;
  wire  line_340_clock;
  wire  line_340_reset;
  wire  line_340_valid;
  reg  line_340_valid_reg;
  wire  line_341_clock;
  wire  line_341_reset;
  wire  line_341_valid;
  reg  line_341_valid_reg;
  wire  line_342_clock;
  wire  line_342_reset;
  wire  line_342_valid;
  reg  line_342_valid_reg;
  wire  line_343_clock;
  wire  line_343_reset;
  wire  line_343_valid;
  reg  line_343_valid_reg;
  wire  line_344_clock;
  wire  line_344_reset;
  wire  line_344_valid;
  reg  line_344_valid_reg;
  wire  line_345_clock;
  wire  line_345_reset;
  wire  line_345_valid;
  reg  line_345_valid_reg;
  wire  line_346_clock;
  wire  line_346_reset;
  wire  line_346_valid;
  reg  line_346_valid_reg;
  wire  line_347_clock;
  wire  line_347_reset;
  wire  line_347_valid;
  reg  line_347_valid_reg;
  wire  line_348_clock;
  wire  line_348_reset;
  wire  line_348_valid;
  reg  line_348_valid_reg;
  wire  line_349_clock;
  wire  line_349_reset;
  wire  line_349_valid;
  reg  line_349_valid_reg;
  wire  line_350_clock;
  wire  line_350_reset;
  wire  line_350_valid;
  reg  line_350_valid_reg;
  wire  line_351_clock;
  wire  line_351_reset;
  wire  line_351_valid;
  reg  line_351_valid_reg;
  wire  line_352_clock;
  wire  line_352_reset;
  wire  line_352_valid;
  reg  line_352_valid_reg;
  wire  line_353_clock;
  wire  line_353_reset;
  wire  line_353_valid;
  reg  line_353_valid_reg;
  wire  line_354_clock;
  wire  line_354_reset;
  wire  line_354_valid;
  reg  line_354_valid_reg;
  wire  _out_arw_valid_T_1 = _nodeIn_a_ready_T & auto_in_a_valid; // @[src/main/scala/tilelink/ToAXI4.scala 200:31]
  wire  _out_arw_valid_T_4 = a_isPut ? ~doneAW & out_w_ready : 1'h1; // @[src/main/scala/tilelink/ToAXI4.scala 200:51]
  wire  out_arw_valid = _nodeIn_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[src/main/scala/tilelink/ToAXI4.scala 200:45]
  reg  r_holds_d; // @[src/main/scala/tilelink/ToAXI4.scala 209:30]
  reg [2:0] b_delay; // @[src/main/scala/tilelink/ToAXI4.scala 212:24]
  wire  r_wins = auto_out_r_valid & b_delay != 3'h7 | r_holds_d; // @[src/main/scala/tilelink/ToAXI4.scala 218:53]
  wire  nodeOut_r_ready = auto_in_d_ready & r_wins; // @[src/main/scala/tilelink/ToAXI4.scala 220:33]
  wire  _T_2 = nodeOut_r_ready & auto_out_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_355_clock;
  wire  line_355_reset;
  wire  line_355_valid;
  reg  line_355_valid_reg;
  wire  nodeOut_b_ready = auto_in_d_ready & ~r_wins; // @[src/main/scala/tilelink/ToAXI4.scala 221:33]
  wire  _T_4 = auto_out_b_valid & ~nodeOut_b_ready; // @[src/main/scala/tilelink/ToAXI4.scala 213:25]
  wire  line_356_clock;
  wire  line_356_reset;
  wire  line_356_valid;
  reg  line_356_valid_reg;
  wire [2:0] _b_delay_T_1 = b_delay + 3'h1; // @[src/main/scala/tilelink/ToAXI4.scala 214:28]
  wire  line_357_clock;
  wire  line_357_reset;
  wire  line_357_valid;
  reg  line_357_valid_reg;
  wire  nodeIn_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[src/main/scala/tilelink/ToAXI4.scala 222:24]
  reg  r_first; // @[src/main/scala/tilelink/ToAXI4.scala 227:28]
  wire  line_358_clock;
  wire  line_358_reset;
  wire  line_358_valid;
  reg  line_358_valid_reg;
  wire  _GEN_155 = _T_2 ? auto_out_r_bits_last : r_first; // @[src/main/scala/tilelink/ToAXI4.scala 228:25 227:28 228:35]
  wire  _r_denied_T = auto_out_r_bits_resp == 2'h3; // @[src/main/scala/tilelink/ToAXI4.scala 229:39]
  reg  r_denied_r; // @[src/main/scala/util/package.scala 80:63]
  wire  line_359_clock;
  wire  line_359_reset;
  wire  line_359_valid;
  reg  line_359_valid_reg;
  wire  _GEN_156 = r_first ? _r_denied_T : r_denied_r; // @[src/main/scala/util/package.scala 80:{63,63,63}]
  wire  r_corrupt = auto_out_r_bits_resp != 2'h0; // @[src/main/scala/tilelink/ToAXI4.scala 230:39]
  wire  b_denied = auto_out_b_bits_resp != 2'h0; // @[src/main/scala/tilelink/ToAXI4.scala 231:39]
  wire  r_d_corrupt = r_corrupt | _GEN_156; // @[src/main/scala/tilelink/ToAXI4.scala 233:96]
  wire [2:0] r_d_size = auto_out_r_bits_echo_tl_state_size[2:0]; // @[src/main/scala/tilelink/Edges.scala 810:17 813:15]
  wire [2:0] b_d_size = auto_out_b_bits_echo_tl_state_size[2:0]; // @[src/main/scala/tilelink/Edges.scala 792:17 795:15]
  wire [15:0] _a_sel_T = 16'h1 << out_arw_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  a_sel_0 = _a_sel_T[0]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_1 = _a_sel_T[1]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_2 = _a_sel_T[2]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_3 = _a_sel_T[3]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_4 = _a_sel_T[4]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_5 = _a_sel_T[5]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_6 = _a_sel_T[6]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_7 = _a_sel_T[7]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_8 = _a_sel_T[8]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_9 = _a_sel_T[9]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_10 = _a_sel_T[10]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_11 = _a_sel_T[11]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_12 = _a_sel_T[12]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_13 = _a_sel_T[13]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_14 = _a_sel_T[14]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire  a_sel_15 = _a_sel_T[15]; // @[src/main/scala/tilelink/ToAXI4.scala 253:58]
  wire [3:0] d_sel_shiftAmount = r_wins ? auto_out_r_bits_id : auto_out_b_bits_id; // @[src/main/scala/tilelink/ToAXI4.scala 254:31]
  wire [15:0] _d_sel_T_1 = 16'h1 << d_sel_shiftAmount; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  d_sel_0 = _d_sel_T_1[0]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_1 = _d_sel_T_1[1]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_2 = _d_sel_T_1[2]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_3 = _d_sel_T_1[3]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_4 = _d_sel_T_1[4]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_5 = _d_sel_T_1[5]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_6 = _d_sel_T_1[6]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_7 = _d_sel_T_1[7]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_8 = _d_sel_T_1[8]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_9 = _d_sel_T_1[9]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_10 = _d_sel_T_1[10]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_11 = _d_sel_T_1[11]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_12 = _d_sel_T_1[12]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_13 = _d_sel_T_1[13]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_14 = _d_sel_T_1[14]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_sel_15 = _d_sel_T_1[15]; // @[src/main/scala/tilelink/ToAXI4.scala 254:93]
  wire  d_last = r_wins ? auto_out_r_bits_last : 1'h1; // @[src/main/scala/tilelink/ToAXI4.scala 255:23]
  wire  _inc_T = out_arw_ready & out_arw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  inc = a_sel_0 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  _dec_T_1 = auto_in_d_ready & nodeIn_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  dec = d_sel_0 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_2 = count_1 + inc; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  _T_10 = ~reset; // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_360_clock;
  wire  line_360_reset;
  wire  line_360_valid;
  reg  line_360_valid_reg;
  wire  _T_11 = ~(~dec | count_1); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_361_clock;
  wire  line_361_reset;
  wire  line_361_valid;
  reg  line_361_valid_reg;
  wire  line_362_clock;
  wire  line_362_reset;
  wire  line_362_valid;
  reg  line_362_valid_reg;
  wire  _T_17 = ~(~inc | idle); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_363_clock;
  wire  line_363_reset;
  wire  line_363_valid;
  reg  line_363_valid_reg;
  wire  line_364_clock;
  wire  line_364_reset;
  wire  line_364_valid;
  reg  line_364_valid_reg;
  wire  inc_1 = a_sel_1 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_1 = d_sel_1 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_6 = count_2 + inc_1; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_365_clock;
  wire  line_365_reset;
  wire  line_365_valid;
  reg  line_365_valid_reg;
  wire  _T_23 = ~(~dec_1 | count_2); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_366_clock;
  wire  line_366_reset;
  wire  line_366_valid;
  reg  line_366_valid_reg;
  wire  line_367_clock;
  wire  line_367_reset;
  wire  line_367_valid;
  reg  line_367_valid_reg;
  wire  _T_29 = ~(~inc_1 | idle_1); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_368_clock;
  wire  line_368_reset;
  wire  line_368_valid;
  reg  line_368_valid_reg;
  wire  line_369_clock;
  wire  line_369_reset;
  wire  line_369_valid;
  reg  line_369_valid_reg;
  wire  inc_2 = a_sel_2 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_2 = d_sel_2 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_10 = count_3 + inc_2; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_370_clock;
  wire  line_370_reset;
  wire  line_370_valid;
  reg  line_370_valid_reg;
  wire  _T_35 = ~(~dec_2 | count_3); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_371_clock;
  wire  line_371_reset;
  wire  line_371_valid;
  reg  line_371_valid_reg;
  wire  line_372_clock;
  wire  line_372_reset;
  wire  line_372_valid;
  reg  line_372_valid_reg;
  wire  _T_41 = ~(~inc_2 | idle_2); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_373_clock;
  wire  line_373_reset;
  wire  line_373_valid;
  reg  line_373_valid_reg;
  wire  line_374_clock;
  wire  line_374_reset;
  wire  line_374_valid;
  reg  line_374_valid_reg;
  wire  inc_3 = a_sel_3 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_3 = d_sel_3 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_14 = count_4 + inc_3; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_375_clock;
  wire  line_375_reset;
  wire  line_375_valid;
  reg  line_375_valid_reg;
  wire  _T_47 = ~(~dec_3 | count_4); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_376_clock;
  wire  line_376_reset;
  wire  line_376_valid;
  reg  line_376_valid_reg;
  wire  line_377_clock;
  wire  line_377_reset;
  wire  line_377_valid;
  reg  line_377_valid_reg;
  wire  _T_53 = ~(~inc_3 | idle_3); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_378_clock;
  wire  line_378_reset;
  wire  line_378_valid;
  reg  line_378_valid_reg;
  wire  line_379_clock;
  wire  line_379_reset;
  wire  line_379_valid;
  reg  line_379_valid_reg;
  wire  inc_4 = a_sel_4 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_4 = d_sel_4 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_18 = count_5 + inc_4; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_380_clock;
  wire  line_380_reset;
  wire  line_380_valid;
  reg  line_380_valid_reg;
  wire  _T_59 = ~(~dec_4 | count_5); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_381_clock;
  wire  line_381_reset;
  wire  line_381_valid;
  reg  line_381_valid_reg;
  wire  line_382_clock;
  wire  line_382_reset;
  wire  line_382_valid;
  reg  line_382_valid_reg;
  wire  _T_65 = ~(~inc_4 | idle_4); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_383_clock;
  wire  line_383_reset;
  wire  line_383_valid;
  reg  line_383_valid_reg;
  wire  line_384_clock;
  wire  line_384_reset;
  wire  line_384_valid;
  reg  line_384_valid_reg;
  wire  inc_5 = a_sel_5 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_5 = d_sel_5 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_22 = count_6 + inc_5; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_385_clock;
  wire  line_385_reset;
  wire  line_385_valid;
  reg  line_385_valid_reg;
  wire  _T_71 = ~(~dec_5 | count_6); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_386_clock;
  wire  line_386_reset;
  wire  line_386_valid;
  reg  line_386_valid_reg;
  wire  line_387_clock;
  wire  line_387_reset;
  wire  line_387_valid;
  reg  line_387_valid_reg;
  wire  _T_77 = ~(~inc_5 | idle_5); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_388_clock;
  wire  line_388_reset;
  wire  line_388_valid;
  reg  line_388_valid_reg;
  wire  line_389_clock;
  wire  line_389_reset;
  wire  line_389_valid;
  reg  line_389_valid_reg;
  wire  inc_6 = a_sel_6 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_6 = d_sel_6 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_26 = count_7 + inc_6; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_390_clock;
  wire  line_390_reset;
  wire  line_390_valid;
  reg  line_390_valid_reg;
  wire  _T_83 = ~(~dec_6 | count_7); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_391_clock;
  wire  line_391_reset;
  wire  line_391_valid;
  reg  line_391_valid_reg;
  wire  line_392_clock;
  wire  line_392_reset;
  wire  line_392_valid;
  reg  line_392_valid_reg;
  wire  _T_89 = ~(~inc_6 | idle_6); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_393_clock;
  wire  line_393_reset;
  wire  line_393_valid;
  reg  line_393_valid_reg;
  wire  line_394_clock;
  wire  line_394_reset;
  wire  line_394_valid;
  reg  line_394_valid_reg;
  wire  inc_7 = a_sel_7 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_7 = d_sel_7 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_30 = count_8 + inc_7; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_395_clock;
  wire  line_395_reset;
  wire  line_395_valid;
  reg  line_395_valid_reg;
  wire  _T_95 = ~(~dec_7 | count_8); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_396_clock;
  wire  line_396_reset;
  wire  line_396_valid;
  reg  line_396_valid_reg;
  wire  line_397_clock;
  wire  line_397_reset;
  wire  line_397_valid;
  reg  line_397_valid_reg;
  wire  _T_101 = ~(~inc_7 | idle_7); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_398_clock;
  wire  line_398_reset;
  wire  line_398_valid;
  reg  line_398_valid_reg;
  wire  line_399_clock;
  wire  line_399_reset;
  wire  line_399_valid;
  reg  line_399_valid_reg;
  wire  inc_8 = a_sel_8 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_8 = d_sel_8 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_34 = count_9 + inc_8; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_400_clock;
  wire  line_400_reset;
  wire  line_400_valid;
  reg  line_400_valid_reg;
  wire  _T_107 = ~(~dec_8 | count_9); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_401_clock;
  wire  line_401_reset;
  wire  line_401_valid;
  reg  line_401_valid_reg;
  wire  line_402_clock;
  wire  line_402_reset;
  wire  line_402_valid;
  reg  line_402_valid_reg;
  wire  _T_113 = ~(~inc_8 | idle_8); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_403_clock;
  wire  line_403_reset;
  wire  line_403_valid;
  reg  line_403_valid_reg;
  wire  line_404_clock;
  wire  line_404_reset;
  wire  line_404_valid;
  reg  line_404_valid_reg;
  wire  inc_9 = a_sel_9 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_9 = d_sel_9 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_38 = count_10 + inc_9; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_405_clock;
  wire  line_405_reset;
  wire  line_405_valid;
  reg  line_405_valid_reg;
  wire  _T_119 = ~(~dec_9 | count_10); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_406_clock;
  wire  line_406_reset;
  wire  line_406_valid;
  reg  line_406_valid_reg;
  wire  line_407_clock;
  wire  line_407_reset;
  wire  line_407_valid;
  reg  line_407_valid_reg;
  wire  _T_125 = ~(~inc_9 | idle_9); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_408_clock;
  wire  line_408_reset;
  wire  line_408_valid;
  reg  line_408_valid_reg;
  wire  line_409_clock;
  wire  line_409_reset;
  wire  line_409_valid;
  reg  line_409_valid_reg;
  wire  inc_10 = a_sel_10 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_10 = d_sel_10 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_42 = count_11 + inc_10; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_410_clock;
  wire  line_410_reset;
  wire  line_410_valid;
  reg  line_410_valid_reg;
  wire  _T_131 = ~(~dec_10 | count_11); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_411_clock;
  wire  line_411_reset;
  wire  line_411_valid;
  reg  line_411_valid_reg;
  wire  line_412_clock;
  wire  line_412_reset;
  wire  line_412_valid;
  reg  line_412_valid_reg;
  wire  _T_137 = ~(~inc_10 | idle_10); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_413_clock;
  wire  line_413_reset;
  wire  line_413_valid;
  reg  line_413_valid_reg;
  wire  line_414_clock;
  wire  line_414_reset;
  wire  line_414_valid;
  reg  line_414_valid_reg;
  wire  inc_11 = a_sel_11 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_11 = d_sel_11 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_46 = count_12 + inc_11; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_415_clock;
  wire  line_415_reset;
  wire  line_415_valid;
  reg  line_415_valid_reg;
  wire  _T_143 = ~(~dec_11 | count_12); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_416_clock;
  wire  line_416_reset;
  wire  line_416_valid;
  reg  line_416_valid_reg;
  wire  line_417_clock;
  wire  line_417_reset;
  wire  line_417_valid;
  reg  line_417_valid_reg;
  wire  _T_149 = ~(~inc_11 | idle_11); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_418_clock;
  wire  line_418_reset;
  wire  line_418_valid;
  reg  line_418_valid_reg;
  wire  line_419_clock;
  wire  line_419_reset;
  wire  line_419_valid;
  reg  line_419_valid_reg;
  wire  inc_12 = a_sel_12 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_12 = d_sel_12 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_50 = count_13 + inc_12; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_420_clock;
  wire  line_420_reset;
  wire  line_420_valid;
  reg  line_420_valid_reg;
  wire  _T_155 = ~(~dec_12 | count_13); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_421_clock;
  wire  line_421_reset;
  wire  line_421_valid;
  reg  line_421_valid_reg;
  wire  line_422_clock;
  wire  line_422_reset;
  wire  line_422_valid;
  reg  line_422_valid_reg;
  wire  _T_161 = ~(~inc_12 | idle_12); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_423_clock;
  wire  line_423_reset;
  wire  line_423_valid;
  reg  line_423_valid_reg;
  wire  line_424_clock;
  wire  line_424_reset;
  wire  line_424_valid;
  reg  line_424_valid_reg;
  wire  inc_13 = a_sel_13 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_13 = d_sel_13 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_54 = count_14 + inc_13; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_425_clock;
  wire  line_425_reset;
  wire  line_425_valid;
  reg  line_425_valid_reg;
  wire  _T_167 = ~(~dec_13 | count_14); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_426_clock;
  wire  line_426_reset;
  wire  line_426_valid;
  reg  line_426_valid_reg;
  wire  line_427_clock;
  wire  line_427_reset;
  wire  line_427_valid;
  reg  line_427_valid_reg;
  wire  _T_173 = ~(~inc_13 | idle_13); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_428_clock;
  wire  line_428_reset;
  wire  line_428_valid;
  reg  line_428_valid_reg;
  wire  line_429_clock;
  wire  line_429_reset;
  wire  line_429_valid;
  reg  line_429_valid_reg;
  wire  inc_14 = a_sel_14 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_14 = d_sel_14 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_58 = count_15 + inc_14; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_430_clock;
  wire  line_430_reset;
  wire  line_430_valid;
  reg  line_430_valid_reg;
  wire  _T_179 = ~(~dec_14 | count_15); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_431_clock;
  wire  line_431_reset;
  wire  line_431_valid;
  reg  line_431_valid_reg;
  wire  line_432_clock;
  wire  line_432_reset;
  wire  line_432_valid;
  reg  line_432_valid_reg;
  wire  _T_185 = ~(~inc_14 | idle_14); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_433_clock;
  wire  line_433_reset;
  wire  line_433_valid;
  reg  line_433_valid_reg;
  wire  line_434_clock;
  wire  line_434_reset;
  wire  line_434_valid;
  reg  line_434_valid_reg;
  wire  inc_15 = a_sel_15 & _inc_T; // @[src/main/scala/tilelink/ToAXI4.scala 269:22]
  wire  dec_15 = d_sel_15 & d_last & _dec_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 270:32]
  wire  _count_T_62 = count_16 + inc_15; // @[src/main/scala/tilelink/ToAXI4.scala 271:24]
  wire  line_435_clock;
  wire  line_435_reset;
  wire  line_435_valid;
  reg  line_435_valid_reg;
  wire  _T_191 = ~(~dec_15 | count_16); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
  wire  line_436_clock;
  wire  line_436_reset;
  wire  line_436_valid;
  reg  line_436_valid_reg;
  wire  line_437_clock;
  wire  line_437_reset;
  wire  line_437_valid;
  reg  line_437_valid_reg;
  wire  _T_197 = ~(~inc_15 | idle_15); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
  wire  line_438_clock;
  wire  line_438_reset;
  wire  line_438_valid;
  reg  line_438_valid_reg;
  wire  line_439_clock;
  wire  line_439_reset;
  wire  line_439_valid;
  reg  line_439_valid_reg;
  Queue_34 nodeOut_w_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_w_deq_q_clock),
    .reset(nodeOut_w_deq_q_reset),
    .io_enq_ready(nodeOut_w_deq_q_io_enq_ready),
    .io_enq_valid(nodeOut_w_deq_q_io_enq_valid),
    .io_enq_bits_data(nodeOut_w_deq_q_io_enq_bits_data),
    .io_enq_bits_strb(nodeOut_w_deq_q_io_enq_bits_strb),
    .io_enq_bits_last(nodeOut_w_deq_q_io_enq_bits_last),
    .io_deq_ready(nodeOut_w_deq_q_io_deq_ready),
    .io_deq_valid(nodeOut_w_deq_q_io_deq_valid),
    .io_deq_bits_data(nodeOut_w_deq_q_io_deq_bits_data),
    .io_deq_bits_strb(nodeOut_w_deq_q_io_deq_bits_strb),
    .io_deq_bits_last(nodeOut_w_deq_q_io_deq_bits_last)
  );
  Queue_35 queue_arw_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(queue_arw_deq_q_clock),
    .reset(queue_arw_deq_q_reset),
    .io_enq_ready(queue_arw_deq_q_io_enq_ready),
    .io_enq_valid(queue_arw_deq_q_io_enq_valid),
    .io_enq_bits_id(queue_arw_deq_q_io_enq_bits_id),
    .io_enq_bits_addr(queue_arw_deq_q_io_enq_bits_addr),
    .io_enq_bits_len(queue_arw_deq_q_io_enq_bits_len),
    .io_enq_bits_size(queue_arw_deq_q_io_enq_bits_size),
    .io_enq_bits_echo_tl_state_size(queue_arw_deq_q_io_enq_bits_echo_tl_state_size),
    .io_enq_bits_echo_tl_state_source(queue_arw_deq_q_io_enq_bits_echo_tl_state_source),
    .io_enq_bits_wen(queue_arw_deq_q_io_enq_bits_wen),
    .io_deq_ready(queue_arw_deq_q_io_deq_ready),
    .io_deq_valid(queue_arw_deq_q_io_deq_valid),
    .io_deq_bits_id(queue_arw_deq_q_io_deq_bits_id),
    .io_deq_bits_addr(queue_arw_deq_q_io_deq_bits_addr),
    .io_deq_bits_len(queue_arw_deq_q_io_deq_bits_len),
    .io_deq_bits_size(queue_arw_deq_q_io_deq_bits_size),
    .io_deq_bits_burst(queue_arw_deq_q_io_deq_bits_burst),
    .io_deq_bits_echo_tl_state_size(queue_arw_deq_q_io_deq_bits_echo_tl_state_size),
    .io_deq_bits_echo_tl_state_source(queue_arw_deq_q_io_deq_bits_echo_tl_state_source),
    .io_deq_bits_wen(queue_arw_deq_q_io_deq_bits_wen)
  );
  GEN_w1_line #(.COVER_INDEX(321)) line_321 (
    .clock(line_321_clock),
    .reset(line_321_reset),
    .valid(line_321_valid)
  );
  GEN_w1_line #(.COVER_INDEX(322)) line_322 (
    .clock(line_322_clock),
    .reset(line_322_reset),
    .valid(line_322_valid)
  );
  GEN_w1_line #(.COVER_INDEX(323)) line_323 (
    .clock(line_323_clock),
    .reset(line_323_reset),
    .valid(line_323_valid)
  );
  GEN_w1_line #(.COVER_INDEX(324)) line_324 (
    .clock(line_324_clock),
    .reset(line_324_reset),
    .valid(line_324_valid)
  );
  GEN_w1_line #(.COVER_INDEX(325)) line_325 (
    .clock(line_325_clock),
    .reset(line_325_reset),
    .valid(line_325_valid)
  );
  GEN_w1_line #(.COVER_INDEX(326)) line_326 (
    .clock(line_326_clock),
    .reset(line_326_reset),
    .valid(line_326_valid)
  );
  GEN_w1_line #(.COVER_INDEX(327)) line_327 (
    .clock(line_327_clock),
    .reset(line_327_reset),
    .valid(line_327_valid)
  );
  GEN_w1_line #(.COVER_INDEX(328)) line_328 (
    .clock(line_328_clock),
    .reset(line_328_reset),
    .valid(line_328_valid)
  );
  GEN_w1_line #(.COVER_INDEX(329)) line_329 (
    .clock(line_329_clock),
    .reset(line_329_reset),
    .valid(line_329_valid)
  );
  GEN_w1_line #(.COVER_INDEX(330)) line_330 (
    .clock(line_330_clock),
    .reset(line_330_reset),
    .valid(line_330_valid)
  );
  GEN_w1_line #(.COVER_INDEX(331)) line_331 (
    .clock(line_331_clock),
    .reset(line_331_reset),
    .valid(line_331_valid)
  );
  GEN_w1_line #(.COVER_INDEX(332)) line_332 (
    .clock(line_332_clock),
    .reset(line_332_reset),
    .valid(line_332_valid)
  );
  GEN_w1_line #(.COVER_INDEX(333)) line_333 (
    .clock(line_333_clock),
    .reset(line_333_reset),
    .valid(line_333_valid)
  );
  GEN_w1_line #(.COVER_INDEX(334)) line_334 (
    .clock(line_334_clock),
    .reset(line_334_reset),
    .valid(line_334_valid)
  );
  GEN_w1_line #(.COVER_INDEX(335)) line_335 (
    .clock(line_335_clock),
    .reset(line_335_reset),
    .valid(line_335_valid)
  );
  GEN_w1_line #(.COVER_INDEX(336)) line_336 (
    .clock(line_336_clock),
    .reset(line_336_reset),
    .valid(line_336_valid)
  );
  GEN_w1_line #(.COVER_INDEX(337)) line_337 (
    .clock(line_337_clock),
    .reset(line_337_reset),
    .valid(line_337_valid)
  );
  GEN_w1_line #(.COVER_INDEX(338)) line_338 (
    .clock(line_338_clock),
    .reset(line_338_reset),
    .valid(line_338_valid)
  );
  GEN_w1_line #(.COVER_INDEX(339)) line_339 (
    .clock(line_339_clock),
    .reset(line_339_reset),
    .valid(line_339_valid)
  );
  GEN_w1_line #(.COVER_INDEX(340)) line_340 (
    .clock(line_340_clock),
    .reset(line_340_reset),
    .valid(line_340_valid)
  );
  GEN_w1_line #(.COVER_INDEX(341)) line_341 (
    .clock(line_341_clock),
    .reset(line_341_reset),
    .valid(line_341_valid)
  );
  GEN_w1_line #(.COVER_INDEX(342)) line_342 (
    .clock(line_342_clock),
    .reset(line_342_reset),
    .valid(line_342_valid)
  );
  GEN_w1_line #(.COVER_INDEX(343)) line_343 (
    .clock(line_343_clock),
    .reset(line_343_reset),
    .valid(line_343_valid)
  );
  GEN_w1_line #(.COVER_INDEX(344)) line_344 (
    .clock(line_344_clock),
    .reset(line_344_reset),
    .valid(line_344_valid)
  );
  GEN_w1_line #(.COVER_INDEX(345)) line_345 (
    .clock(line_345_clock),
    .reset(line_345_reset),
    .valid(line_345_valid)
  );
  GEN_w1_line #(.COVER_INDEX(346)) line_346 (
    .clock(line_346_clock),
    .reset(line_346_reset),
    .valid(line_346_valid)
  );
  GEN_w1_line #(.COVER_INDEX(347)) line_347 (
    .clock(line_347_clock),
    .reset(line_347_reset),
    .valid(line_347_valid)
  );
  GEN_w1_line #(.COVER_INDEX(348)) line_348 (
    .clock(line_348_clock),
    .reset(line_348_reset),
    .valid(line_348_valid)
  );
  GEN_w1_line #(.COVER_INDEX(349)) line_349 (
    .clock(line_349_clock),
    .reset(line_349_reset),
    .valid(line_349_valid)
  );
  GEN_w1_line #(.COVER_INDEX(350)) line_350 (
    .clock(line_350_clock),
    .reset(line_350_reset),
    .valid(line_350_valid)
  );
  GEN_w1_line #(.COVER_INDEX(351)) line_351 (
    .clock(line_351_clock),
    .reset(line_351_reset),
    .valid(line_351_valid)
  );
  GEN_w1_line #(.COVER_INDEX(352)) line_352 (
    .clock(line_352_clock),
    .reset(line_352_reset),
    .valid(line_352_valid)
  );
  GEN_w1_line #(.COVER_INDEX(353)) line_353 (
    .clock(line_353_clock),
    .reset(line_353_reset),
    .valid(line_353_valid)
  );
  GEN_w1_line #(.COVER_INDEX(354)) line_354 (
    .clock(line_354_clock),
    .reset(line_354_reset),
    .valid(line_354_valid)
  );
  GEN_w1_line #(.COVER_INDEX(355)) line_355 (
    .clock(line_355_clock),
    .reset(line_355_reset),
    .valid(line_355_valid)
  );
  GEN_w1_line #(.COVER_INDEX(356)) line_356 (
    .clock(line_356_clock),
    .reset(line_356_reset),
    .valid(line_356_valid)
  );
  GEN_w1_line #(.COVER_INDEX(357)) line_357 (
    .clock(line_357_clock),
    .reset(line_357_reset),
    .valid(line_357_valid)
  );
  GEN_w1_line #(.COVER_INDEX(358)) line_358 (
    .clock(line_358_clock),
    .reset(line_358_reset),
    .valid(line_358_valid)
  );
  GEN_w1_line #(.COVER_INDEX(359)) line_359 (
    .clock(line_359_clock),
    .reset(line_359_reset),
    .valid(line_359_valid)
  );
  GEN_w1_line #(.COVER_INDEX(360)) line_360 (
    .clock(line_360_clock),
    .reset(line_360_reset),
    .valid(line_360_valid)
  );
  GEN_w1_line #(.COVER_INDEX(361)) line_361 (
    .clock(line_361_clock),
    .reset(line_361_reset),
    .valid(line_361_valid)
  );
  GEN_w1_line #(.COVER_INDEX(362)) line_362 (
    .clock(line_362_clock),
    .reset(line_362_reset),
    .valid(line_362_valid)
  );
  GEN_w1_line #(.COVER_INDEX(363)) line_363 (
    .clock(line_363_clock),
    .reset(line_363_reset),
    .valid(line_363_valid)
  );
  GEN_w1_line #(.COVER_INDEX(364)) line_364 (
    .clock(line_364_clock),
    .reset(line_364_reset),
    .valid(line_364_valid)
  );
  GEN_w1_line #(.COVER_INDEX(365)) line_365 (
    .clock(line_365_clock),
    .reset(line_365_reset),
    .valid(line_365_valid)
  );
  GEN_w1_line #(.COVER_INDEX(366)) line_366 (
    .clock(line_366_clock),
    .reset(line_366_reset),
    .valid(line_366_valid)
  );
  GEN_w1_line #(.COVER_INDEX(367)) line_367 (
    .clock(line_367_clock),
    .reset(line_367_reset),
    .valid(line_367_valid)
  );
  GEN_w1_line #(.COVER_INDEX(368)) line_368 (
    .clock(line_368_clock),
    .reset(line_368_reset),
    .valid(line_368_valid)
  );
  GEN_w1_line #(.COVER_INDEX(369)) line_369 (
    .clock(line_369_clock),
    .reset(line_369_reset),
    .valid(line_369_valid)
  );
  GEN_w1_line #(.COVER_INDEX(370)) line_370 (
    .clock(line_370_clock),
    .reset(line_370_reset),
    .valid(line_370_valid)
  );
  GEN_w1_line #(.COVER_INDEX(371)) line_371 (
    .clock(line_371_clock),
    .reset(line_371_reset),
    .valid(line_371_valid)
  );
  GEN_w1_line #(.COVER_INDEX(372)) line_372 (
    .clock(line_372_clock),
    .reset(line_372_reset),
    .valid(line_372_valid)
  );
  GEN_w1_line #(.COVER_INDEX(373)) line_373 (
    .clock(line_373_clock),
    .reset(line_373_reset),
    .valid(line_373_valid)
  );
  GEN_w1_line #(.COVER_INDEX(374)) line_374 (
    .clock(line_374_clock),
    .reset(line_374_reset),
    .valid(line_374_valid)
  );
  GEN_w1_line #(.COVER_INDEX(375)) line_375 (
    .clock(line_375_clock),
    .reset(line_375_reset),
    .valid(line_375_valid)
  );
  GEN_w1_line #(.COVER_INDEX(376)) line_376 (
    .clock(line_376_clock),
    .reset(line_376_reset),
    .valid(line_376_valid)
  );
  GEN_w1_line #(.COVER_INDEX(377)) line_377 (
    .clock(line_377_clock),
    .reset(line_377_reset),
    .valid(line_377_valid)
  );
  GEN_w1_line #(.COVER_INDEX(378)) line_378 (
    .clock(line_378_clock),
    .reset(line_378_reset),
    .valid(line_378_valid)
  );
  GEN_w1_line #(.COVER_INDEX(379)) line_379 (
    .clock(line_379_clock),
    .reset(line_379_reset),
    .valid(line_379_valid)
  );
  GEN_w1_line #(.COVER_INDEX(380)) line_380 (
    .clock(line_380_clock),
    .reset(line_380_reset),
    .valid(line_380_valid)
  );
  GEN_w1_line #(.COVER_INDEX(381)) line_381 (
    .clock(line_381_clock),
    .reset(line_381_reset),
    .valid(line_381_valid)
  );
  GEN_w1_line #(.COVER_INDEX(382)) line_382 (
    .clock(line_382_clock),
    .reset(line_382_reset),
    .valid(line_382_valid)
  );
  GEN_w1_line #(.COVER_INDEX(383)) line_383 (
    .clock(line_383_clock),
    .reset(line_383_reset),
    .valid(line_383_valid)
  );
  GEN_w1_line #(.COVER_INDEX(384)) line_384 (
    .clock(line_384_clock),
    .reset(line_384_reset),
    .valid(line_384_valid)
  );
  GEN_w1_line #(.COVER_INDEX(385)) line_385 (
    .clock(line_385_clock),
    .reset(line_385_reset),
    .valid(line_385_valid)
  );
  GEN_w1_line #(.COVER_INDEX(386)) line_386 (
    .clock(line_386_clock),
    .reset(line_386_reset),
    .valid(line_386_valid)
  );
  GEN_w1_line #(.COVER_INDEX(387)) line_387 (
    .clock(line_387_clock),
    .reset(line_387_reset),
    .valid(line_387_valid)
  );
  GEN_w1_line #(.COVER_INDEX(388)) line_388 (
    .clock(line_388_clock),
    .reset(line_388_reset),
    .valid(line_388_valid)
  );
  GEN_w1_line #(.COVER_INDEX(389)) line_389 (
    .clock(line_389_clock),
    .reset(line_389_reset),
    .valid(line_389_valid)
  );
  GEN_w1_line #(.COVER_INDEX(390)) line_390 (
    .clock(line_390_clock),
    .reset(line_390_reset),
    .valid(line_390_valid)
  );
  GEN_w1_line #(.COVER_INDEX(391)) line_391 (
    .clock(line_391_clock),
    .reset(line_391_reset),
    .valid(line_391_valid)
  );
  GEN_w1_line #(.COVER_INDEX(392)) line_392 (
    .clock(line_392_clock),
    .reset(line_392_reset),
    .valid(line_392_valid)
  );
  GEN_w1_line #(.COVER_INDEX(393)) line_393 (
    .clock(line_393_clock),
    .reset(line_393_reset),
    .valid(line_393_valid)
  );
  GEN_w1_line #(.COVER_INDEX(394)) line_394 (
    .clock(line_394_clock),
    .reset(line_394_reset),
    .valid(line_394_valid)
  );
  GEN_w1_line #(.COVER_INDEX(395)) line_395 (
    .clock(line_395_clock),
    .reset(line_395_reset),
    .valid(line_395_valid)
  );
  GEN_w1_line #(.COVER_INDEX(396)) line_396 (
    .clock(line_396_clock),
    .reset(line_396_reset),
    .valid(line_396_valid)
  );
  GEN_w1_line #(.COVER_INDEX(397)) line_397 (
    .clock(line_397_clock),
    .reset(line_397_reset),
    .valid(line_397_valid)
  );
  GEN_w1_line #(.COVER_INDEX(398)) line_398 (
    .clock(line_398_clock),
    .reset(line_398_reset),
    .valid(line_398_valid)
  );
  GEN_w1_line #(.COVER_INDEX(399)) line_399 (
    .clock(line_399_clock),
    .reset(line_399_reset),
    .valid(line_399_valid)
  );
  GEN_w1_line #(.COVER_INDEX(400)) line_400 (
    .clock(line_400_clock),
    .reset(line_400_reset),
    .valid(line_400_valid)
  );
  GEN_w1_line #(.COVER_INDEX(401)) line_401 (
    .clock(line_401_clock),
    .reset(line_401_reset),
    .valid(line_401_valid)
  );
  GEN_w1_line #(.COVER_INDEX(402)) line_402 (
    .clock(line_402_clock),
    .reset(line_402_reset),
    .valid(line_402_valid)
  );
  GEN_w1_line #(.COVER_INDEX(403)) line_403 (
    .clock(line_403_clock),
    .reset(line_403_reset),
    .valid(line_403_valid)
  );
  GEN_w1_line #(.COVER_INDEX(404)) line_404 (
    .clock(line_404_clock),
    .reset(line_404_reset),
    .valid(line_404_valid)
  );
  GEN_w1_line #(.COVER_INDEX(405)) line_405 (
    .clock(line_405_clock),
    .reset(line_405_reset),
    .valid(line_405_valid)
  );
  GEN_w1_line #(.COVER_INDEX(406)) line_406 (
    .clock(line_406_clock),
    .reset(line_406_reset),
    .valid(line_406_valid)
  );
  GEN_w1_line #(.COVER_INDEX(407)) line_407 (
    .clock(line_407_clock),
    .reset(line_407_reset),
    .valid(line_407_valid)
  );
  GEN_w1_line #(.COVER_INDEX(408)) line_408 (
    .clock(line_408_clock),
    .reset(line_408_reset),
    .valid(line_408_valid)
  );
  GEN_w1_line #(.COVER_INDEX(409)) line_409 (
    .clock(line_409_clock),
    .reset(line_409_reset),
    .valid(line_409_valid)
  );
  GEN_w1_line #(.COVER_INDEX(410)) line_410 (
    .clock(line_410_clock),
    .reset(line_410_reset),
    .valid(line_410_valid)
  );
  GEN_w1_line #(.COVER_INDEX(411)) line_411 (
    .clock(line_411_clock),
    .reset(line_411_reset),
    .valid(line_411_valid)
  );
  GEN_w1_line #(.COVER_INDEX(412)) line_412 (
    .clock(line_412_clock),
    .reset(line_412_reset),
    .valid(line_412_valid)
  );
  GEN_w1_line #(.COVER_INDEX(413)) line_413 (
    .clock(line_413_clock),
    .reset(line_413_reset),
    .valid(line_413_valid)
  );
  GEN_w1_line #(.COVER_INDEX(414)) line_414 (
    .clock(line_414_clock),
    .reset(line_414_reset),
    .valid(line_414_valid)
  );
  GEN_w1_line #(.COVER_INDEX(415)) line_415 (
    .clock(line_415_clock),
    .reset(line_415_reset),
    .valid(line_415_valid)
  );
  GEN_w1_line #(.COVER_INDEX(416)) line_416 (
    .clock(line_416_clock),
    .reset(line_416_reset),
    .valid(line_416_valid)
  );
  GEN_w1_line #(.COVER_INDEX(417)) line_417 (
    .clock(line_417_clock),
    .reset(line_417_reset),
    .valid(line_417_valid)
  );
  GEN_w1_line #(.COVER_INDEX(418)) line_418 (
    .clock(line_418_clock),
    .reset(line_418_reset),
    .valid(line_418_valid)
  );
  GEN_w1_line #(.COVER_INDEX(419)) line_419 (
    .clock(line_419_clock),
    .reset(line_419_reset),
    .valid(line_419_valid)
  );
  GEN_w1_line #(.COVER_INDEX(420)) line_420 (
    .clock(line_420_clock),
    .reset(line_420_reset),
    .valid(line_420_valid)
  );
  GEN_w1_line #(.COVER_INDEX(421)) line_421 (
    .clock(line_421_clock),
    .reset(line_421_reset),
    .valid(line_421_valid)
  );
  GEN_w1_line #(.COVER_INDEX(422)) line_422 (
    .clock(line_422_clock),
    .reset(line_422_reset),
    .valid(line_422_valid)
  );
  GEN_w1_line #(.COVER_INDEX(423)) line_423 (
    .clock(line_423_clock),
    .reset(line_423_reset),
    .valid(line_423_valid)
  );
  GEN_w1_line #(.COVER_INDEX(424)) line_424 (
    .clock(line_424_clock),
    .reset(line_424_reset),
    .valid(line_424_valid)
  );
  GEN_w1_line #(.COVER_INDEX(425)) line_425 (
    .clock(line_425_clock),
    .reset(line_425_reset),
    .valid(line_425_valid)
  );
  GEN_w1_line #(.COVER_INDEX(426)) line_426 (
    .clock(line_426_clock),
    .reset(line_426_reset),
    .valid(line_426_valid)
  );
  GEN_w1_line #(.COVER_INDEX(427)) line_427 (
    .clock(line_427_clock),
    .reset(line_427_reset),
    .valid(line_427_valid)
  );
  GEN_w1_line #(.COVER_INDEX(428)) line_428 (
    .clock(line_428_clock),
    .reset(line_428_reset),
    .valid(line_428_valid)
  );
  GEN_w1_line #(.COVER_INDEX(429)) line_429 (
    .clock(line_429_clock),
    .reset(line_429_reset),
    .valid(line_429_valid)
  );
  GEN_w1_line #(.COVER_INDEX(430)) line_430 (
    .clock(line_430_clock),
    .reset(line_430_reset),
    .valid(line_430_valid)
  );
  GEN_w1_line #(.COVER_INDEX(431)) line_431 (
    .clock(line_431_clock),
    .reset(line_431_reset),
    .valid(line_431_valid)
  );
  GEN_w1_line #(.COVER_INDEX(432)) line_432 (
    .clock(line_432_clock),
    .reset(line_432_reset),
    .valid(line_432_valid)
  );
  GEN_w1_line #(.COVER_INDEX(433)) line_433 (
    .clock(line_433_clock),
    .reset(line_433_reset),
    .valid(line_433_valid)
  );
  GEN_w1_line #(.COVER_INDEX(434)) line_434 (
    .clock(line_434_clock),
    .reset(line_434_reset),
    .valid(line_434_valid)
  );
  GEN_w1_line #(.COVER_INDEX(435)) line_435 (
    .clock(line_435_clock),
    .reset(line_435_reset),
    .valid(line_435_valid)
  );
  GEN_w1_line #(.COVER_INDEX(436)) line_436 (
    .clock(line_436_clock),
    .reset(line_436_reset),
    .valid(line_436_valid)
  );
  GEN_w1_line #(.COVER_INDEX(437)) line_437 (
    .clock(line_437_clock),
    .reset(line_437_reset),
    .valid(line_437_valid)
  );
  GEN_w1_line #(.COVER_INDEX(438)) line_438 (
    .clock(line_438_clock),
    .reset(line_438_reset),
    .valid(line_438_valid)
  );
  GEN_w1_line #(.COVER_INDEX(439)) line_439 (
    .clock(line_439_clock),
    .reset(line_439_reset),
    .valid(line_439_valid)
  );
  assign line_321_clock = clock;
  assign line_321_reset = reset;
  assign line_321_valid = _T ^ line_321_valid_reg;
  assign line_322_clock = clock;
  assign line_322_reset = reset;
  assign line_322_valid = _T ^ line_322_valid_reg;
  assign line_323_clock = clock;
  assign line_323_reset = reset;
  assign line_323_valid = 4'h0 == auto_in_a_bits_source ^ line_323_valid_reg;
  assign line_324_clock = clock;
  assign line_324_reset = reset;
  assign line_324_valid = 4'h1 == auto_in_a_bits_source ^ line_324_valid_reg;
  assign line_325_clock = clock;
  assign line_325_reset = reset;
  assign line_325_valid = 4'h2 == auto_in_a_bits_source ^ line_325_valid_reg;
  assign line_326_clock = clock;
  assign line_326_reset = reset;
  assign line_326_valid = 4'h3 == auto_in_a_bits_source ^ line_326_valid_reg;
  assign line_327_clock = clock;
  assign line_327_reset = reset;
  assign line_327_valid = 4'h4 == auto_in_a_bits_source ^ line_327_valid_reg;
  assign line_328_clock = clock;
  assign line_328_reset = reset;
  assign line_328_valid = 4'h5 == auto_in_a_bits_source ^ line_328_valid_reg;
  assign line_329_clock = clock;
  assign line_329_reset = reset;
  assign line_329_valid = 4'h6 == auto_in_a_bits_source ^ line_329_valid_reg;
  assign line_330_clock = clock;
  assign line_330_reset = reset;
  assign line_330_valid = 4'h7 == auto_in_a_bits_source ^ line_330_valid_reg;
  assign line_331_clock = clock;
  assign line_331_reset = reset;
  assign line_331_valid = 4'h8 == auto_in_a_bits_source ^ line_331_valid_reg;
  assign line_332_clock = clock;
  assign line_332_reset = reset;
  assign line_332_valid = 4'h9 == auto_in_a_bits_source ^ line_332_valid_reg;
  assign line_333_clock = clock;
  assign line_333_reset = reset;
  assign line_333_valid = 4'ha == auto_in_a_bits_source ^ line_333_valid_reg;
  assign line_334_clock = clock;
  assign line_334_reset = reset;
  assign line_334_valid = 4'hb == auto_in_a_bits_source ^ line_334_valid_reg;
  assign line_335_clock = clock;
  assign line_335_reset = reset;
  assign line_335_valid = 4'hc == auto_in_a_bits_source ^ line_335_valid_reg;
  assign line_336_clock = clock;
  assign line_336_reset = reset;
  assign line_336_valid = 4'hd == auto_in_a_bits_source ^ line_336_valid_reg;
  assign line_337_clock = clock;
  assign line_337_reset = reset;
  assign line_337_valid = 4'he == auto_in_a_bits_source ^ line_337_valid_reg;
  assign line_338_clock = clock;
  assign line_338_reset = reset;
  assign line_338_valid = 4'hf == auto_in_a_bits_source ^ line_338_valid_reg;
  assign line_339_clock = clock;
  assign line_339_reset = reset;
  assign line_339_valid = 4'h0 == auto_in_a_bits_source ^ line_339_valid_reg;
  assign line_340_clock = clock;
  assign line_340_reset = reset;
  assign line_340_valid = 4'h1 == auto_in_a_bits_source ^ line_340_valid_reg;
  assign line_341_clock = clock;
  assign line_341_reset = reset;
  assign line_341_valid = 4'h2 == auto_in_a_bits_source ^ line_341_valid_reg;
  assign line_342_clock = clock;
  assign line_342_reset = reset;
  assign line_342_valid = 4'h3 == auto_in_a_bits_source ^ line_342_valid_reg;
  assign line_343_clock = clock;
  assign line_343_reset = reset;
  assign line_343_valid = 4'h4 == auto_in_a_bits_source ^ line_343_valid_reg;
  assign line_344_clock = clock;
  assign line_344_reset = reset;
  assign line_344_valid = 4'h5 == auto_in_a_bits_source ^ line_344_valid_reg;
  assign line_345_clock = clock;
  assign line_345_reset = reset;
  assign line_345_valid = 4'h6 == auto_in_a_bits_source ^ line_345_valid_reg;
  assign line_346_clock = clock;
  assign line_346_reset = reset;
  assign line_346_valid = 4'h7 == auto_in_a_bits_source ^ line_346_valid_reg;
  assign line_347_clock = clock;
  assign line_347_reset = reset;
  assign line_347_valid = 4'h8 == auto_in_a_bits_source ^ line_347_valid_reg;
  assign line_348_clock = clock;
  assign line_348_reset = reset;
  assign line_348_valid = 4'h9 == auto_in_a_bits_source ^ line_348_valid_reg;
  assign line_349_clock = clock;
  assign line_349_reset = reset;
  assign line_349_valid = 4'ha == auto_in_a_bits_source ^ line_349_valid_reg;
  assign line_350_clock = clock;
  assign line_350_reset = reset;
  assign line_350_valid = 4'hb == auto_in_a_bits_source ^ line_350_valid_reg;
  assign line_351_clock = clock;
  assign line_351_reset = reset;
  assign line_351_valid = 4'hc == auto_in_a_bits_source ^ line_351_valid_reg;
  assign line_352_clock = clock;
  assign line_352_reset = reset;
  assign line_352_valid = 4'hd == auto_in_a_bits_source ^ line_352_valid_reg;
  assign line_353_clock = clock;
  assign line_353_reset = reset;
  assign line_353_valid = 4'he == auto_in_a_bits_source ^ line_353_valid_reg;
  assign line_354_clock = clock;
  assign line_354_reset = reset;
  assign line_354_valid = 4'hf == auto_in_a_bits_source ^ line_354_valid_reg;
  assign line_355_clock = clock;
  assign line_355_reset = reset;
  assign line_355_valid = _T_2 ^ line_355_valid_reg;
  assign line_356_clock = clock;
  assign line_356_reset = reset;
  assign line_356_valid = _T_4 ^ line_356_valid_reg;
  assign line_357_clock = clock;
  assign line_357_reset = reset;
  assign line_357_valid = _T_4 ^ line_357_valid_reg;
  assign line_358_clock = clock;
  assign line_358_reset = reset;
  assign line_358_valid = _T_2 ^ line_358_valid_reg;
  assign line_359_clock = clock;
  assign line_359_reset = reset;
  assign line_359_valid = r_first ^ line_359_valid_reg;
  assign line_360_clock = clock;
  assign line_360_reset = reset;
  assign line_360_valid = _T_10 ^ line_360_valid_reg;
  assign line_361_clock = clock;
  assign line_361_reset = reset;
  assign line_361_valid = _T_11 ^ line_361_valid_reg;
  assign line_362_clock = clock;
  assign line_362_reset = reset;
  assign line_362_valid = _T_10 ^ line_362_valid_reg;
  assign line_363_clock = clock;
  assign line_363_reset = reset;
  assign line_363_valid = _T_17 ^ line_363_valid_reg;
  assign line_364_clock = clock;
  assign line_364_reset = reset;
  assign line_364_valid = inc ^ line_364_valid_reg;
  assign line_365_clock = clock;
  assign line_365_reset = reset;
  assign line_365_valid = _T_10 ^ line_365_valid_reg;
  assign line_366_clock = clock;
  assign line_366_reset = reset;
  assign line_366_valid = _T_23 ^ line_366_valid_reg;
  assign line_367_clock = clock;
  assign line_367_reset = reset;
  assign line_367_valid = _T_10 ^ line_367_valid_reg;
  assign line_368_clock = clock;
  assign line_368_reset = reset;
  assign line_368_valid = _T_29 ^ line_368_valid_reg;
  assign line_369_clock = clock;
  assign line_369_reset = reset;
  assign line_369_valid = inc_1 ^ line_369_valid_reg;
  assign line_370_clock = clock;
  assign line_370_reset = reset;
  assign line_370_valid = _T_10 ^ line_370_valid_reg;
  assign line_371_clock = clock;
  assign line_371_reset = reset;
  assign line_371_valid = _T_35 ^ line_371_valid_reg;
  assign line_372_clock = clock;
  assign line_372_reset = reset;
  assign line_372_valid = _T_10 ^ line_372_valid_reg;
  assign line_373_clock = clock;
  assign line_373_reset = reset;
  assign line_373_valid = _T_41 ^ line_373_valid_reg;
  assign line_374_clock = clock;
  assign line_374_reset = reset;
  assign line_374_valid = inc_2 ^ line_374_valid_reg;
  assign line_375_clock = clock;
  assign line_375_reset = reset;
  assign line_375_valid = _T_10 ^ line_375_valid_reg;
  assign line_376_clock = clock;
  assign line_376_reset = reset;
  assign line_376_valid = _T_47 ^ line_376_valid_reg;
  assign line_377_clock = clock;
  assign line_377_reset = reset;
  assign line_377_valid = _T_10 ^ line_377_valid_reg;
  assign line_378_clock = clock;
  assign line_378_reset = reset;
  assign line_378_valid = _T_53 ^ line_378_valid_reg;
  assign line_379_clock = clock;
  assign line_379_reset = reset;
  assign line_379_valid = inc_3 ^ line_379_valid_reg;
  assign line_380_clock = clock;
  assign line_380_reset = reset;
  assign line_380_valid = _T_10 ^ line_380_valid_reg;
  assign line_381_clock = clock;
  assign line_381_reset = reset;
  assign line_381_valid = _T_59 ^ line_381_valid_reg;
  assign line_382_clock = clock;
  assign line_382_reset = reset;
  assign line_382_valid = _T_10 ^ line_382_valid_reg;
  assign line_383_clock = clock;
  assign line_383_reset = reset;
  assign line_383_valid = _T_65 ^ line_383_valid_reg;
  assign line_384_clock = clock;
  assign line_384_reset = reset;
  assign line_384_valid = inc_4 ^ line_384_valid_reg;
  assign line_385_clock = clock;
  assign line_385_reset = reset;
  assign line_385_valid = _T_10 ^ line_385_valid_reg;
  assign line_386_clock = clock;
  assign line_386_reset = reset;
  assign line_386_valid = _T_71 ^ line_386_valid_reg;
  assign line_387_clock = clock;
  assign line_387_reset = reset;
  assign line_387_valid = _T_10 ^ line_387_valid_reg;
  assign line_388_clock = clock;
  assign line_388_reset = reset;
  assign line_388_valid = _T_77 ^ line_388_valid_reg;
  assign line_389_clock = clock;
  assign line_389_reset = reset;
  assign line_389_valid = inc_5 ^ line_389_valid_reg;
  assign line_390_clock = clock;
  assign line_390_reset = reset;
  assign line_390_valid = _T_10 ^ line_390_valid_reg;
  assign line_391_clock = clock;
  assign line_391_reset = reset;
  assign line_391_valid = _T_83 ^ line_391_valid_reg;
  assign line_392_clock = clock;
  assign line_392_reset = reset;
  assign line_392_valid = _T_10 ^ line_392_valid_reg;
  assign line_393_clock = clock;
  assign line_393_reset = reset;
  assign line_393_valid = _T_89 ^ line_393_valid_reg;
  assign line_394_clock = clock;
  assign line_394_reset = reset;
  assign line_394_valid = inc_6 ^ line_394_valid_reg;
  assign line_395_clock = clock;
  assign line_395_reset = reset;
  assign line_395_valid = _T_10 ^ line_395_valid_reg;
  assign line_396_clock = clock;
  assign line_396_reset = reset;
  assign line_396_valid = _T_95 ^ line_396_valid_reg;
  assign line_397_clock = clock;
  assign line_397_reset = reset;
  assign line_397_valid = _T_10 ^ line_397_valid_reg;
  assign line_398_clock = clock;
  assign line_398_reset = reset;
  assign line_398_valid = _T_101 ^ line_398_valid_reg;
  assign line_399_clock = clock;
  assign line_399_reset = reset;
  assign line_399_valid = inc_7 ^ line_399_valid_reg;
  assign line_400_clock = clock;
  assign line_400_reset = reset;
  assign line_400_valid = _T_10 ^ line_400_valid_reg;
  assign line_401_clock = clock;
  assign line_401_reset = reset;
  assign line_401_valid = _T_107 ^ line_401_valid_reg;
  assign line_402_clock = clock;
  assign line_402_reset = reset;
  assign line_402_valid = _T_10 ^ line_402_valid_reg;
  assign line_403_clock = clock;
  assign line_403_reset = reset;
  assign line_403_valid = _T_113 ^ line_403_valid_reg;
  assign line_404_clock = clock;
  assign line_404_reset = reset;
  assign line_404_valid = inc_8 ^ line_404_valid_reg;
  assign line_405_clock = clock;
  assign line_405_reset = reset;
  assign line_405_valid = _T_10 ^ line_405_valid_reg;
  assign line_406_clock = clock;
  assign line_406_reset = reset;
  assign line_406_valid = _T_119 ^ line_406_valid_reg;
  assign line_407_clock = clock;
  assign line_407_reset = reset;
  assign line_407_valid = _T_10 ^ line_407_valid_reg;
  assign line_408_clock = clock;
  assign line_408_reset = reset;
  assign line_408_valid = _T_125 ^ line_408_valid_reg;
  assign line_409_clock = clock;
  assign line_409_reset = reset;
  assign line_409_valid = inc_9 ^ line_409_valid_reg;
  assign line_410_clock = clock;
  assign line_410_reset = reset;
  assign line_410_valid = _T_10 ^ line_410_valid_reg;
  assign line_411_clock = clock;
  assign line_411_reset = reset;
  assign line_411_valid = _T_131 ^ line_411_valid_reg;
  assign line_412_clock = clock;
  assign line_412_reset = reset;
  assign line_412_valid = _T_10 ^ line_412_valid_reg;
  assign line_413_clock = clock;
  assign line_413_reset = reset;
  assign line_413_valid = _T_137 ^ line_413_valid_reg;
  assign line_414_clock = clock;
  assign line_414_reset = reset;
  assign line_414_valid = inc_10 ^ line_414_valid_reg;
  assign line_415_clock = clock;
  assign line_415_reset = reset;
  assign line_415_valid = _T_10 ^ line_415_valid_reg;
  assign line_416_clock = clock;
  assign line_416_reset = reset;
  assign line_416_valid = _T_143 ^ line_416_valid_reg;
  assign line_417_clock = clock;
  assign line_417_reset = reset;
  assign line_417_valid = _T_10 ^ line_417_valid_reg;
  assign line_418_clock = clock;
  assign line_418_reset = reset;
  assign line_418_valid = _T_149 ^ line_418_valid_reg;
  assign line_419_clock = clock;
  assign line_419_reset = reset;
  assign line_419_valid = inc_11 ^ line_419_valid_reg;
  assign line_420_clock = clock;
  assign line_420_reset = reset;
  assign line_420_valid = _T_10 ^ line_420_valid_reg;
  assign line_421_clock = clock;
  assign line_421_reset = reset;
  assign line_421_valid = _T_155 ^ line_421_valid_reg;
  assign line_422_clock = clock;
  assign line_422_reset = reset;
  assign line_422_valid = _T_10 ^ line_422_valid_reg;
  assign line_423_clock = clock;
  assign line_423_reset = reset;
  assign line_423_valid = _T_161 ^ line_423_valid_reg;
  assign line_424_clock = clock;
  assign line_424_reset = reset;
  assign line_424_valid = inc_12 ^ line_424_valid_reg;
  assign line_425_clock = clock;
  assign line_425_reset = reset;
  assign line_425_valid = _T_10 ^ line_425_valid_reg;
  assign line_426_clock = clock;
  assign line_426_reset = reset;
  assign line_426_valid = _T_167 ^ line_426_valid_reg;
  assign line_427_clock = clock;
  assign line_427_reset = reset;
  assign line_427_valid = _T_10 ^ line_427_valid_reg;
  assign line_428_clock = clock;
  assign line_428_reset = reset;
  assign line_428_valid = _T_173 ^ line_428_valid_reg;
  assign line_429_clock = clock;
  assign line_429_reset = reset;
  assign line_429_valid = inc_13 ^ line_429_valid_reg;
  assign line_430_clock = clock;
  assign line_430_reset = reset;
  assign line_430_valid = _T_10 ^ line_430_valid_reg;
  assign line_431_clock = clock;
  assign line_431_reset = reset;
  assign line_431_valid = _T_179 ^ line_431_valid_reg;
  assign line_432_clock = clock;
  assign line_432_reset = reset;
  assign line_432_valid = _T_10 ^ line_432_valid_reg;
  assign line_433_clock = clock;
  assign line_433_reset = reset;
  assign line_433_valid = _T_185 ^ line_433_valid_reg;
  assign line_434_clock = clock;
  assign line_434_reset = reset;
  assign line_434_valid = inc_14 ^ line_434_valid_reg;
  assign line_435_clock = clock;
  assign line_435_reset = reset;
  assign line_435_valid = _T_10 ^ line_435_valid_reg;
  assign line_436_clock = clock;
  assign line_436_reset = reset;
  assign line_436_valid = _T_191 ^ line_436_valid_reg;
  assign line_437_clock = clock;
  assign line_437_reset = reset;
  assign line_437_valid = _T_10 ^ line_437_valid_reg;
  assign line_438_clock = clock;
  assign line_438_reset = reset;
  assign line_438_valid = _T_197 ^ line_438_valid_reg;
  assign line_439_clock = clock;
  assign line_439_reset = reset;
  assign line_439_valid = inc_15 ^ line_439_valid_reg;
  assign auto_in_a_ready = ~stall & _nodeIn_a_ready_T_3; // @[src/main/scala/tilelink/ToAXI4.scala 199:28]
  assign auto_in_d_valid = r_wins ? auto_out_r_valid : auto_out_b_valid; // @[src/main/scala/tilelink/ToAXI4.scala 222:24]
  assign auto_in_d_bits_opcode = r_wins ? 3'h1 : 3'h0; // @[src/main/scala/tilelink/ToAXI4.scala 248:23]
  assign auto_in_d_bits_size = r_wins ? r_d_size : b_d_size; // @[src/main/scala/tilelink/ToAXI4.scala 248:23]
  assign auto_in_d_bits_source = r_wins ? auto_out_r_bits_echo_tl_state_source : auto_out_b_bits_echo_tl_state_source; // @[src/main/scala/tilelink/ToAXI4.scala 248:23]
  assign auto_in_d_bits_denied = r_wins ? _GEN_156 : b_denied; // @[src/main/scala/tilelink/ToAXI4.scala 248:23]
  assign auto_in_d_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = r_wins & r_d_corrupt; // @[src/main/scala/tilelink/ToAXI4.scala 248:23]
  assign auto_out_aw_valid = queue_arw_valid & queue_arw_bits_wen; // @[src/main/scala/tilelink/ToAXI4.scala 155:39]
  assign auto_out_aw_bits_id = queue_arw_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_addr = queue_arw_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_len = queue_arw_deq_q_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_size = queue_arw_deq_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_burst = queue_arw_deq_q_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_echo_tl_state_size = queue_arw_deq_q_io_deq_bits_echo_tl_state_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_echo_tl_state_source = queue_arw_deq_q_io_deq_bits_echo_tl_state_source; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_valid = nodeOut_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_out_w_bits_data = nodeOut_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_bits_strb = nodeOut_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_bits_last = nodeOut_w_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_b_ready = auto_in_d_ready & ~r_wins; // @[src/main/scala/tilelink/ToAXI4.scala 221:33]
  assign auto_out_ar_valid = queue_arw_valid & ~queue_arw_bits_wen; // @[src/main/scala/tilelink/ToAXI4.scala 154:39]
  assign auto_out_ar_bits_id = queue_arw_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_addr = queue_arw_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_len = queue_arw_deq_q_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_size = queue_arw_deq_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_burst = queue_arw_deq_q_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_echo_tl_state_size = queue_arw_deq_q_io_deq_bits_echo_tl_state_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_echo_tl_state_source = queue_arw_deq_q_io_deq_bits_echo_tl_state_source; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_r_ready = auto_in_d_ready & r_wins; // @[src/main/scala/tilelink/ToAXI4.scala 220:33]
  assign nodeOut_w_deq_q_clock = clock;
  assign nodeOut_w_deq_q_reset = reset;
  assign nodeOut_w_deq_q_io_enq_valid = _out_arw_valid_T_1 & a_isPut & _nodeIn_a_ready_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 202:54]
  assign nodeOut_w_deq_q_io_enq_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_w_deq_q_io_enq_bits_strb = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_w_deq_q_io_enq_bits_last = counter == 2'h1 | beats1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  assign nodeOut_w_deq_q_io_deq_ready = auto_out_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign queue_arw_deq_q_clock = clock;
  assign queue_arw_deq_q_reset = reset;
  assign queue_arw_deq_q_io_enq_valid = _nodeIn_a_ready_T & auto_in_a_valid & _out_arw_valid_T_4; // @[src/main/scala/tilelink/ToAXI4.scala 200:45]
  assign queue_arw_deq_q_io_enq_bits_id = 4'hf == auto_in_a_bits_source ? 4'hf : _GEN_135; // @[src/main/scala/tilelink/ToAXI4.scala 165:{17,17}]
  assign queue_arw_deq_q_io_enq_bits_addr = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign queue_arw_deq_q_io_enq_bits_len = _out_arw_bits_len_T_3[10:3]; // @[src/main/scala/tilelink/ToAXI4.scala 167:84]
  assign queue_arw_deq_q_io_enq_bits_size = auto_in_a_bits_size >= 3'h3 ? 3'h3 : auto_in_a_bits_size; // @[src/main/scala/tilelink/ToAXI4.scala 168:23]
  assign queue_arw_deq_q_io_enq_bits_echo_tl_state_size = {{1'd0}, auto_in_a_bits_size}; // @[src/main/scala/tilelink/ToAXI4.scala 146:25 182:22]
  assign queue_arw_deq_q_io_enq_bits_echo_tl_state_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign queue_arw_deq_q_io_enq_bits_wen = ~auto_in_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  assign queue_arw_deq_q_io_deq_ready = queue_arw_bits_wen ? auto_out_aw_ready : auto_out_ar_ready; // @[src/main/scala/tilelink/ToAXI4.scala 156:29]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_16 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_16 <= _count_T_62 - dec_15; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_15 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_15 <= _count_T_58 - dec_14; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_14 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_14 <= _count_T_54 - dec_13; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_13 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_13 <= _count_T_50 - dec_12; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_12 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_12 <= _count_T_46 - dec_11; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_11 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_11 <= _count_T_42 - dec_10; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_10 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_10 <= _count_T_38 - dec_9; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_9 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_9 <= _count_T_34 - dec_8; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_8 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_8 <= _count_T_30 - dec_7; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_7 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_7 <= _count_T_26 - dec_6; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_6 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_6 <= _count_T_22 - dec_5; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_5 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_5 <= _count_T_18 - dec_4; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_4 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_4 <= _count_T_14 - dec_3; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_3 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_3 <= _count_T_10 - dec_2; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_2 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_2 <= _count_T_6 - dec_1; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
      count_1 <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 265:28]
    end else begin
      count_1 <= _count_T_2 - dec; // @[src/main/scala/tilelink/ToAXI4.scala 271:15]
    end
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (a_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (a_isPut) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          counter <= beats1_decode;
        end else begin
          counter <= 2'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 160:30]
      doneAW <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 160:30]
    end else if (_T) begin // @[src/main/scala/tilelink/ToAXI4.scala 161:24]
      doneAW <= ~a_last; // @[src/main/scala/tilelink/ToAXI4.scala 161:33]
    end
    line_321_valid_reg <= _T;
    line_322_valid_reg <= _T;
    line_323_valid_reg <= 4'h0 == auto_in_a_bits_source;
    line_324_valid_reg <= 4'h1 == auto_in_a_bits_source;
    line_325_valid_reg <= 4'h2 == auto_in_a_bits_source;
    line_326_valid_reg <= 4'h3 == auto_in_a_bits_source;
    line_327_valid_reg <= 4'h4 == auto_in_a_bits_source;
    line_328_valid_reg <= 4'h5 == auto_in_a_bits_source;
    line_329_valid_reg <= 4'h6 == auto_in_a_bits_source;
    line_330_valid_reg <= 4'h7 == auto_in_a_bits_source;
    line_331_valid_reg <= 4'h8 == auto_in_a_bits_source;
    line_332_valid_reg <= 4'h9 == auto_in_a_bits_source;
    line_333_valid_reg <= 4'ha == auto_in_a_bits_source;
    line_334_valid_reg <= 4'hb == auto_in_a_bits_source;
    line_335_valid_reg <= 4'hc == auto_in_a_bits_source;
    line_336_valid_reg <= 4'hd == auto_in_a_bits_source;
    line_337_valid_reg <= 4'he == auto_in_a_bits_source;
    line_338_valid_reg <= 4'hf == auto_in_a_bits_source;
    line_339_valid_reg <= 4'h0 == auto_in_a_bits_source;
    line_340_valid_reg <= 4'h1 == auto_in_a_bits_source;
    line_341_valid_reg <= 4'h2 == auto_in_a_bits_source;
    line_342_valid_reg <= 4'h3 == auto_in_a_bits_source;
    line_343_valid_reg <= 4'h4 == auto_in_a_bits_source;
    line_344_valid_reg <= 4'h5 == auto_in_a_bits_source;
    line_345_valid_reg <= 4'h6 == auto_in_a_bits_source;
    line_346_valid_reg <= 4'h7 == auto_in_a_bits_source;
    line_347_valid_reg <= 4'h8 == auto_in_a_bits_source;
    line_348_valid_reg <= 4'h9 == auto_in_a_bits_source;
    line_349_valid_reg <= 4'ha == auto_in_a_bits_source;
    line_350_valid_reg <= 4'hb == auto_in_a_bits_source;
    line_351_valid_reg <= 4'hc == auto_in_a_bits_source;
    line_352_valid_reg <= 4'hd == auto_in_a_bits_source;
    line_353_valid_reg <= 4'he == auto_in_a_bits_source;
    line_354_valid_reg <= 4'hf == auto_in_a_bits_source;
    if (reset) begin // @[src/main/scala/tilelink/ToAXI4.scala 209:30]
      r_holds_d <= 1'h0; // @[src/main/scala/tilelink/ToAXI4.scala 209:30]
    end else if (_T_2) begin // @[src/main/scala/tilelink/ToAXI4.scala 210:25]
      r_holds_d <= ~auto_out_r_bits_last; // @[src/main/scala/tilelink/ToAXI4.scala 210:37]
    end
    if (auto_out_b_valid & ~nodeOut_b_ready) begin // @[src/main/scala/tilelink/ToAXI4.scala 213:42]
      b_delay <= _b_delay_T_1; // @[src/main/scala/tilelink/ToAXI4.scala 214:17]
    end else begin
      b_delay <= 3'h0; // @[src/main/scala/tilelink/ToAXI4.scala 216:17]
    end
    line_355_valid_reg <= _T_2;
    line_356_valid_reg <= _T_4;
    line_357_valid_reg <= _T_4;
    r_first <= reset | _GEN_155; // @[src/main/scala/tilelink/ToAXI4.scala 227:{28,28}]
    line_358_valid_reg <= _T_2;
    if (r_first) begin // @[src/main/scala/util/package.scala 80:63]
      r_denied_r <= _r_denied_T; // @[src/main/scala/util/package.scala 80:63]
    end
    line_359_valid_reg <= r_first;
    line_360_valid_reg <= _T_10;
    line_361_valid_reg <= _T_11;
    line_362_valid_reg <= _T_10;
    line_363_valid_reg <= _T_17;
    line_364_valid_reg <= inc;
    line_365_valid_reg <= _T_10;
    line_366_valid_reg <= _T_23;
    line_367_valid_reg <= _T_10;
    line_368_valid_reg <= _T_29;
    line_369_valid_reg <= inc_1;
    line_370_valid_reg <= _T_10;
    line_371_valid_reg <= _T_35;
    line_372_valid_reg <= _T_10;
    line_373_valid_reg <= _T_41;
    line_374_valid_reg <= inc_2;
    line_375_valid_reg <= _T_10;
    line_376_valid_reg <= _T_47;
    line_377_valid_reg <= _T_10;
    line_378_valid_reg <= _T_53;
    line_379_valid_reg <= inc_3;
    line_380_valid_reg <= _T_10;
    line_381_valid_reg <= _T_59;
    line_382_valid_reg <= _T_10;
    line_383_valid_reg <= _T_65;
    line_384_valid_reg <= inc_4;
    line_385_valid_reg <= _T_10;
    line_386_valid_reg <= _T_71;
    line_387_valid_reg <= _T_10;
    line_388_valid_reg <= _T_77;
    line_389_valid_reg <= inc_5;
    line_390_valid_reg <= _T_10;
    line_391_valid_reg <= _T_83;
    line_392_valid_reg <= _T_10;
    line_393_valid_reg <= _T_89;
    line_394_valid_reg <= inc_6;
    line_395_valid_reg <= _T_10;
    line_396_valid_reg <= _T_95;
    line_397_valid_reg <= _T_10;
    line_398_valid_reg <= _T_101;
    line_399_valid_reg <= inc_7;
    line_400_valid_reg <= _T_10;
    line_401_valid_reg <= _T_107;
    line_402_valid_reg <= _T_10;
    line_403_valid_reg <= _T_113;
    line_404_valid_reg <= inc_8;
    line_405_valid_reg <= _T_10;
    line_406_valid_reg <= _T_119;
    line_407_valid_reg <= _T_10;
    line_408_valid_reg <= _T_125;
    line_409_valid_reg <= inc_9;
    line_410_valid_reg <= _T_10;
    line_411_valid_reg <= _T_131;
    line_412_valid_reg <= _T_10;
    line_413_valid_reg <= _T_137;
    line_414_valid_reg <= inc_10;
    line_415_valid_reg <= _T_10;
    line_416_valid_reg <= _T_143;
    line_417_valid_reg <= _T_10;
    line_418_valid_reg <= _T_149;
    line_419_valid_reg <= inc_11;
    line_420_valid_reg <= _T_10;
    line_421_valid_reg <= _T_155;
    line_422_valid_reg <= _T_10;
    line_423_valid_reg <= _T_161;
    line_424_valid_reg <= inc_12;
    line_425_valid_reg <= _T_10;
    line_426_valid_reg <= _T_167;
    line_427_valid_reg <= _T_10;
    line_428_valid_reg <= _T_173;
    line_429_valid_reg <= inc_13;
    line_430_valid_reg <= _T_10;
    line_431_valid_reg <= _T_179;
    line_432_valid_reg <= _T_10;
    line_433_valid_reg <= _T_185;
    line_434_valid_reg <= inc_14;
    line_435_valid_reg <= _T_10;
    line_436_valid_reg <= _T_191;
    line_437_valid_reg <= _T_10;
    line_438_valid_reg <= _T_197;
    line_439_valid_reg <= inc_15;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec | count_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc | idle)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_1 | count_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_1 | idle_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_2 | count_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_2 | idle_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_3 | count_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_3 | idle_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_4 | count_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_4 | idle_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_5 | count_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_5 | idle_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_6 | count_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_6 | idle_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_7 | count_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_7 | idle_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_8 | count_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_8 | idle_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_9 | count_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_9 | idle_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_10 | count_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_10 | idle_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_11 | count_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_11 | idle_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_12 | count_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_12 | idle_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_13 | count_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_13 | idle_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_14 | count_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_14 | idle_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~dec_15 | count_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~inc_15 | idle_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n"); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count_16 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  count_15 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  count_14 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  count_13 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  count_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  count_11 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  count_10 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  count_9 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  count_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  count_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  count_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  count_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  count_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  count_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  count_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  count_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  counter = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  doneAW = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_321_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_322_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_323_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_324_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_325_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_326_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_327_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_328_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_329_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_330_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_331_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_332_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_333_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_334_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_335_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_336_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_337_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_338_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_339_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_340_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_341_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_342_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_343_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_344_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_345_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_346_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_347_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_348_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_349_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_350_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_351_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_352_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_353_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_354_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_holds_d = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  b_delay = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  line_355_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_356_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_357_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_first = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_358_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_denied_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_359_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_360_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_361_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_362_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_363_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_364_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_365_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_366_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_367_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_368_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_369_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_370_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_371_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_372_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_373_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_374_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_375_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_376_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_377_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_378_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_379_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_380_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_381_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_382_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_383_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_384_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_385_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_386_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_387_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_388_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_389_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_390_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_391_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_392_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_393_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_394_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_395_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_396_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_397_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_398_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_399_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_400_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_401_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_402_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_403_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_404_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_405_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_406_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_407_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_408_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_409_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_410_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_411_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_412_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_413_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_414_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_415_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_416_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_417_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_418_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_419_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_420_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_421_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_422_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_423_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_424_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_425_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_426_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_427_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_428_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_429_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_430_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_431_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_432_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_433_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_434_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_435_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_436_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_437_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_438_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_439_valid_reg = _RAND_140[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~dec | count_1); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc | idle); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_1 | count_2); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_1 | idle_1); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_2 | count_3); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_2 | idle_2); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_3 | count_4); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_3 | idle_3); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_4 | count_5); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_4 | idle_4); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_5 | count_6); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_5 | idle_5); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_6 | count_7); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_6 | idle_6); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_7 | count_8); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_7 | idle_7); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_8 | count_9); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_8 | idle_8); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_9 | count_10); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_9 | idle_9); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_10 | count_11); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_10 | idle_10); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_11 | count_12); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_11 | idle_11); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_12 | count_13); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_12 | idle_12); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_13 | count_14); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_13 | idle_13); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_14 | count_15); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_14 | idle_14); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
    //
    if (~reset) begin
      assert(~dec_15 | count_16); // @[src/main/scala/tilelink/ToAXI4.scala 273:16]
    end
    //
    if (_T_10) begin
      assert(~inc_15 | idle_15); // @[src/main/scala/tilelink/ToAXI4.scala 274:16]
    end
  end
endmodule
module TLWidthWidget_5(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLInterconnectCoupler_7(
  input         clock,
  input         reset,
  output        auto_widget_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_widget_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_widget_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_widget_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_widget_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_widget_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_axi4yank_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_axi4yank_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_axi4yank_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_axi4yank_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_axi4yank_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_axi4yank_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_axi4yank_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_axi4yank_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_axi4yank_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_axi4yank_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_axi4yank_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_axi4yank_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_axi4yank_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_axi4yank_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_axi4yank_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_axi4yank_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_axi4yank_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_axi4yank_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_axi4yank_out_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_tl_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tl_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_tl_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_tl_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_tl_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_tl_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_tl_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  axi4yank_clock; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_reset; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_aw_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_aw_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [31:0] axi4yank_auto_in_aw_bits_addr; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_in_aw_bits_len; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [2:0] axi4yank_auto_in_aw_bits_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_in_aw_bits_burst; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_w_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_w_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [63:0] axi4yank_auto_in_w_bits_data; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_in_w_bits_strb; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_w_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_b_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_b_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_b_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_in_b_bits_resp; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_b_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_b_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_ar_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_ar_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [31:0] axi4yank_auto_in_ar_bits_addr; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_in_ar_bits_len; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [2:0] axi4yank_auto_in_ar_bits_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_in_ar_bits_burst; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_r_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_r_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_r_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [63:0] axi4yank_auto_in_r_bits_data; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_in_r_bits_resp; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_r_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_in_r_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_in_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_aw_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_aw_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_out_aw_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [31:0] axi4yank_auto_out_aw_bits_addr; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_out_aw_bits_len; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [2:0] axi4yank_auto_out_aw_bits_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_out_aw_bits_burst; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_w_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_w_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [63:0] axi4yank_auto_out_w_bits_data; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_out_w_bits_strb; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_w_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_b_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_b_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_out_b_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_ar_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_ar_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_out_ar_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [31:0] axi4yank_auto_out_ar_bits_addr; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [7:0] axi4yank_auto_out_ar_bits_len; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [2:0] axi4yank_auto_out_ar_bits_size; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_out_ar_bits_burst; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_r_ready; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_r_valid; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [3:0] axi4yank_auto_out_r_bits_id; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [63:0] axi4yank_auto_out_r_bits_data; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire [1:0] axi4yank_auto_out_r_bits_resp; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4yank_auto_out_r_bits_last; // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
  wire  axi4index_clock; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_reset; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_aw_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_aw_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [31:0] axi4index_auto_in_aw_bits_addr; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_in_aw_bits_len; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [2:0] axi4index_auto_in_aw_bits_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_in_aw_bits_burst; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_aw_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_aw_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_w_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_w_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [63:0] axi4index_auto_in_w_bits_data; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_in_w_bits_strb; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_w_bits_last; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_b_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_b_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_b_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_in_b_bits_resp; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_b_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_b_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_ar_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_ar_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [31:0] axi4index_auto_in_ar_bits_addr; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_in_ar_bits_len; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [2:0] axi4index_auto_in_ar_bits_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_in_ar_bits_burst; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_ar_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_ar_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_r_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_r_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_r_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [63:0] axi4index_auto_in_r_bits_data; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_in_r_bits_resp; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_r_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_in_r_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_in_r_bits_last; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_aw_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_aw_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_aw_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [31:0] axi4index_auto_out_aw_bits_addr; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_out_aw_bits_len; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [2:0] axi4index_auto_out_aw_bits_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_out_aw_bits_burst; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_aw_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_aw_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_w_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_w_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [63:0] axi4index_auto_out_w_bits_data; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_out_w_bits_strb; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_w_bits_last; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_b_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_b_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_b_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_b_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_b_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_ar_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_ar_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_ar_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [31:0] axi4index_auto_out_ar_bits_addr; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [7:0] axi4index_auto_out_ar_bits_len; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [2:0] axi4index_auto_out_ar_bits_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_out_ar_bits_burst; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_ar_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_ar_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_r_ready; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_r_valid; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_r_bits_id; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [63:0] axi4index_auto_out_r_bits_data; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [1:0] axi4index_auto_out_r_bits_resp; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_r_bits_echo_tl_state_size; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire [3:0] axi4index_auto_out_r_bits_echo_tl_state_source; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  axi4index_auto_out_r_bits_last; // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
  wire  tl2axi4_clock; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_reset; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_a_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_a_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_in_a_bits_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_in_a_bits_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [31:0] tl2axi4_auto_in_a_bits_address; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [7:0] tl2axi4_auto_in_a_bits_mask; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [63:0] tl2axi4_auto_in_a_bits_data; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_d_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_d_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_in_d_bits_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_in_d_bits_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_d_bits_denied; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [63:0] tl2axi4_auto_in_d_bits_data; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_aw_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_aw_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_id; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [31:0] tl2axi4_auto_out_aw_bits_addr; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [7:0] tl2axi4_auto_out_aw_bits_len; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_out_aw_bits_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [1:0] tl2axi4_auto_out_aw_bits_burst; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_echo_tl_state_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_w_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_w_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [63:0] tl2axi4_auto_out_w_bits_data; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [7:0] tl2axi4_auto_out_w_bits_strb; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_w_bits_last; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_b_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_b_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_b_bits_id; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [1:0] tl2axi4_auto_out_b_bits_resp; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_b_bits_echo_tl_state_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_b_bits_echo_tl_state_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_ar_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_ar_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_id; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [31:0] tl2axi4_auto_out_ar_bits_addr; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [7:0] tl2axi4_auto_out_ar_bits_len; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [2:0] tl2axi4_auto_out_ar_bits_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [1:0] tl2axi4_auto_out_ar_bits_burst; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_echo_tl_state_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_r_ready; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_r_valid; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_r_bits_id; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [63:0] tl2axi4_auto_out_r_bits_data; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [1:0] tl2axi4_auto_out_r_bits_resp; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_r_bits_echo_tl_state_size; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire [3:0] tl2axi4_auto_out_r_bits_echo_tl_state_source; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  tl2axi4_auto_out_r_bits_last; // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_in_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_in_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_out_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_out_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_out_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  AXI4UserYanker axi4yank ( // @[src/main/scala/amba/axi4/UserYanker.scala 122:30]
    .clock(axi4yank_clock),
    .reset(axi4yank_reset),
    .auto_in_aw_ready(axi4yank_auto_in_aw_ready),
    .auto_in_aw_valid(axi4yank_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4yank_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4yank_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4yank_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4yank_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4yank_auto_in_aw_bits_burst),
    .auto_in_aw_bits_echo_tl_state_size(axi4yank_auto_in_aw_bits_echo_tl_state_size),
    .auto_in_aw_bits_echo_tl_state_source(axi4yank_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4yank_auto_in_w_ready),
    .auto_in_w_valid(axi4yank_auto_in_w_valid),
    .auto_in_w_bits_data(axi4yank_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4yank_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4yank_auto_in_w_bits_last),
    .auto_in_b_ready(axi4yank_auto_in_b_ready),
    .auto_in_b_valid(axi4yank_auto_in_b_valid),
    .auto_in_b_bits_id(axi4yank_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4yank_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_size(axi4yank_auto_in_b_bits_echo_tl_state_size),
    .auto_in_b_bits_echo_tl_state_source(axi4yank_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4yank_auto_in_ar_ready),
    .auto_in_ar_valid(axi4yank_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4yank_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4yank_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4yank_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4yank_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4yank_auto_in_ar_bits_burst),
    .auto_in_ar_bits_echo_tl_state_size(axi4yank_auto_in_ar_bits_echo_tl_state_size),
    .auto_in_ar_bits_echo_tl_state_source(axi4yank_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4yank_auto_in_r_ready),
    .auto_in_r_valid(axi4yank_auto_in_r_valid),
    .auto_in_r_bits_id(axi4yank_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4yank_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4yank_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_size(axi4yank_auto_in_r_bits_echo_tl_state_size),
    .auto_in_r_bits_echo_tl_state_source(axi4yank_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4yank_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4yank_auto_out_aw_ready),
    .auto_out_aw_valid(axi4yank_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4yank_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4yank_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4yank_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4yank_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4yank_auto_out_aw_bits_burst),
    .auto_out_w_ready(axi4yank_auto_out_w_ready),
    .auto_out_w_valid(axi4yank_auto_out_w_valid),
    .auto_out_w_bits_data(axi4yank_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4yank_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4yank_auto_out_w_bits_last),
    .auto_out_b_ready(axi4yank_auto_out_b_ready),
    .auto_out_b_valid(axi4yank_auto_out_b_valid),
    .auto_out_b_bits_id(axi4yank_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4yank_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4yank_auto_out_ar_ready),
    .auto_out_ar_valid(axi4yank_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4yank_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4yank_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4yank_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4yank_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4yank_auto_out_ar_bits_burst),
    .auto_out_r_ready(axi4yank_auto_out_r_ready),
    .auto_out_r_valid(axi4yank_auto_out_r_valid),
    .auto_out_r_bits_id(axi4yank_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4yank_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4yank_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4yank_auto_out_r_bits_last)
  );
  AXI4IdIndexer axi4index ( // @[src/main/scala/amba/axi4/IdIndexer.scala 104:31]
    .clock(axi4index_clock),
    .reset(axi4index_reset),
    .auto_in_aw_ready(axi4index_auto_in_aw_ready),
    .auto_in_aw_valid(axi4index_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4index_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4index_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4index_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4index_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4index_auto_in_aw_bits_burst),
    .auto_in_aw_bits_echo_tl_state_size(axi4index_auto_in_aw_bits_echo_tl_state_size),
    .auto_in_aw_bits_echo_tl_state_source(axi4index_auto_in_aw_bits_echo_tl_state_source),
    .auto_in_w_ready(axi4index_auto_in_w_ready),
    .auto_in_w_valid(axi4index_auto_in_w_valid),
    .auto_in_w_bits_data(axi4index_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4index_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4index_auto_in_w_bits_last),
    .auto_in_b_ready(axi4index_auto_in_b_ready),
    .auto_in_b_valid(axi4index_auto_in_b_valid),
    .auto_in_b_bits_id(axi4index_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4index_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_tl_state_size(axi4index_auto_in_b_bits_echo_tl_state_size),
    .auto_in_b_bits_echo_tl_state_source(axi4index_auto_in_b_bits_echo_tl_state_source),
    .auto_in_ar_ready(axi4index_auto_in_ar_ready),
    .auto_in_ar_valid(axi4index_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4index_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4index_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4index_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4index_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4index_auto_in_ar_bits_burst),
    .auto_in_ar_bits_echo_tl_state_size(axi4index_auto_in_ar_bits_echo_tl_state_size),
    .auto_in_ar_bits_echo_tl_state_source(axi4index_auto_in_ar_bits_echo_tl_state_source),
    .auto_in_r_ready(axi4index_auto_in_r_ready),
    .auto_in_r_valid(axi4index_auto_in_r_valid),
    .auto_in_r_bits_id(axi4index_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4index_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4index_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_tl_state_size(axi4index_auto_in_r_bits_echo_tl_state_size),
    .auto_in_r_bits_echo_tl_state_source(axi4index_auto_in_r_bits_echo_tl_state_source),
    .auto_in_r_bits_last(axi4index_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4index_auto_out_aw_ready),
    .auto_out_aw_valid(axi4index_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4index_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4index_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4index_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4index_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4index_auto_out_aw_bits_burst),
    .auto_out_aw_bits_echo_tl_state_size(axi4index_auto_out_aw_bits_echo_tl_state_size),
    .auto_out_aw_bits_echo_tl_state_source(axi4index_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(axi4index_auto_out_w_ready),
    .auto_out_w_valid(axi4index_auto_out_w_valid),
    .auto_out_w_bits_data(axi4index_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4index_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4index_auto_out_w_bits_last),
    .auto_out_b_ready(axi4index_auto_out_b_ready),
    .auto_out_b_valid(axi4index_auto_out_b_valid),
    .auto_out_b_bits_id(axi4index_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4index_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_size(axi4index_auto_out_b_bits_echo_tl_state_size),
    .auto_out_b_bits_echo_tl_state_source(axi4index_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(axi4index_auto_out_ar_ready),
    .auto_out_ar_valid(axi4index_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4index_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4index_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4index_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4index_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4index_auto_out_ar_bits_burst),
    .auto_out_ar_bits_echo_tl_state_size(axi4index_auto_out_ar_bits_echo_tl_state_size),
    .auto_out_ar_bits_echo_tl_state_source(axi4index_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(axi4index_auto_out_r_ready),
    .auto_out_r_valid(axi4index_auto_out_r_valid),
    .auto_out_r_bits_id(axi4index_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4index_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4index_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_size(axi4index_auto_out_r_bits_echo_tl_state_size),
    .auto_out_r_bits_echo_tl_state_source(axi4index_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(axi4index_auto_out_r_bits_last)
  );
  TLToAXI4 tl2axi4 ( // @[src/main/scala/tilelink/ToAXI4.scala 294:29]
    .clock(tl2axi4_clock),
    .reset(tl2axi4_reset),
    .auto_in_a_ready(tl2axi4_auto_in_a_ready),
    .auto_in_a_valid(tl2axi4_auto_in_a_valid),
    .auto_in_a_bits_opcode(tl2axi4_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(tl2axi4_auto_in_a_bits_size),
    .auto_in_a_bits_source(tl2axi4_auto_in_a_bits_source),
    .auto_in_a_bits_address(tl2axi4_auto_in_a_bits_address),
    .auto_in_a_bits_mask(tl2axi4_auto_in_a_bits_mask),
    .auto_in_a_bits_data(tl2axi4_auto_in_a_bits_data),
    .auto_in_d_ready(tl2axi4_auto_in_d_ready),
    .auto_in_d_valid(tl2axi4_auto_in_d_valid),
    .auto_in_d_bits_opcode(tl2axi4_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(tl2axi4_auto_in_d_bits_size),
    .auto_in_d_bits_source(tl2axi4_auto_in_d_bits_source),
    .auto_in_d_bits_denied(tl2axi4_auto_in_d_bits_denied),
    .auto_in_d_bits_data(tl2axi4_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(tl2axi4_auto_in_d_bits_corrupt),
    .auto_out_aw_ready(tl2axi4_auto_out_aw_ready),
    .auto_out_aw_valid(tl2axi4_auto_out_aw_valid),
    .auto_out_aw_bits_id(tl2axi4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(tl2axi4_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(tl2axi4_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(tl2axi4_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(tl2axi4_auto_out_aw_bits_burst),
    .auto_out_aw_bits_echo_tl_state_size(tl2axi4_auto_out_aw_bits_echo_tl_state_size),
    .auto_out_aw_bits_echo_tl_state_source(tl2axi4_auto_out_aw_bits_echo_tl_state_source),
    .auto_out_w_ready(tl2axi4_auto_out_w_ready),
    .auto_out_w_valid(tl2axi4_auto_out_w_valid),
    .auto_out_w_bits_data(tl2axi4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(tl2axi4_auto_out_w_bits_strb),
    .auto_out_w_bits_last(tl2axi4_auto_out_w_bits_last),
    .auto_out_b_ready(tl2axi4_auto_out_b_ready),
    .auto_out_b_valid(tl2axi4_auto_out_b_valid),
    .auto_out_b_bits_id(tl2axi4_auto_out_b_bits_id),
    .auto_out_b_bits_resp(tl2axi4_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_tl_state_size(tl2axi4_auto_out_b_bits_echo_tl_state_size),
    .auto_out_b_bits_echo_tl_state_source(tl2axi4_auto_out_b_bits_echo_tl_state_source),
    .auto_out_ar_ready(tl2axi4_auto_out_ar_ready),
    .auto_out_ar_valid(tl2axi4_auto_out_ar_valid),
    .auto_out_ar_bits_id(tl2axi4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(tl2axi4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(tl2axi4_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(tl2axi4_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(tl2axi4_auto_out_ar_bits_burst),
    .auto_out_ar_bits_echo_tl_state_size(tl2axi4_auto_out_ar_bits_echo_tl_state_size),
    .auto_out_ar_bits_echo_tl_state_source(tl2axi4_auto_out_ar_bits_echo_tl_state_source),
    .auto_out_r_ready(tl2axi4_auto_out_r_ready),
    .auto_out_r_valid(tl2axi4_auto_out_r_valid),
    .auto_out_r_bits_id(tl2axi4_auto_out_r_bits_id),
    .auto_out_r_bits_data(tl2axi4_auto_out_r_bits_data),
    .auto_out_r_bits_resp(tl2axi4_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_tl_state_size(tl2axi4_auto_out_r_bits_echo_tl_state_size),
    .auto_out_r_bits_echo_tl_state_source(tl2axi4_auto_out_r_bits_echo_tl_state_source),
    .auto_out_r_bits_last(tl2axi4_auto_out_r_bits_last)
  );
  TLWidthWidget_5 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
  );
  assign auto_widget_in_a_ready = widget_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_valid = widget_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_axi4yank_out_aw_valid = axi4yank_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_aw_bits_id = axi4yank_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_aw_bits_addr = axi4yank_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_aw_bits_len = axi4yank_auto_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_aw_bits_size = axi4yank_auto_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_aw_bits_burst = axi4yank_auto_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_w_valid = axi4yank_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_w_bits_data = axi4yank_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_w_bits_strb = axi4yank_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_w_bits_last = axi4yank_auto_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_b_ready = axi4yank_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_valid = axi4yank_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_bits_id = axi4yank_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_bits_addr = axi4yank_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_bits_len = axi4yank_auto_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_bits_size = axi4yank_auto_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_ar_bits_burst = axi4yank_auto_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_axi4yank_out_r_ready = axi4yank_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_a_ready = auto_tl_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_valid = auto_tl_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_opcode = auto_tl_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_size = auto_tl_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_source = auto_tl_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_denied = auto_tl_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_data = auto_tl_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_in_d_bits_corrupt = auto_tl_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tl_out_a_valid = auto_tl_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_opcode = auto_tl_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_size = auto_tl_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_source = auto_tl_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_address = auto_tl_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_mask = auto_tl_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_a_bits_data = auto_tl_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_tl_out_d_ready = auto_tl_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign axi4yank_clock = clock;
  assign axi4yank_reset = reset;
  assign axi4yank_auto_in_aw_valid = axi4index_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_id = axi4index_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_addr = axi4index_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_len = axi4index_auto_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_size = axi4index_auto_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_burst = axi4index_auto_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_echo_tl_state_size = axi4index_auto_out_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_aw_bits_echo_tl_state_source = axi4index_auto_out_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_w_valid = axi4index_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_w_bits_data = axi4index_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_w_bits_strb = axi4index_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_w_bits_last = axi4index_auto_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_b_ready = axi4index_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_valid = axi4index_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_id = axi4index_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_addr = axi4index_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_len = axi4index_auto_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_size = axi4index_auto_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_burst = axi4index_auto_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_echo_tl_state_size = axi4index_auto_out_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_ar_bits_echo_tl_state_source = axi4index_auto_out_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_in_r_ready = axi4index_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4yank_auto_out_aw_ready = auto_axi4yank_out_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_w_ready = auto_axi4yank_out_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_b_valid = auto_axi4yank_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_b_bits_id = auto_axi4yank_out_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_b_bits_resp = auto_axi4yank_out_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_ar_ready = auto_axi4yank_out_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_r_valid = auto_axi4yank_out_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_r_bits_id = auto_axi4yank_out_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_r_bits_data = auto_axi4yank_out_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_r_bits_resp = auto_axi4yank_out_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4yank_auto_out_r_bits_last = auto_axi4yank_out_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign axi4index_clock = clock;
  assign axi4index_reset = reset;
  assign axi4index_auto_in_aw_valid = tl2axi4_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_id = tl2axi4_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_addr = tl2axi4_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_len = tl2axi4_auto_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_size = tl2axi4_auto_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_burst = tl2axi4_auto_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_echo_tl_state_size = tl2axi4_auto_out_aw_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_aw_bits_echo_tl_state_source = tl2axi4_auto_out_aw_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_w_valid = tl2axi4_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_w_bits_data = tl2axi4_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_w_bits_strb = tl2axi4_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_w_bits_last = tl2axi4_auto_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_b_ready = tl2axi4_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_valid = tl2axi4_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_id = tl2axi4_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_addr = tl2axi4_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_len = tl2axi4_auto_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_size = tl2axi4_auto_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_burst = tl2axi4_auto_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_echo_tl_state_size = tl2axi4_auto_out_ar_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_ar_bits_echo_tl_state_source = tl2axi4_auto_out_ar_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_in_r_ready = tl2axi4_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_aw_ready = axi4yank_auto_in_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_w_ready = axi4yank_auto_in_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_b_valid = axi4yank_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_b_bits_id = axi4yank_auto_in_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_b_bits_resp = axi4yank_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_b_bits_echo_tl_state_size = axi4yank_auto_in_b_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_b_bits_echo_tl_state_source = axi4yank_auto_in_b_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_ar_ready = axi4yank_auto_in_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_valid = axi4yank_auto_in_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_id = axi4yank_auto_in_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_data = axi4yank_auto_in_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_resp = axi4yank_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_echo_tl_state_size = axi4yank_auto_in_r_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_echo_tl_state_source = axi4yank_auto_in_r_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4index_auto_out_r_bits_last = axi4yank_auto_in_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_clock = clock;
  assign tl2axi4_reset = reset;
  assign tl2axi4_auto_in_a_valid = widget_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_size = widget_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_source = widget_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_address = widget_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_mask = widget_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_a_bits_data = widget_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_in_d_ready = widget_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_aw_ready = axi4index_auto_in_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_w_ready = axi4index_auto_in_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_b_valid = axi4index_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_b_bits_id = axi4index_auto_in_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_b_bits_resp = axi4index_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_b_bits_echo_tl_state_size = axi4index_auto_in_b_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_b_bits_echo_tl_state_source = axi4index_auto_in_b_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_ar_ready = axi4index_auto_in_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_valid = axi4index_auto_in_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_id = axi4index_auto_in_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_data = axi4index_auto_in_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_resp = axi4index_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_echo_tl_state_size = axi4index_auto_in_r_bits_echo_tl_state_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_echo_tl_state_source = axi4index_auto_in_r_bits_echo_tl_state_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tl2axi4_auto_out_r_bits_last = axi4index_auto_in_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_opcode = auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_data = auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_d_ready = auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_out_a_ready = tl2axi4_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_valid = tl2axi4_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_opcode = tl2axi4_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_size = tl2axi4_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_source = tl2axi4_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_denied = tl2axi4_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_data = tl2axi4_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_corrupt = tl2axi4_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module MemoryBus(
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_bus_xing_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_bus_xing_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_bus_xing_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_bus_xing_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_bus_xing_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_bus_xing_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_mbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_mbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  subsystem_mbus_xbar_clock; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_reset; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_a_ready; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_a_valid; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_in_a_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_in_a_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [3:0] subsystem_mbus_xbar_auto_in_a_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [31:0] subsystem_mbus_xbar_auto_in_a_bits_address; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [7:0] subsystem_mbus_xbar_auto_in_a_bits_mask; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [63:0] subsystem_mbus_xbar_auto_in_a_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_d_ready; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_d_valid; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_in_d_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_in_d_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [3:0] subsystem_mbus_xbar_auto_in_d_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_d_bits_denied; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [63:0] subsystem_mbus_xbar_auto_in_d_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_a_ready; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_a_valid; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_out_a_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_out_a_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [3:0] subsystem_mbus_xbar_auto_out_a_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [31:0] subsystem_mbus_xbar_auto_out_a_bits_address; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [7:0] subsystem_mbus_xbar_auto_out_a_bits_mask; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [63:0] subsystem_mbus_xbar_auto_out_a_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_d_ready; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_d_valid; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_out_d_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [2:0] subsystem_mbus_xbar_auto_out_d_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [3:0] subsystem_mbus_xbar_auto_out_d_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_d_bits_denied; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire [63:0] subsystem_mbus_xbar_auto_out_d_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  subsystem_mbus_xbar_auto_out_d_bits_corrupt; // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
  wire  fixer_clock; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_reset; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_a_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [3:0] fixer_auto_in_a_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_in_a_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [7:0] fixer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_in_a_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_in_d_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [3:0] fixer_auto_in_d_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_in_d_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_a_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_a_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_a_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [3:0] fixer_auto_out_a_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [31:0] fixer_auto_out_a_bits_address; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [7:0] fixer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_out_a_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_ready; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_valid; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [2:0] fixer_auto_out_d_bits_size; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [3:0] fixer_auto_out_d_bits_source; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_bits_denied; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire [63:0] fixer_auto_out_d_bits_data; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  fixer_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
  wire  picker_clock; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_reset; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_a_ready; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_a_valid; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_in_a_bits_size; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [3:0] picker_auto_in_a_bits_source; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [31:0] picker_auto_in_a_bits_address; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [7:0] picker_auto_in_a_bits_mask; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [63:0] picker_auto_in_a_bits_data; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_d_ready; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_d_valid; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_in_d_bits_size; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [3:0] picker_auto_in_d_bits_source; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_d_bits_denied; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [63:0] picker_auto_in_d_bits_data; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_a_ready; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_a_valid; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_out_a_bits_size; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [3:0] picker_auto_out_a_bits_source; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [31:0] picker_auto_out_a_bits_address; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [7:0] picker_auto_out_a_bits_mask; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [63:0] picker_auto_out_a_bits_data; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_d_ready; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_d_valid; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [2:0] picker_auto_out_d_bits_size; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [3:0] picker_auto_out_d_bits_source; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_d_bits_denied; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire [63:0] picker_auto_out_d_bits_data; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  picker_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [3:0] buffer_auto_in_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [3:0] buffer_auto_out_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  xbar_clock; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_reset; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_a_ready; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_in_a_bits_size; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [3:0] xbar_auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [31:0] xbar_auto_in_a_bits_address; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [63:0] xbar_auto_in_a_bits_data; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_d_ready; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_d_valid; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_in_d_bits_size; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [3:0] xbar_auto_in_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [63:0] xbar_auto_in_d_bits_data; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_a_ready; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_a_valid; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_out_a_bits_size; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [3:0] xbar_auto_out_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [31:0] xbar_auto_out_a_bits_address; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [7:0] xbar_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [63:0] xbar_auto_out_a_bits_data; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_d_ready; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [2:0] xbar_auto_out_d_bits_size; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [3:0] xbar_auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_d_bits_denied; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire [63:0] xbar_auto_out_d_bits_data; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  xbar_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/Xbar.scala 343:26]
  wire  coupler_to_memory_controller_port_named_axi4_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [1:0] coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  ClockGroupAggregator_4 subsystem_mbus_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_mbus_0_clock(subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock),
    .auto_in_member_subsystem_mbus_0_reset(subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset),
    .auto_out_member_subsystem_mbus_0_clock(subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock),
    .auto_out_member_subsystem_mbus_0_reset(subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset)
  );
  ClockGroup_4 clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_mbus_0_clock(clockGroup_auto_in_member_subsystem_mbus_0_clock),
    .auto_in_member_subsystem_mbus_0_reset(clockGroup_auto_in_member_subsystem_mbus_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast_4 fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_clock(fixedClockNode_auto_out_clock),
    .auto_out_reset(fixedClockNode_auto_out_reset)
  );
  BundleBridgeNexus_4 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLXbar_6 subsystem_mbus_xbar ( // @[src/main/scala/subsystem/MemoryBus.scala 42:32]
    .clock(subsystem_mbus_xbar_clock),
    .reset(subsystem_mbus_xbar_reset),
    .auto_in_a_ready(subsystem_mbus_xbar_auto_in_a_ready),
    .auto_in_a_valid(subsystem_mbus_xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(subsystem_mbus_xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(subsystem_mbus_xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(subsystem_mbus_xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(subsystem_mbus_xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(subsystem_mbus_xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(subsystem_mbus_xbar_auto_in_a_bits_data),
    .auto_in_d_ready(subsystem_mbus_xbar_auto_in_d_ready),
    .auto_in_d_valid(subsystem_mbus_xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(subsystem_mbus_xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(subsystem_mbus_xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(subsystem_mbus_xbar_auto_in_d_bits_source),
    .auto_in_d_bits_denied(subsystem_mbus_xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(subsystem_mbus_xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(subsystem_mbus_xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(subsystem_mbus_xbar_auto_out_a_ready),
    .auto_out_a_valid(subsystem_mbus_xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(subsystem_mbus_xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(subsystem_mbus_xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(subsystem_mbus_xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(subsystem_mbus_xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(subsystem_mbus_xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(subsystem_mbus_xbar_auto_out_a_bits_data),
    .auto_out_d_ready(subsystem_mbus_xbar_auto_out_d_ready),
    .auto_out_d_valid(subsystem_mbus_xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(subsystem_mbus_xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(subsystem_mbus_xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(subsystem_mbus_xbar_auto_out_d_bits_source),
    .auto_out_d_bits_denied(subsystem_mbus_xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(subsystem_mbus_xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(subsystem_mbus_xbar_auto_out_d_bits_corrupt)
  );
  TLFIFOFixer_3 fixer ( // @[src/main/scala/tilelink/FIFOFixer.scala 146:27]
    .clock(fixer_clock),
    .reset(fixer_reset),
    .auto_in_a_ready(fixer_auto_in_a_ready),
    .auto_in_a_valid(fixer_auto_in_a_valid),
    .auto_in_a_bits_opcode(fixer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(fixer_auto_in_a_bits_size),
    .auto_in_a_bits_source(fixer_auto_in_a_bits_source),
    .auto_in_a_bits_address(fixer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fixer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fixer_auto_in_a_bits_data),
    .auto_in_d_ready(fixer_auto_in_d_ready),
    .auto_in_d_valid(fixer_auto_in_d_valid),
    .auto_in_d_bits_opcode(fixer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(fixer_auto_in_d_bits_size),
    .auto_in_d_bits_source(fixer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(fixer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fixer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fixer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fixer_auto_out_a_ready),
    .auto_out_a_valid(fixer_auto_out_a_valid),
    .auto_out_a_bits_opcode(fixer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(fixer_auto_out_a_bits_size),
    .auto_out_a_bits_source(fixer_auto_out_a_bits_source),
    .auto_out_a_bits_address(fixer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fixer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fixer_auto_out_a_bits_data),
    .auto_out_d_ready(fixer_auto_out_d_ready),
    .auto_out_d_valid(fixer_auto_out_d_valid),
    .auto_out_d_bits_opcode(fixer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(fixer_auto_out_d_bits_size),
    .auto_out_d_bits_source(fixer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(fixer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fixer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fixer_auto_out_d_bits_corrupt)
  );
  ProbePicker picker ( // @[src/main/scala/tilelink/ProbePicker.scala 66:28]
    .clock(picker_clock),
    .reset(picker_reset),
    .auto_in_a_ready(picker_auto_in_a_ready),
    .auto_in_a_valid(picker_auto_in_a_valid),
    .auto_in_a_bits_opcode(picker_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(picker_auto_in_a_bits_size),
    .auto_in_a_bits_source(picker_auto_in_a_bits_source),
    .auto_in_a_bits_address(picker_auto_in_a_bits_address),
    .auto_in_a_bits_mask(picker_auto_in_a_bits_mask),
    .auto_in_a_bits_data(picker_auto_in_a_bits_data),
    .auto_in_d_ready(picker_auto_in_d_ready),
    .auto_in_d_valid(picker_auto_in_d_valid),
    .auto_in_d_bits_opcode(picker_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(picker_auto_in_d_bits_size),
    .auto_in_d_bits_source(picker_auto_in_d_bits_source),
    .auto_in_d_bits_denied(picker_auto_in_d_bits_denied),
    .auto_in_d_bits_data(picker_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(picker_auto_in_d_bits_corrupt),
    .auto_out_a_ready(picker_auto_out_a_ready),
    .auto_out_a_valid(picker_auto_out_a_valid),
    .auto_out_a_bits_opcode(picker_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(picker_auto_out_a_bits_size),
    .auto_out_a_bits_source(picker_auto_out_a_bits_source),
    .auto_out_a_bits_address(picker_auto_out_a_bits_address),
    .auto_out_a_bits_mask(picker_auto_out_a_bits_mask),
    .auto_out_a_bits_data(picker_auto_out_a_bits_data),
    .auto_out_d_ready(picker_auto_out_d_ready),
    .auto_out_d_valid(picker_auto_out_d_valid),
    .auto_out_d_bits_opcode(picker_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(picker_auto_out_d_bits_size),
    .auto_out_d_bits_source(picker_auto_out_d_bits_source),
    .auto_out_d_bits_denied(picker_auto_out_d_bits_denied),
    .auto_out_d_bits_data(picker_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(picker_auto_out_d_bits_corrupt)
  );
  TLBuffer_5 buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt)
  );
  TLXbar_7 xbar ( // @[src/main/scala/tilelink/Xbar.scala 343:26]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLInterconnectCoupler_7 coupler_to_memory_controller_port_named_axi4 ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_memory_controller_port_named_axi4_clock),
    .reset(coupler_to_memory_controller_port_named_axi4_reset),
    .auto_widget_in_a_ready(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready),
    .auto_widget_in_a_valid(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_valid),
    .auto_widget_in_a_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_opcode),
    .auto_widget_in_a_bits_size(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_size),
    .auto_widget_in_a_bits_source(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_source),
    .auto_widget_in_a_bits_address(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_address),
    .auto_widget_in_a_bits_mask(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_mask),
    .auto_widget_in_a_bits_data(coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_data),
    .auto_widget_in_d_ready(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_ready),
    .auto_widget_in_d_valid(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid),
    .auto_widget_in_d_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode),
    .auto_widget_in_d_bits_size(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size),
    .auto_widget_in_d_bits_source(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source),
    .auto_widget_in_d_bits_denied(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied),
    .auto_widget_in_d_bits_data(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data),
    .auto_widget_in_d_bits_corrupt(coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt),
    .auto_axi4yank_out_aw_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready),
    .auto_axi4yank_out_aw_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid),
    .auto_axi4yank_out_aw_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id),
    .auto_axi4yank_out_aw_bits_addr(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr),
    .auto_axi4yank_out_aw_bits_len(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len),
    .auto_axi4yank_out_aw_bits_size(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size),
    .auto_axi4yank_out_aw_bits_burst(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst),
    .auto_axi4yank_out_w_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready),
    .auto_axi4yank_out_w_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid),
    .auto_axi4yank_out_w_bits_data(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data),
    .auto_axi4yank_out_w_bits_strb(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb),
    .auto_axi4yank_out_w_bits_last(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last),
    .auto_axi4yank_out_b_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready),
    .auto_axi4yank_out_b_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid),
    .auto_axi4yank_out_b_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id),
    .auto_axi4yank_out_b_bits_resp(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp),
    .auto_axi4yank_out_ar_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready),
    .auto_axi4yank_out_ar_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid),
    .auto_axi4yank_out_ar_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id),
    .auto_axi4yank_out_ar_bits_addr(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr),
    .auto_axi4yank_out_ar_bits_len(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len),
    .auto_axi4yank_out_ar_bits_size(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size),
    .auto_axi4yank_out_ar_bits_burst(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst),
    .auto_axi4yank_out_r_ready(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready),
    .auto_axi4yank_out_r_valid(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid),
    .auto_axi4yank_out_r_bits_id(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id),
    .auto_axi4yank_out_r_bits_data(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data),
    .auto_axi4yank_out_r_bits_resp(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp),
    .auto_axi4yank_out_r_bits_last(coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last),
    .auto_tl_in_a_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),
    .auto_tl_in_a_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid),
    .auto_tl_in_a_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode),
    .auto_tl_in_a_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size),
    .auto_tl_in_a_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source),
    .auto_tl_in_a_bits_address(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address),
    .auto_tl_in_a_bits_mask(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask),
    .auto_tl_in_a_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data),
    .auto_tl_in_d_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready),
    .auto_tl_in_d_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),
    .auto_tl_in_d_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),
    .auto_tl_in_d_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),
    .auto_tl_in_d_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),
    .auto_tl_in_d_bits_denied(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),
    .auto_tl_in_d_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data),
    .auto_tl_in_d_bits_corrupt(coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt),
    .auto_tl_out_a_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_ready),
    .auto_tl_out_a_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid),
    .auto_tl_out_a_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode),
    .auto_tl_out_a_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size),
    .auto_tl_out_a_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source),
    .auto_tl_out_a_bits_address(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address),
    .auto_tl_out_a_bits_mask(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask),
    .auto_tl_out_a_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data),
    .auto_tl_out_d_ready(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready),
    .auto_tl_out_d_valid(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_valid),
    .auto_tl_out_d_bits_opcode(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_opcode),
    .auto_tl_out_d_bits_size(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_size),
    .auto_tl_out_d_bits_source(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_source),
    .auto_tl_out_d_bits_denied(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_denied),
    .auto_tl_out_d_bits_data(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_data),
    .auto_tl_out_d_bits_corrupt(coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_corrupt)
  );
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready =
    coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_bus_xing_in_a_ready = buffer_auto_in_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_valid = buffer_auto_in_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_size = buffer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_source = buffer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_denied = buffer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_data = buffer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign auto_bus_xing_in_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_clock =
    auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_mbus_clock_groups_auto_in_member_subsystem_mbus_0_reset =
    auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_mbus_0_clock =
    subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_mbus_0_reset =
    subsystem_mbus_clock_groups_auto_out_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_valid = fixer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_opcode = fixer_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_size = fixer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_source = fixer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_address = fixer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_mask = fixer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_a_bits_data = fixer_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_in_d_ready = fixer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_xbar_auto_out_a_ready = picker_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_valid = picker_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_opcode = picker_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_size = picker_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_source = picker_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_denied = picker_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_data = picker_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_xbar_auto_out_d_bits_corrupt = picker_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixer_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_valid = buffer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_in_d_ready = buffer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_a_ready = subsystem_mbus_xbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_valid = subsystem_mbus_xbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_opcode = subsystem_mbus_xbar_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_size = subsystem_mbus_xbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_source = subsystem_mbus_xbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_denied = subsystem_mbus_xbar_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_data = subsystem_mbus_xbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fixer_auto_out_d_bits_corrupt = subsystem_mbus_xbar_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign picker_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign picker_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign picker_auto_in_a_valid = subsystem_mbus_xbar_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_opcode = subsystem_mbus_xbar_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_size = subsystem_mbus_xbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_source = subsystem_mbus_xbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_address = subsystem_mbus_xbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_mask = subsystem_mbus_xbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_a_bits_data = subsystem_mbus_xbar_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_in_d_ready = subsystem_mbus_xbar_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_a_ready = coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_valid = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_opcode = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_size = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_source = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_denied = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_data = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign picker_auto_out_d_bits_corrupt = coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_valid = auto_bus_xing_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_opcode = auto_bus_xing_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_size = auto_bus_xing_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_source = auto_bus_xing_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_address = auto_bus_xing_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_mask = auto_bus_xing_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_bits_data = auto_bus_xing_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_d_ready = auto_bus_xing_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_out_a_ready = fixer_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_valid = fixer_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_opcode = fixer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_size = fixer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_source = fixer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_denied = fixer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_data = fixer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_d_bits_corrupt = fixer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_valid = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_opcode = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_size = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_source = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_address = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_mask = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_a_bits_data = coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_in_d_ready = coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign xbar_auto_out_a_ready = coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_valid = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_opcode = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_size = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_source = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_denied = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_data = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_auto_out_d_bits_corrupt = coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_valid = xbar_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_size = xbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_source = xbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_address = xbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_bits_data = xbar_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_ready = xbar_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_aw_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_w_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_valid =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_id =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_b_bits_resp =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_ar_ready =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_valid =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_id =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_data =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_resp =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_axi4yank_out_r_bits_last =
    auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_valid = picker_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_opcode = picker_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_size = picker_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_source = picker_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_address = picker_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_mask = picker_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_bits_data = picker_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_ready = picker_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_ready = xbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_valid = xbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_size = xbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_source = xbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_data = xbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module ClockGroupAggregator_5(
  input   auto_in_member_subsystem_l2_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_l2_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_l2_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_1_member_subsystem_mbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_0_member_subsystem_l2_0_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_1_member_subsystem_mbus_0_clock = auto_in_member_subsystem_l2_1_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_1_member_subsystem_mbus_0_reset = auto_in_member_subsystem_l2_1_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_l2_0_clock = auto_in_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_0_member_subsystem_l2_0_reset = auto_in_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ClockGroup_5(
  input   auto_in_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_member_subsystem_l2_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_5(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_5(
  input   clock,
  input   reset
);
endmodule
module BroadcastFilter(
  input         clock,
  input         reset,
  output        io_request_ready, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input         io_request_valid, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input  [1:0]  io_request_bits_mshr, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input  [31:0] io_request_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input         io_request_bits_allocOH, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input         io_request_bits_needT, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  input         io_response_ready, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  output        io_response_valid, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  output [1:0]  io_response_bits_mshr, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  output [31:0] io_response_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  output        io_response_bits_allocOH, // @[src/main/scala/tilelink/Broadcast.scala 356:14]
  output        io_response_bits_needT // @[src/main/scala/tilelink/Broadcast.scala 356:14]
);
  assign io_request_ready = io_response_ready; // @[src/main/scala/tilelink/Broadcast.scala 362:20]
  assign io_response_valid = io_request_valid; // @[src/main/scala/tilelink/Broadcast.scala 363:21]
  assign io_response_bits_mshr = io_request_bits_mshr; // @[src/main/scala/tilelink/Broadcast.scala 365:28]
  assign io_response_bits_address = io_request_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 366:28]
  assign io_response_bits_allocOH = io_request_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 368:28]
  assign io_response_bits_needT = io_request_bits_needT; // @[src/main/scala/tilelink/Broadcast.scala 367:28]
endmodule
module Queue_36(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_mask [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_440_clock;
  wire  line_440_reset;
  wire  line_440_valid;
  reg  line_440_valid_reg;
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_441_clock;
  wire  line_441_reset;
  wire  line_441_valid;
  reg  line_441_valid_reg;
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_442_clock;
  wire  line_442_reset;
  wire  line_442_valid;
  reg  line_442_valid_reg;
  GEN_w1_line #(.COVER_INDEX(440)) line_440 (
    .clock(line_440_clock),
    .reset(line_440_reset),
    .valid(line_440_valid)
  );
  GEN_w1_line #(.COVER_INDEX(441)) line_441 (
    .clock(line_441_clock),
    .reset(line_441_reset),
    .valid(line_441_valid)
  );
  GEN_w1_line #(.COVER_INDEX(442)) line_442 (
    .clock(line_442_clock),
    .reset(line_442_reset),
    .valid(line_442_valid)
  );
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_440_clock = clock;
  assign line_440_reset = reset;
  assign line_440_valid = do_enq ^ line_440_valid_reg;
  assign line_441_clock = clock;
  assign line_441_reset = reset;
  assign line_441_valid = do_deq ^ line_441_valid_reg;
  assign line_442_clock = clock;
  assign line_442_reset = reset;
  assign line_442_valid = _T ^ line_442_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_440_valid_reg <= do_enq;
    line_441_valid_reg <= do_deq;
    line_442_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_440_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_441_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_442_valid_reg = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker(
  input         clock,
  input         reset,
  input         io_in_a_first, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_in_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_in_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [1:0]  io_in_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [31:0] io_in_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [7:0]  io_in_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [63:0] io_in_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_out_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_out_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [3:0]  io_out_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [31:0] io_out_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [7:0]  io_out_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [63:0] io_out_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_bits_count, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probenack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probedack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probesack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_d_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_e_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [1:0]  io_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [26:0] io_line, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_idle, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_need_d // @[src/main/scala/tilelink/Broadcast.scala 401:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  reg  got_e; // @[src/main/scala/tilelink/Broadcast.scala 424:24]
  reg  sent_d; // @[src/main/scala/tilelink/Broadcast.scala 425:24]
  reg  shared; // @[src/main/scala/tilelink/Broadcast.scala 426:20]
  reg [2:0] opcode; // @[src/main/scala/tilelink/Broadcast.scala 427:20]
  reg [2:0] size; // @[src/main/scala/tilelink/Broadcast.scala 429:20]
  reg [1:0] source; // @[src/main/scala/tilelink/Broadcast.scala 430:20]
  reg [31:0] address; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
  reg  count; // @[src/main/scala/tilelink/Broadcast.scala 434:20]
  wire  idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 438:22]
  wire  line_443_clock;
  wire  line_443_reset;
  wire  line_443_valid;
  reg  line_443_valid_reg;
  wire  _T_3 = ~reset; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_444_clock;
  wire  line_444_reset;
  wire  line_444_valid;
  reg  line_444_valid_reg;
  wire  _T_4 = ~idle; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_445_clock;
  wire  line_445_reset;
  wire  line_445_valid;
  reg  line_445_valid_reg;
  wire  _GEN_14 = _T & io_in_a_first ? 1'h0 : sent_d; // @[src/main/scala/tilelink/Broadcast.scala 438:40 440:13 425:24]
  wire  _GEN_15 = _T & io_in_a_first ? 1'h0 : shared; // @[src/main/scala/tilelink/Broadcast.scala 438:40 441:13 426:20]
  wire  _GEN_16 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[src/main/scala/tilelink/Broadcast.scala 438:40 442:13 424:24]
  wire  _GEN_22 = _T & io_in_a_first | count; // @[src/main/scala/tilelink/Broadcast.scala 438:40 450:13 434:20]
  wire  line_446_clock;
  wire  line_446_reset;
  wire  line_446_valid;
  reg  line_446_valid_reg;
  wire  _GEN_23 = io_probe_valid ? io_probe_bits_count : _GEN_22; // @[src/main/scala/tilelink/Broadcast.scala 454:25 455:13]
  wire  line_447_clock;
  wire  line_447_reset;
  wire  line_447_valid;
  reg  line_447_valid_reg;
  wire  line_448_clock;
  wire  line_448_reset;
  wire  line_448_valid;
  reg  line_448_valid_reg;
  wire  _T_8 = ~(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
  wire  line_449_clock;
  wire  line_449_reset;
  wire  line_449_valid;
  reg  line_449_valid_reg;
  wire  _GEN_25 = io_d_last | _GEN_14; // @[src/main/scala/tilelink/Broadcast.scala 459:20 461:12]
  wire  line_450_clock;
  wire  line_450_reset;
  wire  line_450_valid;
  reg  line_450_valid_reg;
  wire  line_451_clock;
  wire  line_451_reset;
  wire  line_451_valid;
  reg  line_451_valid_reg;
  wire  _T_12 = ~(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
  wire  line_452_clock;
  wire  line_452_reset;
  wire  line_452_valid;
  reg  line_452_valid_reg;
  wire  _GEN_26 = io_e_last | _GEN_16; // @[src/main/scala/tilelink/Broadcast.scala 463:20 465:11]
  wire  _T_13 = io_probenack | io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 468:22]
  wire  line_453_clock;
  wire  line_453_reset;
  wire  line_453_valid;
  reg  line_453_valid_reg;
  wire  line_454_clock;
  wire  line_454_reset;
  wire  line_454_valid;
  reg  line_454_valid_reg;
  wire  _T_17 = ~(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
  wire  line_455_clock;
  wire  line_455_reset;
  wire  line_455_valid;
  reg  line_455_valid_reg;
  wire [1:0] _count_T_1 = io_probenack & io_probedack ? 2'h2 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 470:25]
  wire [1:0] _GEN_29 = {{1'd0}, count}; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _count_T_3 = _GEN_29 - _count_T_1; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _GEN_27 = io_probenack | io_probedack ? _count_T_3 : {{1'd0}, _GEN_23}; // @[src/main/scala/tilelink/Broadcast.scala 468:39 470:11]
  wire  line_456_clock;
  wire  line_456_reset;
  wire  line_456_valid;
  reg  line_456_valid_reg;
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 486:26]
  wire  i_data_ready = o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 385:17 src/main/scala/tilelink/Broadcast.scala 483:20]
  wire  probe_done = ~count; // @[src/main/scala/tilelink/Broadcast.scala 491:26]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[src/main/scala/tilelink/Broadcast.scala 492:52]
  wire [1:0] transform = shared ? 2'h2 : 2'h3; // @[src/main/scala/tilelink/Broadcast.scala 494:22]
  wire [1:0] _io_out_a_bits_source_T = acquire ? transform : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 501:35]
  Queue_36 o_data_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(o_data_q_clock),
    .reset(o_data_q_reset),
    .io_enq_ready(o_data_q_io_enq_ready),
    .io_enq_valid(o_data_q_io_enq_valid),
    .io_enq_bits_mask(o_data_q_io_enq_bits_mask),
    .io_enq_bits_data(o_data_q_io_enq_bits_data),
    .io_deq_ready(o_data_q_io_deq_ready),
    .io_deq_valid(o_data_q_io_deq_valid),
    .io_deq_bits_mask(o_data_q_io_deq_bits_mask),
    .io_deq_bits_data(o_data_q_io_deq_bits_data)
  );
  GEN_w1_line #(.COVER_INDEX(443)) line_443 (
    .clock(line_443_clock),
    .reset(line_443_reset),
    .valid(line_443_valid)
  );
  GEN_w1_line #(.COVER_INDEX(444)) line_444 (
    .clock(line_444_clock),
    .reset(line_444_reset),
    .valid(line_444_valid)
  );
  GEN_w1_line #(.COVER_INDEX(445)) line_445 (
    .clock(line_445_clock),
    .reset(line_445_reset),
    .valid(line_445_valid)
  );
  GEN_w1_line #(.COVER_INDEX(446)) line_446 (
    .clock(line_446_clock),
    .reset(line_446_reset),
    .valid(line_446_valid)
  );
  GEN_w1_line #(.COVER_INDEX(447)) line_447 (
    .clock(line_447_clock),
    .reset(line_447_reset),
    .valid(line_447_valid)
  );
  GEN_w1_line #(.COVER_INDEX(448)) line_448 (
    .clock(line_448_clock),
    .reset(line_448_reset),
    .valid(line_448_valid)
  );
  GEN_w1_line #(.COVER_INDEX(449)) line_449 (
    .clock(line_449_clock),
    .reset(line_449_reset),
    .valid(line_449_valid)
  );
  GEN_w1_line #(.COVER_INDEX(450)) line_450 (
    .clock(line_450_clock),
    .reset(line_450_reset),
    .valid(line_450_valid)
  );
  GEN_w1_line #(.COVER_INDEX(451)) line_451 (
    .clock(line_451_clock),
    .reset(line_451_reset),
    .valid(line_451_valid)
  );
  GEN_w1_line #(.COVER_INDEX(452)) line_452 (
    .clock(line_452_clock),
    .reset(line_452_reset),
    .valid(line_452_valid)
  );
  GEN_w1_line #(.COVER_INDEX(453)) line_453 (
    .clock(line_453_clock),
    .reset(line_453_reset),
    .valid(line_453_valid)
  );
  GEN_w1_line #(.COVER_INDEX(454)) line_454 (
    .clock(line_454_clock),
    .reset(line_454_reset),
    .valid(line_454_valid)
  );
  GEN_w1_line #(.COVER_INDEX(455)) line_455 (
    .clock(line_455_clock),
    .reset(line_455_reset),
    .valid(line_455_valid)
  );
  GEN_w1_line #(.COVER_INDEX(456)) line_456 (
    .clock(line_456_clock),
    .reset(line_456_reset),
    .valid(line_456_valid)
  );
  assign line_443_clock = clock;
  assign line_443_reset = reset;
  assign line_443_valid = _T_1 ^ line_443_valid_reg;
  assign line_444_clock = clock;
  assign line_444_reset = reset;
  assign line_444_valid = _T_3 ^ line_444_valid_reg;
  assign line_445_clock = clock;
  assign line_445_reset = reset;
  assign line_445_valid = _T_4 ^ line_445_valid_reg;
  assign line_446_clock = clock;
  assign line_446_reset = reset;
  assign line_446_valid = io_probe_valid ^ line_446_valid_reg;
  assign line_447_clock = clock;
  assign line_447_reset = reset;
  assign line_447_valid = io_d_last ^ line_447_valid_reg;
  assign line_448_clock = clock;
  assign line_448_reset = reset;
  assign line_448_valid = _T_3 ^ line_448_valid_reg;
  assign line_449_clock = clock;
  assign line_449_reset = reset;
  assign line_449_valid = _T_8 ^ line_449_valid_reg;
  assign line_450_clock = clock;
  assign line_450_reset = reset;
  assign line_450_valid = io_e_last ^ line_450_valid_reg;
  assign line_451_clock = clock;
  assign line_451_reset = reset;
  assign line_451_valid = _T_3 ^ line_451_valid_reg;
  assign line_452_clock = clock;
  assign line_452_reset = reset;
  assign line_452_valid = _T_12 ^ line_452_valid_reg;
  assign line_453_clock = clock;
  assign line_453_reset = reset;
  assign line_453_valid = _T_13 ^ line_453_valid_reg;
  assign line_454_clock = clock;
  assign line_454_reset = reset;
  assign line_454_valid = _T_3 ^ line_454_valid_reg;
  assign line_455_clock = clock;
  assign line_455_reset = reset;
  assign line_455_valid = _T_17 ^ line_455_valid_reg;
  assign line_456_clock = clock;
  assign line_456_reset = reset;
  assign line_456_valid = io_probesack ^ line_456_valid_reg;
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[src/main/scala/tilelink/Broadcast.scala 486:45]
  assign io_out_a_valid = o_data_q_io_deq_valid & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 497:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[src/main/scala/tilelink/Broadcast.scala 498:31]
  assign io_out_a_bits_size = size; // @[src/main/scala/tilelink/Broadcast.scala 500:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[src/main/scala/tilelink/Broadcast.scala 501:31]
  assign io_out_a_bits_address = address; // @[src/main/scala/tilelink/Broadcast.scala 502:25]
  assign io_out_a_bits_mask = o_data_q_io_deq_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 503:25]
  assign io_out_a_bits_data = o_data_q_io_deq_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 504:25]
  assign io_source = source; // @[src/main/scala/tilelink/Broadcast.scala 479:13]
  assign io_line = address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 480:22]
  assign io_idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  assign io_need_d = ~sent_d; // @[src/main/scala/tilelink/Broadcast.scala 478:16]
  assign o_data_q_clock = clock;
  assign o_data_q_reset = reset;
  assign o_data_q_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 487:44]
  assign o_data_q_io_enq_bits_mask = io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 483:20 488:20]
  assign o_data_q_io_enq_bits_data = io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 483:20 489:20]
  assign o_data_q_io_deq_ready = io_out_a_ready & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 496:34]
  always @(posedge clock) begin
    got_e <= reset | _GEN_26; // @[src/main/scala/tilelink/Broadcast.scala 424:{24,24}]
    sent_d <= reset | _GEN_25; // @[src/main/scala/tilelink/Broadcast.scala 425:{24,24}]
    shared <= io_probesack | _GEN_15; // @[src/main/scala/tilelink/Broadcast.scala 473:23 474:12]
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      opcode <= io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 443:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      size <= io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      source <= io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 446:13]
    end
    if (reset) begin // @[src/main/scala/tilelink/Broadcast.scala 433:24]
      address <= 32'h0; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
    end else if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      address <= io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 449:13]
    end
    count <= _GEN_27[0];
    line_443_valid_reg <= _T_1;
    line_444_valid_reg <= _T_3;
    line_445_valid_reg <= _T_4;
    line_446_valid_reg <= io_probe_valid;
    line_447_valid_reg <= io_d_last;
    line_448_valid_reg <= _T_3;
    line_449_valid_reg <= _T_8;
    line_450_valid_reg <= io_e_last;
    line_451_valid_reg <= _T_3;
    line_452_valid_reg <= _T_12;
    line_453_valid_reg <= _T_13;
    line_454_valid_reg <= _T_3;
    line_455_valid_reg <= _T_17;
    line_456_valid_reg <= io_probesack;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:439 assert (idle)\n"); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n"); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_e_last & _T_3 & ~(~got_e)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n"); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_3 & ~(count > 1'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n"); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shared = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  opcode = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  source = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  address = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  count = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_443_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_444_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_445_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_446_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_447_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_448_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_449_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_450_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_451_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_452_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_453_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_454_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_455_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_456_valid_reg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_1 & ~reset) begin
      assert(idle); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
    end
    //
    if (io_d_last & _T_3) begin
      assert(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
    end
    //
    if (io_e_last & _T_3) begin
      assert(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
    end
    //
    if (_T_13 & _T_3) begin
      assert(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
    end
  end
endmodule
module Queue_37(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_mask [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_457_clock;
  wire  line_457_reset;
  wire  line_457_valid;
  reg  line_457_valid_reg;
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_458_clock;
  wire  line_458_reset;
  wire  line_458_valid;
  reg  line_458_valid_reg;
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_459_clock;
  wire  line_459_reset;
  wire  line_459_valid;
  reg  line_459_valid_reg;
  GEN_w1_line #(.COVER_INDEX(457)) line_457 (
    .clock(line_457_clock),
    .reset(line_457_reset),
    .valid(line_457_valid)
  );
  GEN_w1_line #(.COVER_INDEX(458)) line_458 (
    .clock(line_458_clock),
    .reset(line_458_reset),
    .valid(line_458_valid)
  );
  GEN_w1_line #(.COVER_INDEX(459)) line_459 (
    .clock(line_459_clock),
    .reset(line_459_reset),
    .valid(line_459_valid)
  );
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_457_clock = clock;
  assign line_457_reset = reset;
  assign line_457_valid = do_enq ^ line_457_valid_reg;
  assign line_458_clock = clock;
  assign line_458_reset = reset;
  assign line_458_valid = do_deq ^ line_458_valid_reg;
  assign line_459_clock = clock;
  assign line_459_reset = reset;
  assign line_459_valid = _T ^ line_459_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_457_valid_reg <= do_enq;
    line_458_valid_reg <= do_deq;
    line_459_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_457_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_458_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_459_valid_reg = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_1(
  input         clock,
  input         reset,
  input         io_in_a_first, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_in_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_in_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [1:0]  io_in_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [31:0] io_in_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [7:0]  io_in_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [63:0] io_in_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_out_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_out_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [3:0]  io_out_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [31:0] io_out_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [7:0]  io_out_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [63:0] io_out_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_bits_count, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probenack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probedack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probesack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_d_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_e_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [1:0]  io_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [26:0] io_line, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_idle, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_need_d // @[src/main/scala/tilelink/Broadcast.scala 401:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  reg  got_e; // @[src/main/scala/tilelink/Broadcast.scala 424:24]
  reg  sent_d; // @[src/main/scala/tilelink/Broadcast.scala 425:24]
  reg  shared; // @[src/main/scala/tilelink/Broadcast.scala 426:20]
  reg [2:0] opcode; // @[src/main/scala/tilelink/Broadcast.scala 427:20]
  reg [2:0] size; // @[src/main/scala/tilelink/Broadcast.scala 429:20]
  reg [1:0] source; // @[src/main/scala/tilelink/Broadcast.scala 430:20]
  reg [31:0] address; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
  reg  count; // @[src/main/scala/tilelink/Broadcast.scala 434:20]
  wire  idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 438:22]
  wire  line_460_clock;
  wire  line_460_reset;
  wire  line_460_valid;
  reg  line_460_valid_reg;
  wire  _T_3 = ~reset; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_461_clock;
  wire  line_461_reset;
  wire  line_461_valid;
  reg  line_461_valid_reg;
  wire  _T_4 = ~idle; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_462_clock;
  wire  line_462_reset;
  wire  line_462_valid;
  reg  line_462_valid_reg;
  wire  _GEN_14 = _T & io_in_a_first ? 1'h0 : sent_d; // @[src/main/scala/tilelink/Broadcast.scala 438:40 440:13 425:24]
  wire  _GEN_15 = _T & io_in_a_first ? 1'h0 : shared; // @[src/main/scala/tilelink/Broadcast.scala 438:40 441:13 426:20]
  wire  _GEN_16 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[src/main/scala/tilelink/Broadcast.scala 438:40 442:13 424:24]
  wire  _GEN_22 = _T & io_in_a_first | count; // @[src/main/scala/tilelink/Broadcast.scala 438:40 450:13 434:20]
  wire  line_463_clock;
  wire  line_463_reset;
  wire  line_463_valid;
  reg  line_463_valid_reg;
  wire  _GEN_23 = io_probe_valid ? io_probe_bits_count : _GEN_22; // @[src/main/scala/tilelink/Broadcast.scala 454:25 455:13]
  wire  line_464_clock;
  wire  line_464_reset;
  wire  line_464_valid;
  reg  line_464_valid_reg;
  wire  line_465_clock;
  wire  line_465_reset;
  wire  line_465_valid;
  reg  line_465_valid_reg;
  wire  _T_8 = ~(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
  wire  line_466_clock;
  wire  line_466_reset;
  wire  line_466_valid;
  reg  line_466_valid_reg;
  wire  _GEN_25 = io_d_last | _GEN_14; // @[src/main/scala/tilelink/Broadcast.scala 459:20 461:12]
  wire  line_467_clock;
  wire  line_467_reset;
  wire  line_467_valid;
  reg  line_467_valid_reg;
  wire  line_468_clock;
  wire  line_468_reset;
  wire  line_468_valid;
  reg  line_468_valid_reg;
  wire  _T_12 = ~(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
  wire  line_469_clock;
  wire  line_469_reset;
  wire  line_469_valid;
  reg  line_469_valid_reg;
  wire  _GEN_26 = io_e_last | _GEN_16; // @[src/main/scala/tilelink/Broadcast.scala 463:20 465:11]
  wire  _T_13 = io_probenack | io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 468:22]
  wire  line_470_clock;
  wire  line_470_reset;
  wire  line_470_valid;
  reg  line_470_valid_reg;
  wire  line_471_clock;
  wire  line_471_reset;
  wire  line_471_valid;
  reg  line_471_valid_reg;
  wire  _T_17 = ~(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
  wire  line_472_clock;
  wire  line_472_reset;
  wire  line_472_valid;
  reg  line_472_valid_reg;
  wire [1:0] _count_T_1 = io_probenack & io_probedack ? 2'h2 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 470:25]
  wire [1:0] _GEN_29 = {{1'd0}, count}; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _count_T_3 = _GEN_29 - _count_T_1; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _GEN_27 = io_probenack | io_probedack ? _count_T_3 : {{1'd0}, _GEN_23}; // @[src/main/scala/tilelink/Broadcast.scala 468:39 470:11]
  wire  line_473_clock;
  wire  line_473_reset;
  wire  line_473_valid;
  reg  line_473_valid_reg;
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 486:26]
  wire  i_data_ready = o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 385:17 src/main/scala/tilelink/Broadcast.scala 483:20]
  wire  probe_done = ~count; // @[src/main/scala/tilelink/Broadcast.scala 491:26]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[src/main/scala/tilelink/Broadcast.scala 492:52]
  wire [1:0] transform = shared ? 2'h2 : 2'h3; // @[src/main/scala/tilelink/Broadcast.scala 494:22]
  wire [1:0] _io_out_a_bits_source_T = acquire ? transform : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 501:35]
  Queue_37 o_data_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(o_data_q_clock),
    .reset(o_data_q_reset),
    .io_enq_ready(o_data_q_io_enq_ready),
    .io_enq_valid(o_data_q_io_enq_valid),
    .io_enq_bits_mask(o_data_q_io_enq_bits_mask),
    .io_enq_bits_data(o_data_q_io_enq_bits_data),
    .io_deq_ready(o_data_q_io_deq_ready),
    .io_deq_valid(o_data_q_io_deq_valid),
    .io_deq_bits_mask(o_data_q_io_deq_bits_mask),
    .io_deq_bits_data(o_data_q_io_deq_bits_data)
  );
  GEN_w1_line #(.COVER_INDEX(460)) line_460 (
    .clock(line_460_clock),
    .reset(line_460_reset),
    .valid(line_460_valid)
  );
  GEN_w1_line #(.COVER_INDEX(461)) line_461 (
    .clock(line_461_clock),
    .reset(line_461_reset),
    .valid(line_461_valid)
  );
  GEN_w1_line #(.COVER_INDEX(462)) line_462 (
    .clock(line_462_clock),
    .reset(line_462_reset),
    .valid(line_462_valid)
  );
  GEN_w1_line #(.COVER_INDEX(463)) line_463 (
    .clock(line_463_clock),
    .reset(line_463_reset),
    .valid(line_463_valid)
  );
  GEN_w1_line #(.COVER_INDEX(464)) line_464 (
    .clock(line_464_clock),
    .reset(line_464_reset),
    .valid(line_464_valid)
  );
  GEN_w1_line #(.COVER_INDEX(465)) line_465 (
    .clock(line_465_clock),
    .reset(line_465_reset),
    .valid(line_465_valid)
  );
  GEN_w1_line #(.COVER_INDEX(466)) line_466 (
    .clock(line_466_clock),
    .reset(line_466_reset),
    .valid(line_466_valid)
  );
  GEN_w1_line #(.COVER_INDEX(467)) line_467 (
    .clock(line_467_clock),
    .reset(line_467_reset),
    .valid(line_467_valid)
  );
  GEN_w1_line #(.COVER_INDEX(468)) line_468 (
    .clock(line_468_clock),
    .reset(line_468_reset),
    .valid(line_468_valid)
  );
  GEN_w1_line #(.COVER_INDEX(469)) line_469 (
    .clock(line_469_clock),
    .reset(line_469_reset),
    .valid(line_469_valid)
  );
  GEN_w1_line #(.COVER_INDEX(470)) line_470 (
    .clock(line_470_clock),
    .reset(line_470_reset),
    .valid(line_470_valid)
  );
  GEN_w1_line #(.COVER_INDEX(471)) line_471 (
    .clock(line_471_clock),
    .reset(line_471_reset),
    .valid(line_471_valid)
  );
  GEN_w1_line #(.COVER_INDEX(472)) line_472 (
    .clock(line_472_clock),
    .reset(line_472_reset),
    .valid(line_472_valid)
  );
  GEN_w1_line #(.COVER_INDEX(473)) line_473 (
    .clock(line_473_clock),
    .reset(line_473_reset),
    .valid(line_473_valid)
  );
  assign line_460_clock = clock;
  assign line_460_reset = reset;
  assign line_460_valid = _T_1 ^ line_460_valid_reg;
  assign line_461_clock = clock;
  assign line_461_reset = reset;
  assign line_461_valid = _T_3 ^ line_461_valid_reg;
  assign line_462_clock = clock;
  assign line_462_reset = reset;
  assign line_462_valid = _T_4 ^ line_462_valid_reg;
  assign line_463_clock = clock;
  assign line_463_reset = reset;
  assign line_463_valid = io_probe_valid ^ line_463_valid_reg;
  assign line_464_clock = clock;
  assign line_464_reset = reset;
  assign line_464_valid = io_d_last ^ line_464_valid_reg;
  assign line_465_clock = clock;
  assign line_465_reset = reset;
  assign line_465_valid = _T_3 ^ line_465_valid_reg;
  assign line_466_clock = clock;
  assign line_466_reset = reset;
  assign line_466_valid = _T_8 ^ line_466_valid_reg;
  assign line_467_clock = clock;
  assign line_467_reset = reset;
  assign line_467_valid = io_e_last ^ line_467_valid_reg;
  assign line_468_clock = clock;
  assign line_468_reset = reset;
  assign line_468_valid = _T_3 ^ line_468_valid_reg;
  assign line_469_clock = clock;
  assign line_469_reset = reset;
  assign line_469_valid = _T_12 ^ line_469_valid_reg;
  assign line_470_clock = clock;
  assign line_470_reset = reset;
  assign line_470_valid = _T_13 ^ line_470_valid_reg;
  assign line_471_clock = clock;
  assign line_471_reset = reset;
  assign line_471_valid = _T_3 ^ line_471_valid_reg;
  assign line_472_clock = clock;
  assign line_472_reset = reset;
  assign line_472_valid = _T_17 ^ line_472_valid_reg;
  assign line_473_clock = clock;
  assign line_473_reset = reset;
  assign line_473_valid = io_probesack ^ line_473_valid_reg;
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[src/main/scala/tilelink/Broadcast.scala 486:45]
  assign io_out_a_valid = o_data_q_io_deq_valid & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 497:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[src/main/scala/tilelink/Broadcast.scala 498:31]
  assign io_out_a_bits_size = size; // @[src/main/scala/tilelink/Broadcast.scala 500:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[src/main/scala/tilelink/Broadcast.scala 501:31]
  assign io_out_a_bits_address = address; // @[src/main/scala/tilelink/Broadcast.scala 502:25]
  assign io_out_a_bits_mask = o_data_q_io_deq_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 503:25]
  assign io_out_a_bits_data = o_data_q_io_deq_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 504:25]
  assign io_source = source; // @[src/main/scala/tilelink/Broadcast.scala 479:13]
  assign io_line = address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 480:22]
  assign io_idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  assign io_need_d = ~sent_d; // @[src/main/scala/tilelink/Broadcast.scala 478:16]
  assign o_data_q_clock = clock;
  assign o_data_q_reset = reset;
  assign o_data_q_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 487:44]
  assign o_data_q_io_enq_bits_mask = io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 483:20 488:20]
  assign o_data_q_io_enq_bits_data = io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 483:20 489:20]
  assign o_data_q_io_deq_ready = io_out_a_ready & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 496:34]
  always @(posedge clock) begin
    got_e <= reset | _GEN_26; // @[src/main/scala/tilelink/Broadcast.scala 424:{24,24}]
    sent_d <= reset | _GEN_25; // @[src/main/scala/tilelink/Broadcast.scala 425:{24,24}]
    shared <= io_probesack | _GEN_15; // @[src/main/scala/tilelink/Broadcast.scala 473:23 474:12]
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      opcode <= io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 443:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      size <= io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      source <= io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 446:13]
    end
    if (reset) begin // @[src/main/scala/tilelink/Broadcast.scala 433:24]
      address <= 32'h20; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
    end else if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      address <= io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 449:13]
    end
    count <= _GEN_27[0];
    line_460_valid_reg <= _T_1;
    line_461_valid_reg <= _T_3;
    line_462_valid_reg <= _T_4;
    line_463_valid_reg <= io_probe_valid;
    line_464_valid_reg <= io_d_last;
    line_465_valid_reg <= _T_3;
    line_466_valid_reg <= _T_8;
    line_467_valid_reg <= io_e_last;
    line_468_valid_reg <= _T_3;
    line_469_valid_reg <= _T_12;
    line_470_valid_reg <= _T_13;
    line_471_valid_reg <= _T_3;
    line_472_valid_reg <= _T_17;
    line_473_valid_reg <= io_probesack;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:439 assert (idle)\n"); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n"); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_e_last & _T_3 & ~(~got_e)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n"); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_3 & ~(count > 1'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n"); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shared = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  opcode = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  source = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  address = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  count = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_460_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_461_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_462_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_463_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_464_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_465_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_466_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_467_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_468_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_469_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_470_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_471_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_472_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_473_valid_reg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_1 & ~reset) begin
      assert(idle); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
    end
    //
    if (io_d_last & _T_3) begin
      assert(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
    end
    //
    if (io_e_last & _T_3) begin
      assert(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
    end
    //
    if (_T_13 & _T_3) begin
      assert(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
    end
  end
endmodule
module Queue_38(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_mask [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_474_clock;
  wire  line_474_reset;
  wire  line_474_valid;
  reg  line_474_valid_reg;
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_475_clock;
  wire  line_475_reset;
  wire  line_475_valid;
  reg  line_475_valid_reg;
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_476_clock;
  wire  line_476_reset;
  wire  line_476_valid;
  reg  line_476_valid_reg;
  GEN_w1_line #(.COVER_INDEX(474)) line_474 (
    .clock(line_474_clock),
    .reset(line_474_reset),
    .valid(line_474_valid)
  );
  GEN_w1_line #(.COVER_INDEX(475)) line_475 (
    .clock(line_475_clock),
    .reset(line_475_reset),
    .valid(line_475_valid)
  );
  GEN_w1_line #(.COVER_INDEX(476)) line_476 (
    .clock(line_476_clock),
    .reset(line_476_reset),
    .valid(line_476_valid)
  );
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_474_clock = clock;
  assign line_474_reset = reset;
  assign line_474_valid = do_enq ^ line_474_valid_reg;
  assign line_475_clock = clock;
  assign line_475_reset = reset;
  assign line_475_valid = do_deq ^ line_475_valid_reg;
  assign line_476_clock = clock;
  assign line_476_reset = reset;
  assign line_476_valid = _T ^ line_476_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_474_valid_reg <= do_enq;
    line_475_valid_reg <= do_deq;
    line_476_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_474_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_475_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_476_valid_reg = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_2(
  input         clock,
  input         reset,
  input         io_in_a_first, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_in_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_in_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [1:0]  io_in_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [31:0] io_in_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [7:0]  io_in_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [63:0] io_in_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_out_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_out_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [3:0]  io_out_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [31:0] io_out_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [7:0]  io_out_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [63:0] io_out_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_bits_count, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probenack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probedack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probesack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_d_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_e_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [1:0]  io_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [26:0] io_line, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_idle, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_need_d // @[src/main/scala/tilelink/Broadcast.scala 401:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  reg  got_e; // @[src/main/scala/tilelink/Broadcast.scala 424:24]
  reg  sent_d; // @[src/main/scala/tilelink/Broadcast.scala 425:24]
  reg  shared; // @[src/main/scala/tilelink/Broadcast.scala 426:20]
  reg [2:0] opcode; // @[src/main/scala/tilelink/Broadcast.scala 427:20]
  reg [2:0] size; // @[src/main/scala/tilelink/Broadcast.scala 429:20]
  reg [1:0] source; // @[src/main/scala/tilelink/Broadcast.scala 430:20]
  reg [31:0] address; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
  reg  count; // @[src/main/scala/tilelink/Broadcast.scala 434:20]
  wire  idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 438:22]
  wire  line_477_clock;
  wire  line_477_reset;
  wire  line_477_valid;
  reg  line_477_valid_reg;
  wire  _T_3 = ~reset; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_478_clock;
  wire  line_478_reset;
  wire  line_478_valid;
  reg  line_478_valid_reg;
  wire  _T_4 = ~idle; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_479_clock;
  wire  line_479_reset;
  wire  line_479_valid;
  reg  line_479_valid_reg;
  wire  _GEN_14 = _T & io_in_a_first ? 1'h0 : sent_d; // @[src/main/scala/tilelink/Broadcast.scala 438:40 440:13 425:24]
  wire  _GEN_15 = _T & io_in_a_first ? 1'h0 : shared; // @[src/main/scala/tilelink/Broadcast.scala 438:40 441:13 426:20]
  wire  _GEN_16 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[src/main/scala/tilelink/Broadcast.scala 438:40 442:13 424:24]
  wire  _GEN_22 = _T & io_in_a_first | count; // @[src/main/scala/tilelink/Broadcast.scala 438:40 450:13 434:20]
  wire  line_480_clock;
  wire  line_480_reset;
  wire  line_480_valid;
  reg  line_480_valid_reg;
  wire  _GEN_23 = io_probe_valid ? io_probe_bits_count : _GEN_22; // @[src/main/scala/tilelink/Broadcast.scala 454:25 455:13]
  wire  line_481_clock;
  wire  line_481_reset;
  wire  line_481_valid;
  reg  line_481_valid_reg;
  wire  line_482_clock;
  wire  line_482_reset;
  wire  line_482_valid;
  reg  line_482_valid_reg;
  wire  _T_8 = ~(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
  wire  line_483_clock;
  wire  line_483_reset;
  wire  line_483_valid;
  reg  line_483_valid_reg;
  wire  _GEN_25 = io_d_last | _GEN_14; // @[src/main/scala/tilelink/Broadcast.scala 459:20 461:12]
  wire  line_484_clock;
  wire  line_484_reset;
  wire  line_484_valid;
  reg  line_484_valid_reg;
  wire  line_485_clock;
  wire  line_485_reset;
  wire  line_485_valid;
  reg  line_485_valid_reg;
  wire  _T_12 = ~(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
  wire  line_486_clock;
  wire  line_486_reset;
  wire  line_486_valid;
  reg  line_486_valid_reg;
  wire  _GEN_26 = io_e_last | _GEN_16; // @[src/main/scala/tilelink/Broadcast.scala 463:20 465:11]
  wire  _T_13 = io_probenack | io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 468:22]
  wire  line_487_clock;
  wire  line_487_reset;
  wire  line_487_valid;
  reg  line_487_valid_reg;
  wire  line_488_clock;
  wire  line_488_reset;
  wire  line_488_valid;
  reg  line_488_valid_reg;
  wire  _T_17 = ~(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
  wire  line_489_clock;
  wire  line_489_reset;
  wire  line_489_valid;
  reg  line_489_valid_reg;
  wire [1:0] _count_T_1 = io_probenack & io_probedack ? 2'h2 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 470:25]
  wire [1:0] _GEN_29 = {{1'd0}, count}; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _count_T_3 = _GEN_29 - _count_T_1; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _GEN_27 = io_probenack | io_probedack ? _count_T_3 : {{1'd0}, _GEN_23}; // @[src/main/scala/tilelink/Broadcast.scala 468:39 470:11]
  wire  line_490_clock;
  wire  line_490_reset;
  wire  line_490_valid;
  reg  line_490_valid_reg;
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 486:26]
  wire  i_data_ready = o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 385:17 src/main/scala/tilelink/Broadcast.scala 483:20]
  wire  probe_done = ~count; // @[src/main/scala/tilelink/Broadcast.scala 491:26]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[src/main/scala/tilelink/Broadcast.scala 492:52]
  wire [1:0] transform = shared ? 2'h2 : 2'h3; // @[src/main/scala/tilelink/Broadcast.scala 494:22]
  wire [1:0] _io_out_a_bits_source_T = acquire ? transform : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 501:35]
  Queue_38 o_data_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(o_data_q_clock),
    .reset(o_data_q_reset),
    .io_enq_ready(o_data_q_io_enq_ready),
    .io_enq_valid(o_data_q_io_enq_valid),
    .io_enq_bits_mask(o_data_q_io_enq_bits_mask),
    .io_enq_bits_data(o_data_q_io_enq_bits_data),
    .io_deq_ready(o_data_q_io_deq_ready),
    .io_deq_valid(o_data_q_io_deq_valid),
    .io_deq_bits_mask(o_data_q_io_deq_bits_mask),
    .io_deq_bits_data(o_data_q_io_deq_bits_data)
  );
  GEN_w1_line #(.COVER_INDEX(477)) line_477 (
    .clock(line_477_clock),
    .reset(line_477_reset),
    .valid(line_477_valid)
  );
  GEN_w1_line #(.COVER_INDEX(478)) line_478 (
    .clock(line_478_clock),
    .reset(line_478_reset),
    .valid(line_478_valid)
  );
  GEN_w1_line #(.COVER_INDEX(479)) line_479 (
    .clock(line_479_clock),
    .reset(line_479_reset),
    .valid(line_479_valid)
  );
  GEN_w1_line #(.COVER_INDEX(480)) line_480 (
    .clock(line_480_clock),
    .reset(line_480_reset),
    .valid(line_480_valid)
  );
  GEN_w1_line #(.COVER_INDEX(481)) line_481 (
    .clock(line_481_clock),
    .reset(line_481_reset),
    .valid(line_481_valid)
  );
  GEN_w1_line #(.COVER_INDEX(482)) line_482 (
    .clock(line_482_clock),
    .reset(line_482_reset),
    .valid(line_482_valid)
  );
  GEN_w1_line #(.COVER_INDEX(483)) line_483 (
    .clock(line_483_clock),
    .reset(line_483_reset),
    .valid(line_483_valid)
  );
  GEN_w1_line #(.COVER_INDEX(484)) line_484 (
    .clock(line_484_clock),
    .reset(line_484_reset),
    .valid(line_484_valid)
  );
  GEN_w1_line #(.COVER_INDEX(485)) line_485 (
    .clock(line_485_clock),
    .reset(line_485_reset),
    .valid(line_485_valid)
  );
  GEN_w1_line #(.COVER_INDEX(486)) line_486 (
    .clock(line_486_clock),
    .reset(line_486_reset),
    .valid(line_486_valid)
  );
  GEN_w1_line #(.COVER_INDEX(487)) line_487 (
    .clock(line_487_clock),
    .reset(line_487_reset),
    .valid(line_487_valid)
  );
  GEN_w1_line #(.COVER_INDEX(488)) line_488 (
    .clock(line_488_clock),
    .reset(line_488_reset),
    .valid(line_488_valid)
  );
  GEN_w1_line #(.COVER_INDEX(489)) line_489 (
    .clock(line_489_clock),
    .reset(line_489_reset),
    .valid(line_489_valid)
  );
  GEN_w1_line #(.COVER_INDEX(490)) line_490 (
    .clock(line_490_clock),
    .reset(line_490_reset),
    .valid(line_490_valid)
  );
  assign line_477_clock = clock;
  assign line_477_reset = reset;
  assign line_477_valid = _T_1 ^ line_477_valid_reg;
  assign line_478_clock = clock;
  assign line_478_reset = reset;
  assign line_478_valid = _T_3 ^ line_478_valid_reg;
  assign line_479_clock = clock;
  assign line_479_reset = reset;
  assign line_479_valid = _T_4 ^ line_479_valid_reg;
  assign line_480_clock = clock;
  assign line_480_reset = reset;
  assign line_480_valid = io_probe_valid ^ line_480_valid_reg;
  assign line_481_clock = clock;
  assign line_481_reset = reset;
  assign line_481_valid = io_d_last ^ line_481_valid_reg;
  assign line_482_clock = clock;
  assign line_482_reset = reset;
  assign line_482_valid = _T_3 ^ line_482_valid_reg;
  assign line_483_clock = clock;
  assign line_483_reset = reset;
  assign line_483_valid = _T_8 ^ line_483_valid_reg;
  assign line_484_clock = clock;
  assign line_484_reset = reset;
  assign line_484_valid = io_e_last ^ line_484_valid_reg;
  assign line_485_clock = clock;
  assign line_485_reset = reset;
  assign line_485_valid = _T_3 ^ line_485_valid_reg;
  assign line_486_clock = clock;
  assign line_486_reset = reset;
  assign line_486_valid = _T_12 ^ line_486_valid_reg;
  assign line_487_clock = clock;
  assign line_487_reset = reset;
  assign line_487_valid = _T_13 ^ line_487_valid_reg;
  assign line_488_clock = clock;
  assign line_488_reset = reset;
  assign line_488_valid = _T_3 ^ line_488_valid_reg;
  assign line_489_clock = clock;
  assign line_489_reset = reset;
  assign line_489_valid = _T_17 ^ line_489_valid_reg;
  assign line_490_clock = clock;
  assign line_490_reset = reset;
  assign line_490_valid = io_probesack ^ line_490_valid_reg;
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[src/main/scala/tilelink/Broadcast.scala 486:45]
  assign io_out_a_valid = o_data_q_io_deq_valid & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 497:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[src/main/scala/tilelink/Broadcast.scala 498:31]
  assign io_out_a_bits_size = size; // @[src/main/scala/tilelink/Broadcast.scala 500:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[src/main/scala/tilelink/Broadcast.scala 501:31]
  assign io_out_a_bits_address = address; // @[src/main/scala/tilelink/Broadcast.scala 502:25]
  assign io_out_a_bits_mask = o_data_q_io_deq_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 503:25]
  assign io_out_a_bits_data = o_data_q_io_deq_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 504:25]
  assign io_source = source; // @[src/main/scala/tilelink/Broadcast.scala 479:13]
  assign io_line = address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 480:22]
  assign io_idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  assign io_need_d = ~sent_d; // @[src/main/scala/tilelink/Broadcast.scala 478:16]
  assign o_data_q_clock = clock;
  assign o_data_q_reset = reset;
  assign o_data_q_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 487:44]
  assign o_data_q_io_enq_bits_mask = io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 483:20 488:20]
  assign o_data_q_io_enq_bits_data = io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 483:20 489:20]
  assign o_data_q_io_deq_ready = io_out_a_ready & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 496:34]
  always @(posedge clock) begin
    got_e <= reset | _GEN_26; // @[src/main/scala/tilelink/Broadcast.scala 424:{24,24}]
    sent_d <= reset | _GEN_25; // @[src/main/scala/tilelink/Broadcast.scala 425:{24,24}]
    shared <= io_probesack | _GEN_15; // @[src/main/scala/tilelink/Broadcast.scala 473:23 474:12]
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      opcode <= io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 443:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      size <= io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      source <= io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 446:13]
    end
    if (reset) begin // @[src/main/scala/tilelink/Broadcast.scala 433:24]
      address <= 32'h40; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
    end else if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      address <= io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 449:13]
    end
    count <= _GEN_27[0];
    line_477_valid_reg <= _T_1;
    line_478_valid_reg <= _T_3;
    line_479_valid_reg <= _T_4;
    line_480_valid_reg <= io_probe_valid;
    line_481_valid_reg <= io_d_last;
    line_482_valid_reg <= _T_3;
    line_483_valid_reg <= _T_8;
    line_484_valid_reg <= io_e_last;
    line_485_valid_reg <= _T_3;
    line_486_valid_reg <= _T_12;
    line_487_valid_reg <= _T_13;
    line_488_valid_reg <= _T_3;
    line_489_valid_reg <= _T_17;
    line_490_valid_reg <= io_probesack;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:439 assert (idle)\n"); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n"); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_e_last & _T_3 & ~(~got_e)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n"); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_3 & ~(count > 1'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n"); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shared = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  opcode = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  source = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  address = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  count = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_477_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_478_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_479_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_480_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_481_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_482_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_483_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_484_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_485_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_486_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_487_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_488_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_489_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_490_valid_reg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_1 & ~reset) begin
      assert(idle); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
    end
    //
    if (io_d_last & _T_3) begin
      assert(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
    end
    //
    if (io_e_last & _T_3) begin
      assert(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
    end
    //
    if (_T_13 & _T_3) begin
      assert(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
    end
  end
endmodule
module Queue_39(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_mask [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:3]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_491_clock;
  wire  line_491_reset;
  wire  line_491_valid;
  reg  line_491_valid_reg;
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  line_492_clock;
  wire  line_492_reset;
  wire  line_492_valid;
  reg  line_492_valid_reg;
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_493_clock;
  wire  line_493_reset;
  wire  line_493_valid;
  reg  line_493_valid_reg;
  GEN_w1_line #(.COVER_INDEX(491)) line_491 (
    .clock(line_491_clock),
    .reset(line_491_reset),
    .valid(line_491_valid)
  );
  GEN_w1_line #(.COVER_INDEX(492)) line_492 (
    .clock(line_492_clock),
    .reset(line_492_reset),
    .valid(line_492_valid)
  );
  GEN_w1_line #(.COVER_INDEX(493)) line_493 (
    .clock(line_493_clock),
    .reset(line_493_reset),
    .valid(line_493_valid)
  );
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_491_clock = clock;
  assign line_491_reset = reset;
  assign line_491_valid = do_enq ^ line_491_valid_reg;
  assign line_492_clock = clock;
  assign line_492_reset = reset;
  assign line_492_valid = do_deq ^ line_492_valid_reg;
  assign line_493_clock = clock;
  assign line_493_reset = reset;
  assign line_493_valid = _T ^ line_493_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_491_valid_reg <= do_enq;
    line_492_valid_reg <= do_deq;
    line_493_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_mask[initvar] = _RAND_0[7:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_491_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_492_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_493_valid_reg = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBroadcastTracker_3(
  input         clock,
  input         reset,
  input         io_in_a_first, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_in_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_in_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [2:0]  io_in_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [1:0]  io_in_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [31:0] io_in_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [7:0]  io_in_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input  [63:0] io_in_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_out_a_ready, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_out_a_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_opcode, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [2:0]  io_out_a_bits_size, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [3:0]  io_out_a_bits_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [31:0] io_out_a_bits_address, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [7:0]  io_out_a_bits_mask, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [63:0] io_out_a_bits_data, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_valid, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probe_bits_count, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probenack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probedack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_probesack, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_d_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  input         io_e_last, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [1:0]  io_source, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output [26:0] io_line, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_idle, // @[src/main/scala/tilelink/Broadcast.scala 401:14]
  output        io_need_d // @[src/main/scala/tilelink/Broadcast.scala 401:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  o_data_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  o_data_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] o_data_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] o_data_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  reg  got_e; // @[src/main/scala/tilelink/Broadcast.scala 424:24]
  reg  sent_d; // @[src/main/scala/tilelink/Broadcast.scala 425:24]
  reg  shared; // @[src/main/scala/tilelink/Broadcast.scala 426:20]
  reg [2:0] opcode; // @[src/main/scala/tilelink/Broadcast.scala 427:20]
  reg [2:0] size; // @[src/main/scala/tilelink/Broadcast.scala 429:20]
  reg [1:0] source; // @[src/main/scala/tilelink/Broadcast.scala 430:20]
  reg [31:0] address; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
  reg  count; // @[src/main/scala/tilelink/Broadcast.scala 434:20]
  wire  idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  wire  _T = io_in_a_ready & io_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = _T & io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 438:22]
  wire  line_494_clock;
  wire  line_494_reset;
  wire  line_494_valid;
  reg  line_494_valid_reg;
  wire  _T_3 = ~reset; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_495_clock;
  wire  line_495_reset;
  wire  line_495_valid;
  reg  line_495_valid_reg;
  wire  _T_4 = ~idle; // @[src/main/scala/tilelink/Broadcast.scala 439:12]
  wire  line_496_clock;
  wire  line_496_reset;
  wire  line_496_valid;
  reg  line_496_valid_reg;
  wire  _GEN_14 = _T & io_in_a_first ? 1'h0 : sent_d; // @[src/main/scala/tilelink/Broadcast.scala 438:40 440:13 425:24]
  wire  _GEN_15 = _T & io_in_a_first ? 1'h0 : shared; // @[src/main/scala/tilelink/Broadcast.scala 438:40 441:13 426:20]
  wire  _GEN_16 = _T & io_in_a_first ? io_in_a_bits_opcode != 3'h6 & io_in_a_bits_opcode != 3'h7 : got_e; // @[src/main/scala/tilelink/Broadcast.scala 438:40 442:13 424:24]
  wire  _GEN_22 = _T & io_in_a_first | count; // @[src/main/scala/tilelink/Broadcast.scala 438:40 450:13 434:20]
  wire  line_497_clock;
  wire  line_497_reset;
  wire  line_497_valid;
  reg  line_497_valid_reg;
  wire  _GEN_23 = io_probe_valid ? io_probe_bits_count : _GEN_22; // @[src/main/scala/tilelink/Broadcast.scala 454:25 455:13]
  wire  line_498_clock;
  wire  line_498_reset;
  wire  line_498_valid;
  reg  line_498_valid_reg;
  wire  line_499_clock;
  wire  line_499_reset;
  wire  line_499_valid;
  reg  line_499_valid_reg;
  wire  _T_8 = ~(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
  wire  line_500_clock;
  wire  line_500_reset;
  wire  line_500_valid;
  reg  line_500_valid_reg;
  wire  _GEN_25 = io_d_last | _GEN_14; // @[src/main/scala/tilelink/Broadcast.scala 459:20 461:12]
  wire  line_501_clock;
  wire  line_501_reset;
  wire  line_501_valid;
  reg  line_501_valid_reg;
  wire  line_502_clock;
  wire  line_502_reset;
  wire  line_502_valid;
  reg  line_502_valid_reg;
  wire  _T_12 = ~(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
  wire  line_503_clock;
  wire  line_503_reset;
  wire  line_503_valid;
  reg  line_503_valid_reg;
  wire  _GEN_26 = io_e_last | _GEN_16; // @[src/main/scala/tilelink/Broadcast.scala 463:20 465:11]
  wire  _T_13 = io_probenack | io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 468:22]
  wire  line_504_clock;
  wire  line_504_reset;
  wire  line_504_valid;
  reg  line_504_valid_reg;
  wire  line_505_clock;
  wire  line_505_reset;
  wire  line_505_valid;
  reg  line_505_valid_reg;
  wire  _T_17 = ~(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
  wire  line_506_clock;
  wire  line_506_reset;
  wire  line_506_valid;
  reg  line_506_valid_reg;
  wire [1:0] _count_T_1 = io_probenack & io_probedack ? 2'h2 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 470:25]
  wire [1:0] _GEN_29 = {{1'd0}, count}; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _count_T_3 = _GEN_29 - _count_T_1; // @[src/main/scala/tilelink/Broadcast.scala 470:20]
  wire [1:0] _GEN_27 = io_probenack | io_probedack ? _count_T_3 : {{1'd0}, _GEN_23}; // @[src/main/scala/tilelink/Broadcast.scala 468:39 470:11]
  wire  line_507_clock;
  wire  line_507_reset;
  wire  line_507_valid;
  reg  line_507_valid_reg;
  wire  _io_in_a_ready_T_1 = idle | ~io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 486:26]
  wire  i_data_ready = o_data_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 385:17 src/main/scala/tilelink/Broadcast.scala 483:20]
  wire  probe_done = ~count; // @[src/main/scala/tilelink/Broadcast.scala 491:26]
  wire  acquire = opcode == 3'h6 | opcode == 3'h7; // @[src/main/scala/tilelink/Broadcast.scala 492:52]
  wire [1:0] transform = shared ? 2'h2 : 2'h3; // @[src/main/scala/tilelink/Broadcast.scala 494:22]
  wire [1:0] _io_out_a_bits_source_T = acquire ? transform : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 501:35]
  Queue_39 o_data_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(o_data_q_clock),
    .reset(o_data_q_reset),
    .io_enq_ready(o_data_q_io_enq_ready),
    .io_enq_valid(o_data_q_io_enq_valid),
    .io_enq_bits_mask(o_data_q_io_enq_bits_mask),
    .io_enq_bits_data(o_data_q_io_enq_bits_data),
    .io_deq_ready(o_data_q_io_deq_ready),
    .io_deq_valid(o_data_q_io_deq_valid),
    .io_deq_bits_mask(o_data_q_io_deq_bits_mask),
    .io_deq_bits_data(o_data_q_io_deq_bits_data)
  );
  GEN_w1_line #(.COVER_INDEX(494)) line_494 (
    .clock(line_494_clock),
    .reset(line_494_reset),
    .valid(line_494_valid)
  );
  GEN_w1_line #(.COVER_INDEX(495)) line_495 (
    .clock(line_495_clock),
    .reset(line_495_reset),
    .valid(line_495_valid)
  );
  GEN_w1_line #(.COVER_INDEX(496)) line_496 (
    .clock(line_496_clock),
    .reset(line_496_reset),
    .valid(line_496_valid)
  );
  GEN_w1_line #(.COVER_INDEX(497)) line_497 (
    .clock(line_497_clock),
    .reset(line_497_reset),
    .valid(line_497_valid)
  );
  GEN_w1_line #(.COVER_INDEX(498)) line_498 (
    .clock(line_498_clock),
    .reset(line_498_reset),
    .valid(line_498_valid)
  );
  GEN_w1_line #(.COVER_INDEX(499)) line_499 (
    .clock(line_499_clock),
    .reset(line_499_reset),
    .valid(line_499_valid)
  );
  GEN_w1_line #(.COVER_INDEX(500)) line_500 (
    .clock(line_500_clock),
    .reset(line_500_reset),
    .valid(line_500_valid)
  );
  GEN_w1_line #(.COVER_INDEX(501)) line_501 (
    .clock(line_501_clock),
    .reset(line_501_reset),
    .valid(line_501_valid)
  );
  GEN_w1_line #(.COVER_INDEX(502)) line_502 (
    .clock(line_502_clock),
    .reset(line_502_reset),
    .valid(line_502_valid)
  );
  GEN_w1_line #(.COVER_INDEX(503)) line_503 (
    .clock(line_503_clock),
    .reset(line_503_reset),
    .valid(line_503_valid)
  );
  GEN_w1_line #(.COVER_INDEX(504)) line_504 (
    .clock(line_504_clock),
    .reset(line_504_reset),
    .valid(line_504_valid)
  );
  GEN_w1_line #(.COVER_INDEX(505)) line_505 (
    .clock(line_505_clock),
    .reset(line_505_reset),
    .valid(line_505_valid)
  );
  GEN_w1_line #(.COVER_INDEX(506)) line_506 (
    .clock(line_506_clock),
    .reset(line_506_reset),
    .valid(line_506_valid)
  );
  GEN_w1_line #(.COVER_INDEX(507)) line_507 (
    .clock(line_507_clock),
    .reset(line_507_reset),
    .valid(line_507_valid)
  );
  assign line_494_clock = clock;
  assign line_494_reset = reset;
  assign line_494_valid = _T_1 ^ line_494_valid_reg;
  assign line_495_clock = clock;
  assign line_495_reset = reset;
  assign line_495_valid = _T_3 ^ line_495_valid_reg;
  assign line_496_clock = clock;
  assign line_496_reset = reset;
  assign line_496_valid = _T_4 ^ line_496_valid_reg;
  assign line_497_clock = clock;
  assign line_497_reset = reset;
  assign line_497_valid = io_probe_valid ^ line_497_valid_reg;
  assign line_498_clock = clock;
  assign line_498_reset = reset;
  assign line_498_valid = io_d_last ^ line_498_valid_reg;
  assign line_499_clock = clock;
  assign line_499_reset = reset;
  assign line_499_valid = _T_3 ^ line_499_valid_reg;
  assign line_500_clock = clock;
  assign line_500_reset = reset;
  assign line_500_valid = _T_8 ^ line_500_valid_reg;
  assign line_501_clock = clock;
  assign line_501_reset = reset;
  assign line_501_valid = io_e_last ^ line_501_valid_reg;
  assign line_502_clock = clock;
  assign line_502_reset = reset;
  assign line_502_valid = _T_3 ^ line_502_valid_reg;
  assign line_503_clock = clock;
  assign line_503_reset = reset;
  assign line_503_valid = _T_12 ^ line_503_valid_reg;
  assign line_504_clock = clock;
  assign line_504_reset = reset;
  assign line_504_valid = _T_13 ^ line_504_valid_reg;
  assign line_505_clock = clock;
  assign line_505_reset = reset;
  assign line_505_valid = _T_3 ^ line_505_valid_reg;
  assign line_506_clock = clock;
  assign line_506_reset = reset;
  assign line_506_valid = _T_17 ^ line_506_valid_reg;
  assign line_507_clock = clock;
  assign line_507_reset = reset;
  assign line_507_valid = io_probesack ^ line_507_valid_reg;
  assign io_in_a_ready = (idle | ~io_in_a_first) & i_data_ready; // @[src/main/scala/tilelink/Broadcast.scala 486:45]
  assign io_out_a_valid = o_data_q_io_deq_valid & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 497:34]
  assign io_out_a_bits_opcode = acquire ? 3'h4 : opcode; // @[src/main/scala/tilelink/Broadcast.scala 498:31]
  assign io_out_a_bits_size = size; // @[src/main/scala/tilelink/Broadcast.scala 500:25]
  assign io_out_a_bits_source = {_io_out_a_bits_source_T,source}; // @[src/main/scala/tilelink/Broadcast.scala 501:31]
  assign io_out_a_bits_address = address; // @[src/main/scala/tilelink/Broadcast.scala 502:25]
  assign io_out_a_bits_mask = o_data_q_io_deq_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 503:25]
  assign io_out_a_bits_data = o_data_q_io_deq_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 504:25]
  assign io_source = source; // @[src/main/scala/tilelink/Broadcast.scala 479:13]
  assign io_line = address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 480:22]
  assign io_idle = got_e & sent_d; // @[src/main/scala/tilelink/Broadcast.scala 436:23]
  assign io_need_d = ~sent_d; // @[src/main/scala/tilelink/Broadcast.scala 478:16]
  assign o_data_q_clock = clock;
  assign o_data_q_reset = reset;
  assign o_data_q_io_enq_valid = _io_in_a_ready_T_1 & io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 487:44]
  assign o_data_q_io_enq_bits_mask = io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 483:20 488:20]
  assign o_data_q_io_enq_bits_data = io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 483:20 489:20]
  assign o_data_q_io_deq_ready = io_out_a_ready & probe_done; // @[src/main/scala/tilelink/Broadcast.scala 496:34]
  always @(posedge clock) begin
    got_e <= reset | _GEN_26; // @[src/main/scala/tilelink/Broadcast.scala 424:{24,24}]
    sent_d <= reset | _GEN_25; // @[src/main/scala/tilelink/Broadcast.scala 425:{24,24}]
    shared <= io_probesack | _GEN_15; // @[src/main/scala/tilelink/Broadcast.scala 473:23 474:12]
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      opcode <= io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 443:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      size <= io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 445:13]
    end
    if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      source <= io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 446:13]
    end
    if (reset) begin // @[src/main/scala/tilelink/Broadcast.scala 433:24]
      address <= 32'h60; // @[src/main/scala/tilelink/Broadcast.scala 433:24]
    end else if (_T & io_in_a_first) begin // @[src/main/scala/tilelink/Broadcast.scala 438:40]
      address <= io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 449:13]
    end
    count <= _GEN_27[0];
    line_494_valid_reg <= _T_1;
    line_495_valid_reg <= _T_3;
    line_496_valid_reg <= _T_4;
    line_497_valid_reg <= io_probe_valid;
    line_498_valid_reg <= io_d_last;
    line_499_valid_reg <= _T_3;
    line_500_valid_reg <= _T_8;
    line_501_valid_reg <= io_e_last;
    line_502_valid_reg <= _T_3;
    line_503_valid_reg <= _T_12;
    line_504_valid_reg <= _T_13;
    line_505_valid_reg <= _T_3;
    line_506_valid_reg <= _T_17;
    line_507_valid_reg <= io_probesack;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~reset & ~idle) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:439 assert (idle)\n"); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_d_last & _T_3 & ~(~sent_d)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n"); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_e_last & _T_3 & ~(~got_e)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n"); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_3 & ~(count > 1'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n"); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  got_e = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sent_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shared = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  opcode = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  source = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  address = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  count = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_494_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_495_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_496_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_497_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_498_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_499_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_500_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_501_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_502_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_503_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_504_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_505_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_506_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_507_valid_reg = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_1 & ~reset) begin
      assert(idle); // @[src/main/scala/tilelink/Broadcast.scala 439:12]
    end
    //
    if (io_d_last & _T_3) begin
      assert(~sent_d); // @[src/main/scala/tilelink/Broadcast.scala 460:12]
    end
    //
    if (io_e_last & _T_3) begin
      assert(~got_e); // @[src/main/scala/tilelink/Broadcast.scala 464:12]
    end
    //
    if (_T_13 & _T_3) begin
      assert(count > 1'h0); // @[src/main/scala/tilelink/Broadcast.scala 469:12]
    end
  end
endmodule
module TLBroadcast(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  filter_clock; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_reset; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_request_ready; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_request_valid; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire [1:0] filter_io_request_bits_mshr; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire [31:0] filter_io_request_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_request_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_request_bits_needT; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_response_ready; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_response_valid; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire [1:0] filter_io_response_bits_mshr; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire [31:0] filter_io_response_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  filter_io_response_bits_needT; // @[src/main/scala/tilelink/Broadcast.scala 99:26]
  wire  TLBroadcastTracker_clock; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_reset; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_out_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_out_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_io_out_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [3:0] TLBroadcastTracker_io_out_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_io_out_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_io_out_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_io_out_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probe_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probe_bits_count; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probenack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_probesack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_d_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_e_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_io_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [26:0] TLBroadcastTracker_io_line; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_io_need_d; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_clock; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_reset; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_1_io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_1_io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_1_io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_1_io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_out_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_out_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_1_io_out_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [3:0] TLBroadcastTracker_1_io_out_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_1_io_out_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_1_io_out_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_1_io_out_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probe_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probe_bits_count; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probenack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_probesack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_d_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_e_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_1_io_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [26:0] TLBroadcastTracker_1_io_line; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_1_io_need_d; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_clock; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_reset; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_2_io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_2_io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_2_io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_2_io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_out_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_out_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_2_io_out_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [3:0] TLBroadcastTracker_2_io_out_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_2_io_out_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_2_io_out_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_2_io_out_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probe_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probe_bits_count; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probenack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_probesack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_d_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_e_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_2_io_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [26:0] TLBroadcastTracker_2_io_line; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_2_io_need_d; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_clock; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_reset; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_first; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_in_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_in_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_in_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_3_io_in_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_3_io_in_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_3_io_in_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_3_io_in_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_out_a_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_out_a_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [2:0] TLBroadcastTracker_3_io_out_a_bits_size; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [3:0] TLBroadcastTracker_3_io_out_a_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [31:0] TLBroadcastTracker_3_io_out_a_bits_address; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [7:0] TLBroadcastTracker_3_io_out_a_bits_mask; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [63:0] TLBroadcastTracker_3_io_out_a_bits_data; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probe_valid; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probe_bits_count; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probenack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probedack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_probesack; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_d_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_e_last; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [1:0] TLBroadcastTracker_3_io_source; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [26:0] TLBroadcastTracker_3_io_line; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire  TLBroadcastTracker_3_io_need_d; // @[src/main/scala/tilelink/Broadcast.scala 107:15]
  wire [3:0] _T = 4'h1 << auto_in_e_bits_sink; // @[src/main/scala/chisel3/util/OneHot.scala 58:35]
  wire [1:0] d_what = auto_out_d_bits_source[3:2]; // @[src/main/scala/tilelink/Broadcast.scala 118:37]
  wire  d_drop = d_what == 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 119:27]
  wire  d_hasData = auto_out_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  reg [1:0] beatsLeft; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
  wire  idle = beatsLeft == 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 61:28]
  wire  d_response = d_hasData | ~d_what[1]; // @[src/main/scala/tilelink/Broadcast.scala 140:34]
  reg [1:0] counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [2:0] _d_normal_bits_opcode_T = d_hasData ? 3'h5 : 3'h6; // @[src/main/scala/tilelink/Broadcast.scala 132:36]
  wire [2:0] d_normal_bits_opcode = d_what[1] ? _d_normal_bits_opcode_T : auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Broadcast.scala 130:21 131:24 132:30]
  wire  beats1_opdata = d_normal_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  wire [11:0] _beats1_decode_T_1 = 12'h1f << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beats1_decode = _beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire [1:0] beats1 = beats1_opdata ? beats1_decode : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire  d_last = counter == 2'h1 | beats1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  _d_normal_valid_T_1 = ~d_drop; // @[src/main/scala/tilelink/Broadcast.scala 129:51]
  wire  d_normal_valid = auto_out_d_valid & ~d_drop; // @[src/main/scala/tilelink/Broadcast.scala 129:48]
  wire  c_release = auto_in_c_bits_opcode == 3'h6; // @[src/main/scala/tilelink/Broadcast.scala 161:45]
  wire  releaseack_valid = auto_in_c_valid & c_release; // @[src/main/scala/tilelink/Broadcast.scala 192:79]
  wire [1:0] _readys_T = {d_normal_valid,releaseack_valid}; // @[src/main/scala/tilelink/Arbiter.scala 68:51]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[src/main/scala/tilelink/Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[src/main/scala/tilelink/Arbiter.scala 16:61]
  wire  readys__1 = _readys_T_7[1]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  reg  state__1; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  allowed__1 = idle ? readys__1 : state__1; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  d_normal_ready = auto_in_d_ready & allowed__1; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  wire  _T_13 = d_normal_ready & d_normal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] counter1 = counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  d_first = counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  line_508_clock;
  wire  line_508_reset;
  wire  line_508_valid;
  reg  line_508_valid_reg;
  wire [1:0] d_normal_bits_source = auto_out_d_bits_source[1:0]; // @[src/main/scala/tilelink/Broadcast.scala 121:26 130:21]
  wire  _d_trackerOH_T_1 = TLBroadcastTracker_io_need_d & TLBroadcastTracker_io_source == d_normal_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 123:62]
  wire  _d_trackerOH_T_3 = TLBroadcastTracker_1_io_need_d & TLBroadcastTracker_1_io_source == d_normal_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 123:62]
  wire  _d_trackerOH_T_5 = TLBroadcastTracker_2_io_need_d & TLBroadcastTracker_2_io_source == d_normal_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 123:62]
  wire  _d_trackerOH_T_7 = TLBroadcastTracker_3_io_need_d & TLBroadcastTracker_3_io_source == d_normal_bits_source; // @[src/main/scala/tilelink/Broadcast.scala 123:62]
  wire [3:0] _d_trackerOH_T_8 = {_d_trackerOH_T_7,_d_trackerOH_T_5,_d_trackerOH_T_3,_d_trackerOH_T_1}; // @[src/main/scala/tilelink/Broadcast.scala 123:102]
  reg [3:0] d_trackerOH_r; // @[src/main/scala/util/package.scala 80:63]
  wire  line_509_clock;
  wire  line_509_reset;
  wire  line_509_valid;
  reg  line_509_valid_reg;
  wire [3:0] _GEN_24 = d_first ? _d_trackerOH_T_8 : d_trackerOH_r; // @[src/main/scala/util/package.scala 80:{63,63,63}]
  wire  _T_20 = ~reset; // @[src/main/scala/tilelink/Broadcast.scala 125:14]
  wire  line_510_clock;
  wire  line_510_reset;
  wire  line_510_valid;
  reg  line_510_valid_reg;
  wire  _T_21 = ~(~auto_out_d_valid | _d_normal_valid_T_1 | auto_out_d_bits_opcode == 3'h0); // @[src/main/scala/tilelink/Broadcast.scala 125:14]
  wire  line_511_clock;
  wire  line_511_reset;
  wire  line_511_valid;
  reg  line_511_valid_reg;
  wire  nodeOut_d_ready = d_normal_ready | d_drop; // @[src/main/scala/tilelink/Broadcast.scala 128:50]
  wire  line_512_clock;
  wire  line_512_reset;
  wire  line_512_valid;
  reg  line_512_valid_reg;
  wire [1:0] _d_normal_bits_param_T_1 = d_what[0] ? 2'h0 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 133:51]
  wire [1:0] _d_normal_bits_param_T_2 = d_hasData ? _d_normal_bits_param_T_1 : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 133:36]
  wire [1:0] d_normal_bits_param = d_what[1] ? _d_normal_bits_param_T_2 : 2'h0; // @[src/main/scala/tilelink/Broadcast.scala 130:21 131:24 133:30]
  wire [1:0] d_mshr_hi = _GEN_24[3:2]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [1:0] d_mshr_lo = _GEN_24[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [1:0] _d_mshr_T_1 = d_mshr_hi | d_mshr_lo; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [1:0] d_mshr = {|d_mshr_hi,_d_mshr_T_1[1]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:10]
  wire  line_513_clock;
  wire  line_513_reset;
  wire  line_513_valid;
  reg  line_513_valid_reg;
  wire  _T_30 = ~(~d_normal_valid | (|_GEN_24 | d_normal_bits_opcode == 3'h6)); // @[src/main/scala/tilelink/Broadcast.scala 137:14]
  wire  line_514_clock;
  wire  line_514_reset;
  wire  line_514_valid;
  reg  line_514_valid_reg;
  wire  _T_39 = nodeOut_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  c_probeack = auto_in_c_bits_opcode == 3'h4; // @[src/main/scala/tilelink/Broadcast.scala 158:45]
  wire  c_probeackdata = auto_in_c_bits_opcode == 3'h5; // @[src/main/scala/tilelink/Broadcast.scala 159:45]
  wire  c_releasedata = auto_in_c_bits_opcode == 3'h7; // @[src/main/scala/tilelink/Broadcast.scala 160:45]
  wire  c_trackerOH_0 = TLBroadcastTracker_io_line == auto_in_c_bits_address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 162:55]
  wire  c_trackerOH_1 = TLBroadcastTracker_1_io_line == auto_in_c_bits_address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 162:55]
  wire  c_trackerOH_2 = TLBroadcastTracker_2_io_line == auto_in_c_bits_address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 162:55]
  wire  c_trackerOH_3 = TLBroadcastTracker_3_io_line == auto_in_c_bits_address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 162:55]
  wire [1:0] _c_trackerSrc_T = c_trackerOH_0 ? TLBroadcastTracker_io_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _c_trackerSrc_T_1 = c_trackerOH_1 ? TLBroadcastTracker_1_io_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _c_trackerSrc_T_2 = c_trackerOH_2 ? TLBroadcastTracker_2_io_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _c_trackerSrc_T_3 = c_trackerOH_3 ? TLBroadcastTracker_3_io_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _c_trackerSrc_T_4 = _c_trackerSrc_T | _c_trackerSrc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _c_trackerSrc_T_5 = _c_trackerSrc_T_4 | _c_trackerSrc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] c_trackerSrc = _c_trackerSrc_T_5 | _c_trackerSrc_T_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  readys__0 = _readys_T_7[0]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  reg  state__0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  allowed__0 = idle ? readys__0 : state__0; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  releaseack_ready = auto_in_d_ready & allowed__0; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  reg [1:0] beatsLeft_1; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
  wire  idle_1 = beatsLeft_1 == 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 61:28]
  wire  putfull_valid = auto_in_c_valid & (c_probeackdata | c_releasedata); // @[src/main/scala/tilelink/Broadcast.scala 197:35]
  wire [4:0] _readys_T_10 = {TLBroadcastTracker_3_io_out_a_valid,TLBroadcastTracker_2_io_out_a_valid,
    TLBroadcastTracker_1_io_out_a_valid,TLBroadcastTracker_io_out_a_valid,putfull_valid}; // @[src/main/scala/tilelink/Arbiter.scala 68:51]
  wire [5:0] _readys_T_11 = {_readys_T_10, 1'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [4:0] _readys_T_13 = _readys_T_10 | _readys_T_11[4:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [6:0] _readys_T_14 = {_readys_T_13, 2'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [4:0] _readys_T_16 = _readys_T_13 | _readys_T_14[4:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [8:0] _readys_T_17 = {_readys_T_16, 4'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [4:0] _readys_T_19 = _readys_T_16 | _readys_T_17[4:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [5:0] _readys_T_21 = {_readys_T_19, 1'h0}; // @[src/main/scala/tilelink/Arbiter.scala 16:78]
  wire [4:0] _readys_T_23 = ~_readys_T_21[4:0]; // @[src/main/scala/tilelink/Arbiter.scala 16:61]
  wire  readys_1_0 = _readys_T_23[0]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  reg  state_1_0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  allowed_1_0 = idle_1 ? readys_1_0 : state_1_0; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  putfull_ready = auto_out_a_ready & allowed_1_0; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  wire  _nodeIn_c_ready_T = c_release ? releaseack_ready : putfull_ready; // @[src/main/scala/tilelink/Broadcast.scala 184:38]
  wire  nodeIn_c_ready = c_probeack | _nodeIn_c_ready_T; // @[src/main/scala/tilelink/Broadcast.scala 184:32]
  wire  _clearOH_T = nodeIn_c_ready & auto_in_c_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _clearOH_T_1 = c_probeack | c_probeackdata; // @[src/main/scala/tilelink/Broadcast.scala 170:50]
  wire  _T_72 = auto_in_c_bits_param == 3'h4; // @[src/main/scala/tilelink/Broadcast.scala 178:27]
  wire  _T_73 = auto_in_c_bits_param == 3'h0 | _T_72; // @[src/main/scala/tilelink/Broadcast.scala 177:50]
  wire [11:0] _c_first_beats1_decode_T_1 = 12'h1f << auto_in_c_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _c_first_beats1_decode_T_3 = ~_c_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] c_first_beats1_decode = _c_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  line_515_clock;
  wire  line_515_reset;
  wire  line_515_valid;
  reg  line_515_valid_reg;
  wire [1:0] put_what = c_releasedata ? 2'h2 : 2'h1; // @[src/main/scala/tilelink/Broadcast.scala 195:25]
  wire [1:0] put_who = c_releasedata ? auto_in_c_bits_source : c_trackerSrc; // @[src/main/scala/tilelink/Broadcast.scala 196:25]
  wire [3:0] putfull_bits_a_source = {put_what,put_who}; // @[src/main/scala/tilelink/Broadcast.scala 198:38]
  wire [1:0] putfull_bits_a_mask_sizeOH_shiftAmount = auto_in_c_bits_size[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 64:49]
  wire [3:0] _putfull_bits_a_mask_sizeOH_T_1 = 4'h1 << putfull_bits_a_mask_sizeOH_shiftAmount; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire [2:0] putfull_bits_a_mask_sizeOH = _putfull_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[src/main/scala/util/Misc.scala 202:81]
  wire  _putfull_bits_a_mask_T = auto_in_c_bits_size >= 3'h3; // @[src/main/scala/util/Misc.scala 206:21]
  wire  putfull_bits_a_mask_size = putfull_bits_a_mask_sizeOH[2]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  putfull_bits_a_mask_bit = auto_in_c_bits_address[2]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  putfull_bits_a_mask_nbit = ~putfull_bits_a_mask_bit; // @[src/main/scala/util/Misc.scala 211:20]
  wire  putfull_bits_a_mask_acc = _putfull_bits_a_mask_T | putfull_bits_a_mask_size & putfull_bits_a_mask_nbit; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_acc_1 = _putfull_bits_a_mask_T | putfull_bits_a_mask_size & putfull_bits_a_mask_bit; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_size_1 = putfull_bits_a_mask_sizeOH[1]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  putfull_bits_a_mask_bit_1 = auto_in_c_bits_address[1]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  putfull_bits_a_mask_nbit_1 = ~putfull_bits_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 211:20]
  wire  putfull_bits_a_mask_eq_2 = putfull_bits_a_mask_nbit & putfull_bits_a_mask_nbit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_2 = putfull_bits_a_mask_acc | putfull_bits_a_mask_size_1 & putfull_bits_a_mask_eq_2; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_3 = putfull_bits_a_mask_nbit & putfull_bits_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_3 = putfull_bits_a_mask_acc | putfull_bits_a_mask_size_1 & putfull_bits_a_mask_eq_3; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_4 = putfull_bits_a_mask_bit & putfull_bits_a_mask_nbit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_4 = putfull_bits_a_mask_acc_1 | putfull_bits_a_mask_size_1 & putfull_bits_a_mask_eq_4; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_5 = putfull_bits_a_mask_bit & putfull_bits_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_5 = putfull_bits_a_mask_acc_1 | putfull_bits_a_mask_size_1 & putfull_bits_a_mask_eq_5; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_size_2 = putfull_bits_a_mask_sizeOH[0]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  putfull_bits_a_mask_bit_2 = auto_in_c_bits_address[0]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  putfull_bits_a_mask_nbit_2 = ~putfull_bits_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 211:20]
  wire  putfull_bits_a_mask_eq_6 = putfull_bits_a_mask_eq_2 & putfull_bits_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_6 = putfull_bits_a_mask_acc_2 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_6; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_7 = putfull_bits_a_mask_eq_2 & putfull_bits_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_7 = putfull_bits_a_mask_acc_2 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_7; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_8 = putfull_bits_a_mask_eq_3 & putfull_bits_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_8 = putfull_bits_a_mask_acc_3 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_8; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_9 = putfull_bits_a_mask_eq_3 & putfull_bits_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_9 = putfull_bits_a_mask_acc_3 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_9; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_10 = putfull_bits_a_mask_eq_4 & putfull_bits_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_10 = putfull_bits_a_mask_acc_4 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_10; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_11 = putfull_bits_a_mask_eq_4 & putfull_bits_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_11 = putfull_bits_a_mask_acc_4 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_11; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_12 = putfull_bits_a_mask_eq_5 & putfull_bits_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_12 = putfull_bits_a_mask_acc_5 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_12; // @[src/main/scala/util/Misc.scala 215:29]
  wire  putfull_bits_a_mask_eq_13 = putfull_bits_a_mask_eq_5 & putfull_bits_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  putfull_bits_a_mask_acc_13 = putfull_bits_a_mask_acc_5 | putfull_bits_a_mask_size_2 & putfull_bits_a_mask_eq_13; // @[src/main/scala/util/Misc.scala 215:29]
  wire [7:0] putfull_bits_a_mask = {putfull_bits_a_mask_acc_13,putfull_bits_a_mask_acc_12,putfull_bits_a_mask_acc_11,
    putfull_bits_a_mask_acc_10,putfull_bits_a_mask_acc_9,putfull_bits_a_mask_acc_8,putfull_bits_a_mask_acc_7,
    putfull_bits_a_mask_acc_6}; // @[src/main/scala/util/Misc.scala 222:10]
  wire  latch = idle & auto_in_d_ready; // @[src/main/scala/tilelink/Arbiter.scala 62:24]
  wire  winner__0 = readys__0 & releaseack_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner__1 = readys__1 & d_normal_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  _prefixOR_T = winner__0 | winner__1; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  line_516_clock;
  wire  line_516_reset;
  wire  line_516_valid;
  reg  line_516_valid_reg;
  wire  _T_122 = ~(~winner__0 | ~winner__1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
  wire  line_517_clock;
  wire  line_517_reset;
  wire  line_517_valid;
  reg  line_517_valid_reg;
  wire  _T_123 = releaseack_valid | d_normal_valid; // @[src/main/scala/tilelink/Arbiter.scala 79:31]
  wire  line_518_clock;
  wire  line_518_reset;
  wire  line_518_valid;
  reg  line_518_valid_reg;
  wire  _T_129 = ~(~(releaseack_valid | d_normal_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
  wire  line_519_clock;
  wire  line_519_reset;
  wire  line_519_valid;
  reg  line_519_valid_reg;
  wire  _nodeIn_d_valid_T_3 = state__0 & releaseack_valid | state__1 & d_normal_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  nodeIn_d_valid = idle ? _T_123 : _nodeIn_d_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  wire  _beatsLeft_T = auto_in_d_ready & nodeIn_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_37 = {{1'd0}, _beatsLeft_T}; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire [1:0] _beatsLeft_T_2 = beatsLeft - _GEN_37; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire  muxState__0 = idle ? winner__0 : state__0; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState__1 = idle ? winner__1 : state__1; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire [1:0] _nodeIn_d_bits_T_12 = muxState__0 ? auto_in_c_bits_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _nodeIn_d_bits_T_13 = muxState__1 ? d_normal_bits_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeIn_d_bits_T_15 = muxState__0 ? auto_in_c_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeIn_d_bits_T_16 = muxState__1 ? auto_out_d_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeIn_d_bits_T_21 = muxState__0 ? 3'h6 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeIn_d_bits_T_22 = muxState__1 ? d_normal_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [11:0] _decode_T_13 = 12'h1f << TLBroadcastTracker_io_out_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _decode_T_15 = ~_decode_T_13[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] decode_3 = _decode_T_15[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  opdata_3 = ~TLBroadcastTracker_io_out_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  wire [1:0] _T_131 = opdata_3 ? decode_3 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire [11:0] _decode_T_17 = 12'h1f << TLBroadcastTracker_1_io_out_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _decode_T_19 = ~_decode_T_17[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] decode_4 = _decode_T_19[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  opdata_4 = ~TLBroadcastTracker_1_io_out_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  wire [1:0] _T_132 = opdata_4 ? decode_4 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire [11:0] _decode_T_21 = 12'h1f << TLBroadcastTracker_2_io_out_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _decode_T_23 = ~_decode_T_21[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] decode_5 = _decode_T_23[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  opdata_5 = ~TLBroadcastTracker_2_io_out_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  wire [1:0] _T_133 = opdata_5 ? decode_5 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire [11:0] _decode_T_25 = 12'h1f << TLBroadcastTracker_3_io_out_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _decode_T_27 = ~_decode_T_25[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] decode_6 = _decode_T_27[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  opdata_6 = ~TLBroadcastTracker_3_io_out_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  wire [1:0] _T_134 = opdata_6 ? decode_6 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire  latch_1 = idle_1 & auto_out_a_ready; // @[src/main/scala/tilelink/Arbiter.scala 62:24]
  wire  readys_1_1 = _readys_T_23[1]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  readys_1_2 = _readys_T_23[2]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  readys_1_3 = _readys_T_23[3]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  readys_1_4 = _readys_T_23[4]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  winner_1_0 = readys_1_0 & putfull_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner_1_1 = readys_1_1 & TLBroadcastTracker_io_out_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner_1_2 = readys_1_2 & TLBroadcastTracker_1_io_out_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner_1_3 = readys_1_3 & TLBroadcastTracker_2_io_out_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner_1_4 = readys_1_4 & TLBroadcastTracker_3_io_out_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  prefixOR_2 = winner_1_0 | winner_1_1; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  prefixOR_3 = prefixOR_2 | winner_1_2; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  prefixOR_4 = prefixOR_3 | winner_1_3; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  _prefixOR_T_1 = prefixOR_4 | winner_1_4; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  line_520_clock;
  wire  line_520_reset;
  wire  line_520_valid;
  reg  line_520_valid_reg;
  wire  _T_156 = ~((~winner_1_0 | ~winner_1_1) & (~prefixOR_2 | ~winner_1_2) & (~prefixOR_3 | ~winner_1_3) & (~
    prefixOR_4 | ~winner_1_4)); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
  wire  line_521_clock;
  wire  line_521_reset;
  wire  line_521_valid;
  reg  line_521_valid_reg;
  wire  _T_160 = putfull_valid | TLBroadcastTracker_io_out_a_valid | TLBroadcastTracker_1_io_out_a_valid |
    TLBroadcastTracker_2_io_out_a_valid | TLBroadcastTracker_3_io_out_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 79:31]
  wire  line_522_clock;
  wire  line_522_reset;
  wire  line_522_valid;
  reg  line_522_valid_reg;
  wire  _T_169 = ~(~(putfull_valid | TLBroadcastTracker_io_out_a_valid | TLBroadcastTracker_1_io_out_a_valid |
    TLBroadcastTracker_2_io_out_a_valid | TLBroadcastTracker_3_io_out_a_valid) | _prefixOR_T_1); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
  wire  line_523_clock;
  wire  line_523_reset;
  wire  line_523_valid;
  reg  line_523_valid_reg;
  wire [1:0] maskedBeats_0_1 = winner_1_0 ? c_first_beats1_decode : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] maskedBeats_1_1 = winner_1_1 ? _T_131 : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] maskedBeats_2 = winner_1_2 ? _T_132 : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] maskedBeats_3 = winner_1_3 ? _T_133 : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] maskedBeats_4 = winner_1_4 ? _T_134 : 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 82:69]
  wire [1:0] _initBeats_T = maskedBeats_0_1 | maskedBeats_1_1; // @[src/main/scala/tilelink/Arbiter.scala 84:44]
  wire [1:0] _initBeats_T_1 = _initBeats_T | maskedBeats_2; // @[src/main/scala/tilelink/Arbiter.scala 84:44]
  wire [1:0] _initBeats_T_2 = _initBeats_T_1 | maskedBeats_3; // @[src/main/scala/tilelink/Arbiter.scala 84:44]
  wire [1:0] initBeats_1 = _initBeats_T_2 | maskedBeats_4; // @[src/main/scala/tilelink/Arbiter.scala 84:44]
  reg  state_1_1; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  reg  state_1_2; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  reg  state_1_3; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  reg  state_1_4; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  _nodeOut_a_valid_T_12 = state_1_0 & putfull_valid | state_1_1 & TLBroadcastTracker_io_out_a_valid | state_1_2 &
    TLBroadcastTracker_1_io_out_a_valid | state_1_3 & TLBroadcastTracker_2_io_out_a_valid | state_1_4 &
    TLBroadcastTracker_3_io_out_a_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  nodeOut_a_valid = idle_1 ? _T_160 : _nodeOut_a_valid_T_12; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  wire  _beatsLeft_T_4 = auto_out_a_ready & nodeOut_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_38 = {{1'd0}, _beatsLeft_T_4}; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire [1:0] _beatsLeft_T_6 = beatsLeft_1 - _GEN_38; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire  muxState_1_0 = idle_1 ? winner_1_0 : state_1_0; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState_1_1 = idle_1 ? winner_1_1 : state_1_1; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState_1_2 = idle_1 ? winner_1_2 : state_1_2; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState_1_3 = idle_1 ? winner_1_3 : state_1_3; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState_1_4 = idle_1 ? winner_1_4 : state_1_4; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  allowed_1_1 = idle_1 ? readys_1_1 : state_1_1; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  allowed_1_2 = idle_1 ? readys_1_2 : state_1_2; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  allowed_1_3 = idle_1 ? readys_1_3 : state_1_3; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  allowed_1_4 = idle_1 ? readys_1_4 : state_1_4; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire [63:0] _nodeOut_a_bits_T_9 = muxState_1_0 ? auto_in_c_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_10 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_11 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_12 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_13 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_14 = _nodeOut_a_bits_T_9 | _nodeOut_a_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_15 = _nodeOut_a_bits_T_14 | _nodeOut_a_bits_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _nodeOut_a_bits_T_16 = _nodeOut_a_bits_T_15 | _nodeOut_a_bits_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_18 = muxState_1_0 ? putfull_bits_a_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_19 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_20 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_21 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_22 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_23 = _nodeOut_a_bits_T_18 | _nodeOut_a_bits_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_24 = _nodeOut_a_bits_T_23 | _nodeOut_a_bits_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _nodeOut_a_bits_T_25 = _nodeOut_a_bits_T_24 | _nodeOut_a_bits_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_27 = muxState_1_0 ? auto_in_c_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_28 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_29 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_30 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_31 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_32 = _nodeOut_a_bits_T_27 | _nodeOut_a_bits_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_33 = _nodeOut_a_bits_T_32 | _nodeOut_a_bits_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _nodeOut_a_bits_T_34 = _nodeOut_a_bits_T_33 | _nodeOut_a_bits_T_30; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_36 = muxState_1_0 ? putfull_bits_a_source : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_37 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_source : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_38 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_source : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_39 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_source : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_40 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_source : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_41 = _nodeOut_a_bits_T_36 | _nodeOut_a_bits_T_37; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_42 = _nodeOut_a_bits_T_41 | _nodeOut_a_bits_T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _nodeOut_a_bits_T_43 = _nodeOut_a_bits_T_42 | _nodeOut_a_bits_T_39; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_45 = muxState_1_0 ? auto_in_c_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_46 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_47 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_48 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_49 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_50 = _nodeOut_a_bits_T_45 | _nodeOut_a_bits_T_46; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_51 = _nodeOut_a_bits_T_50 | _nodeOut_a_bits_T_47; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_52 = _nodeOut_a_bits_T_51 | _nodeOut_a_bits_T_48; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_64 = muxState_1_1 ? TLBroadcastTracker_io_out_a_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_65 = muxState_1_2 ? TLBroadcastTracker_1_io_out_a_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_66 = muxState_1_3 ? TLBroadcastTracker_2_io_out_a_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_67 = muxState_1_4 ? TLBroadcastTracker_3_io_out_a_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_69 = _nodeOut_a_bits_T_64 | _nodeOut_a_bits_T_65; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _nodeOut_a_bits_T_70 = _nodeOut_a_bits_T_69 | _nodeOut_a_bits_T_66; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  probe_todo; // @[src/main/scala/tilelink/Broadcast.scala 215:31]
  reg [26:0] probe_line; // @[src/main/scala/tilelink/Broadcast.scala 216:27]
  reg [1:0] probe_perms; // @[src/main/scala/tilelink/Broadcast.scala 217:28]
  wire [1:0] _probe_next_T_1 = {probe_todo, 1'h0}; // @[src/main/scala/tilelink/Broadcast.scala 218:58]
  wire [1:0] _probe_next_T_2 = ~_probe_next_T_1; // @[src/main/scala/tilelink/Broadcast.scala 218:37]
  wire [1:0] _GEN_39 = {{1'd0}, probe_todo}; // @[src/main/scala/tilelink/Broadcast.scala 218:35]
  wire [1:0] probe_next = _GEN_39 & _probe_next_T_2; // @[src/main/scala/tilelink/Broadcast.scala 218:35]
  wire  probe_busy = |probe_todo; // @[src/main/scala/tilelink/Broadcast.scala 219:35]
  wire  _T_174 = auto_in_b_ready & probe_busy; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_524_clock;
  wire  line_524_reset;
  wire  line_524_valid;
  reg  line_524_valid_reg;
  wire [1:0] _probe_todo_T = ~probe_next; // @[src/main/scala/tilelink/Broadcast.scala 227:53]
  wire [1:0] _probe_todo_T_1 = _GEN_39 & _probe_todo_T; // @[src/main/scala/tilelink/Broadcast.scala 227:51]
  wire [1:0] _GEN_28 = _T_174 ? _probe_todo_T_1 : {{1'd0}, probe_todo}; // @[src/main/scala/tilelink/Broadcast.scala 227:24 215:31 227:37]
  reg [1:0] a_first_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire  a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  _nodeIn_a_ready_T_1 = ~a_first | filter_io_request_ready; // @[src/main/scala/tilelink/Broadcast.scala 243:31]
  wire [3:0] matchTrackers = {TLBroadcastTracker_3_io_line == auto_in_a_bits_address[31:5],TLBroadcastTracker_2_io_line
     == auto_in_a_bits_address[31:5],TLBroadcastTracker_1_io_line == auto_in_a_bits_address[31:5],
    TLBroadcastTracker_io_line == auto_in_a_bits_address[31:5]}; // @[src/main/scala/tilelink/Broadcast.scala 236:100]
  wire  matchTracker = |matchTrackers; // @[src/main/scala/tilelink/Broadcast.scala 237:40]
  wire  _freeTrackers_WIRE_3 = TLBroadcastTracker_3_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 234:{33,33}]
  wire  _freeTrackers_WIRE_2 = TLBroadcastTracker_2_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 234:{33,33}]
  wire  _freeTrackers_WIRE_1 = TLBroadcastTracker_1_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 234:{33,33}]
  wire  _freeTrackers_WIRE_0 = TLBroadcastTracker_io_idle; // @[src/main/scala/tilelink/Broadcast.scala 234:{33,33}]
  wire [3:0] freeTrackers = {_freeTrackers_WIRE_3,_freeTrackers_WIRE_2,_freeTrackers_WIRE_1,_freeTrackers_WIRE_0}; // @[src/main/scala/tilelink/Broadcast.scala 234:64]
  wire [4:0] _allocTracker_T = {freeTrackers, 1'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [3:0] _allocTracker_T_2 = freeTrackers | _allocTracker_T[3:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [5:0] _allocTracker_T_3 = {_allocTracker_T_2, 2'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [3:0] _allocTracker_T_5 = _allocTracker_T_2 | _allocTracker_T_3[3:0]; // @[src/main/scala/util/package.scala 245:43]
  wire [4:0] _allocTracker_T_7 = {_allocTracker_T_5, 1'h0}; // @[src/main/scala/tilelink/Broadcast.scala 238:64]
  wire [4:0] _allocTracker_T_8 = ~_allocTracker_T_7; // @[src/main/scala/tilelink/Broadcast.scala 238:41]
  wire [4:0] _GEN_41 = {{1'd0}, freeTrackers}; // @[src/main/scala/tilelink/Broadcast.scala 238:39]
  wire [4:0] allocTracker = _GEN_41 & _allocTracker_T_8; // @[src/main/scala/tilelink/Broadcast.scala 238:39]
  wire [4:0] selectTracker = matchTracker ? {{1'd0}, matchTrackers} : allocTracker; // @[src/main/scala/tilelink/Broadcast.scala 239:30]
  wire  _trackerReadys_WIRE_3 = TLBroadcastTracker_3_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 240:{34,34}]
  wire  _trackerReadys_WIRE_2 = TLBroadcastTracker_2_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 240:{34,34}]
  wire  _trackerReadys_WIRE_1 = TLBroadcastTracker_1_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 240:{34,34}]
  wire  _trackerReadys_WIRE_0 = TLBroadcastTracker_io_in_a_ready; // @[src/main/scala/tilelink/Broadcast.scala 240:{34,34}]
  wire [3:0] trackerReadys = {_trackerReadys_WIRE_3,_trackerReadys_WIRE_2,_trackerReadys_WIRE_1,_trackerReadys_WIRE_0}; // @[src/main/scala/tilelink/Broadcast.scala 240:63]
  wire [4:0] _GEN_42 = {{1'd0}, trackerReadys}; // @[src/main/scala/tilelink/Broadcast.scala 241:41]
  wire [4:0] _trackerReady_T = selectTracker & _GEN_42; // @[src/main/scala/tilelink/Broadcast.scala 241:41]
  wire  trackerReady = |_trackerReady_T; // @[src/main/scala/tilelink/Broadcast.scala 241:58]
  wire  nodeIn_a_ready = (~a_first | filter_io_request_ready) & trackerReady; // @[src/main/scala/tilelink/Broadcast.scala 243:59]
  wire  _a_first_T = nodeIn_a_ready & auto_in_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [11:0] _a_first_beats1_decode_T_1 = 12'h1f << auto_in_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _a_first_beats1_decode_T_3 = ~_a_first_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] a_first_beats1_decode = _a_first_beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  a_first_beats1_opdata = ~auto_in_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  wire [1:0] a_first_counter1 = a_first_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  line_525_clock;
  wire  line_525_reset;
  wire  line_525_valid;
  reg  line_525_valid_reg;
  wire [3:0] filter_io_request_bits_mshr_lo = selectTracker[3:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [3:0] _GEN_43 = {{3'd0}, selectTracker[4]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [3:0] _filter_io_request_bits_mshr_T_1 = _GEN_43 | filter_io_request_bits_mshr_lo; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [1:0] filter_io_request_bits_mshr_hi_1 = _filter_io_request_bits_mshr_T_1[3:2]; // @[src/main/scala/chisel3/util/OneHot.scala 30:18]
  wire [1:0] filter_io_request_bits_mshr_lo_1 = _filter_io_request_bits_mshr_T_1[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 31:18]
  wire [1:0] _filter_io_request_bits_mshr_T_3 = filter_io_request_bits_mshr_hi_1 | filter_io_request_bits_mshr_lo_1; // @[src/main/scala/chisel3/util/OneHot.scala 32:28]
  wire [2:0] _filter_io_request_bits_mshr_T_6 = {|selectTracker[4],|filter_io_request_bits_mshr_hi_1,
    _filter_io_request_bits_mshr_T_3[1]}; // @[src/main/scala/chisel3/util/OneHot.scala 32:10]
  wire  _filter_io_request_bits_needT_acq_needT_T_2 = 3'h1 == auto_in_a_bits_param; // @[src/main/scala/tilelink/Edges.scala 276:70]
  wire  filter_io_request_bits_needT_acq_needT = 3'h2 == auto_in_a_bits_param | 3'h1 == auto_in_a_bits_param; // @[src/main/scala/tilelink/Edges.scala 276:70]
  wire  _filter_io_request_bits_needT_T_11 = 3'h4 == auto_in_a_bits_opcode ? 1'h0 : 1'h1; // @[src/main/scala/tilelink/Edges.scala 280:55]
  wire  _filter_io_request_bits_needT_T_13 = 3'h5 == auto_in_a_bits_opcode ? _filter_io_request_bits_needT_acq_needT_T_2
     : _filter_io_request_bits_needT_T_11; // @[src/main/scala/tilelink/Edges.scala 280:55]
  wire  _filter_io_request_bits_needT_T_15 = 3'h6 == auto_in_a_bits_opcode ? filter_io_request_bits_needT_acq_needT :
    _filter_io_request_bits_needT_T_13; // @[src/main/scala/tilelink/Edges.scala 280:55]
  wire  others = ~filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 257:54]
  wire  _T_196 = filter_io_response_ready & filter_io_response_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_526_clock;
  wire  line_526_reset;
  wire  line_526_valid;
  reg  line_526_valid_reg;
  wire [1:0] _GEN_30 = _T_196 ? {{1'd0}, others} : _GEN_28; // @[src/main/scala/tilelink/Broadcast.scala 260:38 261:21]
  wire [1:0] responseMSHR_shiftAmount = filter_io_response_bits_mshr; // @[src/main/scala/chisel3/util/OneHot.scala 64:49]
  wire [3:0] _responseMSHR_T = 4'h1 << responseMSHR_shiftAmount; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  responseMSHR_0 = _responseMSHR_T[0]; // @[src/main/scala/tilelink/Broadcast.scala 269:85]
  wire  responseMSHR_1 = _responseMSHR_T[1]; // @[src/main/scala/tilelink/Broadcast.scala 269:85]
  wire  responseMSHR_2 = _responseMSHR_T[2]; // @[src/main/scala/tilelink/Broadcast.scala 269:85]
  wire  responseMSHR_3 = _responseMSHR_T[3]; // @[src/main/scala/tilelink/Broadcast.scala 269:85]
  wire [1:0] _GEN_44 = reset ? 2'h0 : _GEN_30; // @[src/main/scala/tilelink/Broadcast.scala 215:{31,31}]
  BroadcastFilter filter ( // @[src/main/scala/tilelink/Broadcast.scala 99:26]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_request_ready(filter_io_request_ready),
    .io_request_valid(filter_io_request_valid),
    .io_request_bits_mshr(filter_io_request_bits_mshr),
    .io_request_bits_address(filter_io_request_bits_address),
    .io_request_bits_allocOH(filter_io_request_bits_allocOH),
    .io_request_bits_needT(filter_io_request_bits_needT),
    .io_response_ready(filter_io_response_ready),
    .io_response_valid(filter_io_response_valid),
    .io_response_bits_mshr(filter_io_response_bits_mshr),
    .io_response_bits_address(filter_io_response_bits_address),
    .io_response_bits_allocOH(filter_io_response_bits_allocOH),
    .io_response_bits_needT(filter_io_response_bits_needT)
  );
  TLBroadcastTracker TLBroadcastTracker ( // @[src/main/scala/tilelink/Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_clock),
    .reset(TLBroadcastTracker_reset),
    .io_in_a_first(TLBroadcastTracker_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_io_in_a_bits_address),
    .io_in_a_bits_mask(TLBroadcastTracker_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_io_out_a_bits_address),
    .io_out_a_bits_mask(TLBroadcastTracker_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_io_out_a_bits_data),
    .io_probe_valid(TLBroadcastTracker_io_probe_valid),
    .io_probe_bits_count(TLBroadcastTracker_io_probe_bits_count),
    .io_probenack(TLBroadcastTracker_io_probenack),
    .io_probedack(TLBroadcastTracker_io_probedack),
    .io_probesack(TLBroadcastTracker_io_probesack),
    .io_d_last(TLBroadcastTracker_io_d_last),
    .io_e_last(TLBroadcastTracker_io_e_last),
    .io_source(TLBroadcastTracker_io_source),
    .io_line(TLBroadcastTracker_io_line),
    .io_idle(TLBroadcastTracker_io_idle),
    .io_need_d(TLBroadcastTracker_io_need_d)
  );
  TLBroadcastTracker_1 TLBroadcastTracker_1 ( // @[src/main/scala/tilelink/Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_1_clock),
    .reset(TLBroadcastTracker_1_reset),
    .io_in_a_first(TLBroadcastTracker_1_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_1_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_1_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_1_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_1_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_1_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_1_io_in_a_bits_address),
    .io_in_a_bits_mask(TLBroadcastTracker_1_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_1_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_1_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_1_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_1_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_1_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_1_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_1_io_out_a_bits_address),
    .io_out_a_bits_mask(TLBroadcastTracker_1_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_1_io_out_a_bits_data),
    .io_probe_valid(TLBroadcastTracker_1_io_probe_valid),
    .io_probe_bits_count(TLBroadcastTracker_1_io_probe_bits_count),
    .io_probenack(TLBroadcastTracker_1_io_probenack),
    .io_probedack(TLBroadcastTracker_1_io_probedack),
    .io_probesack(TLBroadcastTracker_1_io_probesack),
    .io_d_last(TLBroadcastTracker_1_io_d_last),
    .io_e_last(TLBroadcastTracker_1_io_e_last),
    .io_source(TLBroadcastTracker_1_io_source),
    .io_line(TLBroadcastTracker_1_io_line),
    .io_idle(TLBroadcastTracker_1_io_idle),
    .io_need_d(TLBroadcastTracker_1_io_need_d)
  );
  TLBroadcastTracker_2 TLBroadcastTracker_2 ( // @[src/main/scala/tilelink/Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_2_clock),
    .reset(TLBroadcastTracker_2_reset),
    .io_in_a_first(TLBroadcastTracker_2_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_2_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_2_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_2_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_2_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_2_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_2_io_in_a_bits_address),
    .io_in_a_bits_mask(TLBroadcastTracker_2_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_2_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_2_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_2_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_2_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_2_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_2_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_2_io_out_a_bits_address),
    .io_out_a_bits_mask(TLBroadcastTracker_2_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_2_io_out_a_bits_data),
    .io_probe_valid(TLBroadcastTracker_2_io_probe_valid),
    .io_probe_bits_count(TLBroadcastTracker_2_io_probe_bits_count),
    .io_probenack(TLBroadcastTracker_2_io_probenack),
    .io_probedack(TLBroadcastTracker_2_io_probedack),
    .io_probesack(TLBroadcastTracker_2_io_probesack),
    .io_d_last(TLBroadcastTracker_2_io_d_last),
    .io_e_last(TLBroadcastTracker_2_io_e_last),
    .io_source(TLBroadcastTracker_2_io_source),
    .io_line(TLBroadcastTracker_2_io_line),
    .io_idle(TLBroadcastTracker_2_io_idle),
    .io_need_d(TLBroadcastTracker_2_io_need_d)
  );
  TLBroadcastTracker_3 TLBroadcastTracker_3 ( // @[src/main/scala/tilelink/Broadcast.scala 107:15]
    .clock(TLBroadcastTracker_3_clock),
    .reset(TLBroadcastTracker_3_reset),
    .io_in_a_first(TLBroadcastTracker_3_io_in_a_first),
    .io_in_a_ready(TLBroadcastTracker_3_io_in_a_ready),
    .io_in_a_valid(TLBroadcastTracker_3_io_in_a_valid),
    .io_in_a_bits_opcode(TLBroadcastTracker_3_io_in_a_bits_opcode),
    .io_in_a_bits_size(TLBroadcastTracker_3_io_in_a_bits_size),
    .io_in_a_bits_source(TLBroadcastTracker_3_io_in_a_bits_source),
    .io_in_a_bits_address(TLBroadcastTracker_3_io_in_a_bits_address),
    .io_in_a_bits_mask(TLBroadcastTracker_3_io_in_a_bits_mask),
    .io_in_a_bits_data(TLBroadcastTracker_3_io_in_a_bits_data),
    .io_out_a_ready(TLBroadcastTracker_3_io_out_a_ready),
    .io_out_a_valid(TLBroadcastTracker_3_io_out_a_valid),
    .io_out_a_bits_opcode(TLBroadcastTracker_3_io_out_a_bits_opcode),
    .io_out_a_bits_size(TLBroadcastTracker_3_io_out_a_bits_size),
    .io_out_a_bits_source(TLBroadcastTracker_3_io_out_a_bits_source),
    .io_out_a_bits_address(TLBroadcastTracker_3_io_out_a_bits_address),
    .io_out_a_bits_mask(TLBroadcastTracker_3_io_out_a_bits_mask),
    .io_out_a_bits_data(TLBroadcastTracker_3_io_out_a_bits_data),
    .io_probe_valid(TLBroadcastTracker_3_io_probe_valid),
    .io_probe_bits_count(TLBroadcastTracker_3_io_probe_bits_count),
    .io_probenack(TLBroadcastTracker_3_io_probenack),
    .io_probedack(TLBroadcastTracker_3_io_probedack),
    .io_probesack(TLBroadcastTracker_3_io_probesack),
    .io_d_last(TLBroadcastTracker_3_io_d_last),
    .io_e_last(TLBroadcastTracker_3_io_e_last),
    .io_source(TLBroadcastTracker_3_io_source),
    .io_line(TLBroadcastTracker_3_io_line),
    .io_idle(TLBroadcastTracker_3_io_idle),
    .io_need_d(TLBroadcastTracker_3_io_need_d)
  );
  GEN_w1_line #(.COVER_INDEX(508)) line_508 (
    .clock(line_508_clock),
    .reset(line_508_reset),
    .valid(line_508_valid)
  );
  GEN_w1_line #(.COVER_INDEX(509)) line_509 (
    .clock(line_509_clock),
    .reset(line_509_reset),
    .valid(line_509_valid)
  );
  GEN_w1_line #(.COVER_INDEX(510)) line_510 (
    .clock(line_510_clock),
    .reset(line_510_reset),
    .valid(line_510_valid)
  );
  GEN_w1_line #(.COVER_INDEX(511)) line_511 (
    .clock(line_511_clock),
    .reset(line_511_reset),
    .valid(line_511_valid)
  );
  GEN_w1_line #(.COVER_INDEX(512)) line_512 (
    .clock(line_512_clock),
    .reset(line_512_reset),
    .valid(line_512_valid)
  );
  GEN_w1_line #(.COVER_INDEX(513)) line_513 (
    .clock(line_513_clock),
    .reset(line_513_reset),
    .valid(line_513_valid)
  );
  GEN_w1_line #(.COVER_INDEX(514)) line_514 (
    .clock(line_514_clock),
    .reset(line_514_reset),
    .valid(line_514_valid)
  );
  GEN_w1_line #(.COVER_INDEX(515)) line_515 (
    .clock(line_515_clock),
    .reset(line_515_reset),
    .valid(line_515_valid)
  );
  GEN_w1_line #(.COVER_INDEX(516)) line_516 (
    .clock(line_516_clock),
    .reset(line_516_reset),
    .valid(line_516_valid)
  );
  GEN_w1_line #(.COVER_INDEX(517)) line_517 (
    .clock(line_517_clock),
    .reset(line_517_reset),
    .valid(line_517_valid)
  );
  GEN_w1_line #(.COVER_INDEX(518)) line_518 (
    .clock(line_518_clock),
    .reset(line_518_reset),
    .valid(line_518_valid)
  );
  GEN_w1_line #(.COVER_INDEX(519)) line_519 (
    .clock(line_519_clock),
    .reset(line_519_reset),
    .valid(line_519_valid)
  );
  GEN_w1_line #(.COVER_INDEX(520)) line_520 (
    .clock(line_520_clock),
    .reset(line_520_reset),
    .valid(line_520_valid)
  );
  GEN_w1_line #(.COVER_INDEX(521)) line_521 (
    .clock(line_521_clock),
    .reset(line_521_reset),
    .valid(line_521_valid)
  );
  GEN_w1_line #(.COVER_INDEX(522)) line_522 (
    .clock(line_522_clock),
    .reset(line_522_reset),
    .valid(line_522_valid)
  );
  GEN_w1_line #(.COVER_INDEX(523)) line_523 (
    .clock(line_523_clock),
    .reset(line_523_reset),
    .valid(line_523_valid)
  );
  GEN_w1_line #(.COVER_INDEX(524)) line_524 (
    .clock(line_524_clock),
    .reset(line_524_reset),
    .valid(line_524_valid)
  );
  GEN_w1_line #(.COVER_INDEX(525)) line_525 (
    .clock(line_525_clock),
    .reset(line_525_reset),
    .valid(line_525_valid)
  );
  GEN_w1_line #(.COVER_INDEX(526)) line_526 (
    .clock(line_526_clock),
    .reset(line_526_reset),
    .valid(line_526_valid)
  );
  assign line_508_clock = clock;
  assign line_508_reset = reset;
  assign line_508_valid = _T_13 ^ line_508_valid_reg;
  assign line_509_clock = clock;
  assign line_509_reset = reset;
  assign line_509_valid = d_first ^ line_509_valid_reg;
  assign line_510_clock = clock;
  assign line_510_reset = reset;
  assign line_510_valid = _T_20 ^ line_510_valid_reg;
  assign line_511_clock = clock;
  assign line_511_reset = reset;
  assign line_511_valid = _T_21 ^ line_511_valid_reg;
  assign line_512_clock = clock;
  assign line_512_reset = reset;
  assign line_512_valid = d_what[1] ^ line_512_valid_reg;
  assign line_513_clock = clock;
  assign line_513_reset = reset;
  assign line_513_valid = _T_20 ^ line_513_valid_reg;
  assign line_514_clock = clock;
  assign line_514_reset = reset;
  assign line_514_valid = _T_30 ^ line_514_valid_reg;
  assign line_515_clock = clock;
  assign line_515_reset = reset;
  assign line_515_valid = _clearOH_T ^ line_515_valid_reg;
  assign line_516_clock = clock;
  assign line_516_reset = reset;
  assign line_516_valid = _T_20 ^ line_516_valid_reg;
  assign line_517_clock = clock;
  assign line_517_reset = reset;
  assign line_517_valid = _T_122 ^ line_517_valid_reg;
  assign line_518_clock = clock;
  assign line_518_reset = reset;
  assign line_518_valid = _T_20 ^ line_518_valid_reg;
  assign line_519_clock = clock;
  assign line_519_reset = reset;
  assign line_519_valid = _T_129 ^ line_519_valid_reg;
  assign line_520_clock = clock;
  assign line_520_reset = reset;
  assign line_520_valid = _T_20 ^ line_520_valid_reg;
  assign line_521_clock = clock;
  assign line_521_reset = reset;
  assign line_521_valid = _T_156 ^ line_521_valid_reg;
  assign line_522_clock = clock;
  assign line_522_reset = reset;
  assign line_522_valid = _T_20 ^ line_522_valid_reg;
  assign line_523_clock = clock;
  assign line_523_reset = reset;
  assign line_523_valid = _T_169 ^ line_523_valid_reg;
  assign line_524_clock = clock;
  assign line_524_reset = reset;
  assign line_524_valid = _T_174 ^ line_524_valid_reg;
  assign line_525_clock = clock;
  assign line_525_reset = reset;
  assign line_525_valid = _a_first_T ^ line_525_valid_reg;
  assign line_526_clock = clock;
  assign line_526_reset = reset;
  assign line_526_valid = _T_196 ^ line_526_valid_reg;
  assign auto_in_a_ready = (~a_first | filter_io_request_ready) & trackerReady; // @[src/main/scala/tilelink/Broadcast.scala 243:59]
  assign auto_in_b_valid = |probe_todo; // @[src/main/scala/tilelink/Broadcast.scala 219:35]
  assign auto_in_b_bits_param = probe_perms; // @[src/main/scala/tilelink/Edges.scala 631:17 633:15]
  assign auto_in_b_bits_address = {probe_line, 5'h0}; // @[src/main/scala/tilelink/Broadcast.scala 225:46]
  assign auto_in_c_ready = c_probeack | _nodeIn_c_ready_T; // @[src/main/scala/tilelink/Broadcast.scala 184:32]
  assign auto_in_d_valid = idle ? _T_123 : _nodeIn_d_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  assign auto_in_d_bits_opcode = _nodeIn_d_bits_T_21 | _nodeIn_d_bits_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_param = muxState__1 ? d_normal_bits_param : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_size = _nodeIn_d_bits_T_15 | _nodeIn_d_bits_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_source = _nodeIn_d_bits_T_12 | _nodeIn_d_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_sink = muxState__1 ? d_mshr : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_denied = muxState__1 & auto_out_d_bits_denied; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_data = muxState__1 ? auto_out_d_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_in_d_bits_corrupt = muxState__1 & auto_out_d_bits_corrupt; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_valid = idle_1 ? _T_160 : _nodeOut_a_valid_T_12; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  assign auto_out_a_bits_opcode = _nodeOut_a_bits_T_70 | _nodeOut_a_bits_T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_size = _nodeOut_a_bits_T_52 | _nodeOut_a_bits_T_49; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_source = _nodeOut_a_bits_T_43 | _nodeOut_a_bits_T_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_address = _nodeOut_a_bits_T_34 | _nodeOut_a_bits_T_31; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_mask = _nodeOut_a_bits_T_25 | _nodeOut_a_bits_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_data = _nodeOut_a_bits_T_16 | _nodeOut_a_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_d_ready = d_normal_ready | d_drop; // @[src/main/scala/tilelink/Broadcast.scala 128:50]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_request_valid = auto_in_a_valid & a_first & trackerReady; // @[src/main/scala/tilelink/Broadcast.scala 250:56]
  assign filter_io_request_bits_mshr = _filter_io_request_bits_mshr_T_6[1:0]; // @[src/main/scala/tilelink/Broadcast.scala 251:38]
  assign filter_io_request_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign filter_io_request_bits_allocOH = auto_in_a_bits_source == 2'h0; // @[src/main/scala/diplomacy/Parameters.scala 46:9]
  assign filter_io_request_bits_needT = 3'h7 == auto_in_a_bits_opcode ? filter_io_request_bits_needT_acq_needT :
    _filter_io_request_bits_needT_T_15; // @[src/main/scala/tilelink/Edges.scala 280:55]
  assign filter_io_response_ready = ~probe_busy; // @[src/main/scala/tilelink/Broadcast.scala 259:35]
  assign TLBroadcastTracker_clock = clock;
  assign TLBroadcastTracker_reset = reset;
  assign TLBroadcastTracker_io_in_a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  assign TLBroadcastTracker_io_in_a_valid = auto_in_a_valid & selectTracker[0] & _nodeIn_a_ready_T_1; // @[src/main/scala/tilelink/Broadcast.scala 245:46]
  assign TLBroadcastTracker_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_in_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_in_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_in_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_in_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_in_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_io_out_a_ready = auto_out_a_ready & allowed_1_1; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign TLBroadcastTracker_io_probe_valid = _T_196 & responseMSHR_0; // @[src/main/scala/tilelink/Broadcast.scala 272:56]
  assign TLBroadcastTracker_io_probe_bits_count = ~filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 257:54]
  assign TLBroadcastTracker_io_probenack = _clearOH_T & c_probeack & c_trackerOH_0; // @[src/main/scala/tilelink/Broadcast.scala 175:54]
  assign TLBroadcastTracker_io_probedack = _GEN_24[0] & _T_39 & d_drop; // @[src/main/scala/tilelink/Broadcast.scala 143:51]
  assign TLBroadcastTracker_io_probesack = _clearOH_T & c_trackerOH_0 & _clearOH_T_1 & _T_73; // @[src/main/scala/tilelink/Broadcast.scala 176:84]
  assign TLBroadcastTracker_io_d_last = _GEN_24[0] & _T_13 & d_response & d_last; // @[src/main/scala/tilelink/Broadcast.scala 142:65]
  assign TLBroadcastTracker_io_e_last = _T[0] & auto_in_e_valid; // @[src/main/scala/tilelink/Broadcast.scala 113:34]
  assign TLBroadcastTracker_1_clock = clock;
  assign TLBroadcastTracker_1_reset = reset;
  assign TLBroadcastTracker_1_io_in_a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  assign TLBroadcastTracker_1_io_in_a_valid = auto_in_a_valid & selectTracker[1] & _nodeIn_a_ready_T_1; // @[src/main/scala/tilelink/Broadcast.scala 245:46]
  assign TLBroadcastTracker_1_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_in_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_in_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_in_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_in_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_in_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_1_io_out_a_ready = auto_out_a_ready & allowed_1_2; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign TLBroadcastTracker_1_io_probe_valid = _T_196 & responseMSHR_1; // @[src/main/scala/tilelink/Broadcast.scala 272:56]
  assign TLBroadcastTracker_1_io_probe_bits_count = ~filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 257:54]
  assign TLBroadcastTracker_1_io_probenack = _clearOH_T & c_probeack & c_trackerOH_1; // @[src/main/scala/tilelink/Broadcast.scala 175:54]
  assign TLBroadcastTracker_1_io_probedack = _GEN_24[1] & _T_39 & d_drop; // @[src/main/scala/tilelink/Broadcast.scala 143:51]
  assign TLBroadcastTracker_1_io_probesack = _clearOH_T & c_trackerOH_1 & _clearOH_T_1 & _T_73; // @[src/main/scala/tilelink/Broadcast.scala 176:84]
  assign TLBroadcastTracker_1_io_d_last = _GEN_24[1] & _T_13 & d_response & d_last; // @[src/main/scala/tilelink/Broadcast.scala 142:65]
  assign TLBroadcastTracker_1_io_e_last = _T[1] & auto_in_e_valid; // @[src/main/scala/tilelink/Broadcast.scala 113:34]
  assign TLBroadcastTracker_2_clock = clock;
  assign TLBroadcastTracker_2_reset = reset;
  assign TLBroadcastTracker_2_io_in_a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  assign TLBroadcastTracker_2_io_in_a_valid = auto_in_a_valid & selectTracker[2] & _nodeIn_a_ready_T_1; // @[src/main/scala/tilelink/Broadcast.scala 245:46]
  assign TLBroadcastTracker_2_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_in_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_in_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_in_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_in_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_in_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_2_io_out_a_ready = auto_out_a_ready & allowed_1_3; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign TLBroadcastTracker_2_io_probe_valid = _T_196 & responseMSHR_2; // @[src/main/scala/tilelink/Broadcast.scala 272:56]
  assign TLBroadcastTracker_2_io_probe_bits_count = ~filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 257:54]
  assign TLBroadcastTracker_2_io_probenack = _clearOH_T & c_probeack & c_trackerOH_2; // @[src/main/scala/tilelink/Broadcast.scala 175:54]
  assign TLBroadcastTracker_2_io_probedack = _GEN_24[2] & _T_39 & d_drop; // @[src/main/scala/tilelink/Broadcast.scala 143:51]
  assign TLBroadcastTracker_2_io_probesack = _clearOH_T & c_trackerOH_2 & _clearOH_T_1 & _T_73; // @[src/main/scala/tilelink/Broadcast.scala 176:84]
  assign TLBroadcastTracker_2_io_d_last = _GEN_24[2] & _T_13 & d_response & d_last; // @[src/main/scala/tilelink/Broadcast.scala 142:65]
  assign TLBroadcastTracker_2_io_e_last = _T[2] & auto_in_e_valid; // @[src/main/scala/tilelink/Broadcast.scala 113:34]
  assign TLBroadcastTracker_3_clock = clock;
  assign TLBroadcastTracker_3_reset = reset;
  assign TLBroadcastTracker_3_io_in_a_first = a_first_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  assign TLBroadcastTracker_3_io_in_a_valid = auto_in_a_valid & selectTracker[3] & _nodeIn_a_ready_T_1; // @[src/main/scala/tilelink/Broadcast.scala 245:46]
  assign TLBroadcastTracker_3_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_in_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_in_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_in_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_in_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_in_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign TLBroadcastTracker_3_io_out_a_ready = auto_out_a_ready & allowed_1_4; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign TLBroadcastTracker_3_io_probe_valid = _T_196 & responseMSHR_3; // @[src/main/scala/tilelink/Broadcast.scala 272:56]
  assign TLBroadcastTracker_3_io_probe_bits_count = ~filter_io_response_bits_allocOH; // @[src/main/scala/tilelink/Broadcast.scala 257:54]
  assign TLBroadcastTracker_3_io_probenack = _clearOH_T & c_probeack & c_trackerOH_3; // @[src/main/scala/tilelink/Broadcast.scala 175:54]
  assign TLBroadcastTracker_3_io_probedack = _GEN_24[3] & _T_39 & d_drop; // @[src/main/scala/tilelink/Broadcast.scala 143:51]
  assign TLBroadcastTracker_3_io_probesack = _clearOH_T & c_trackerOH_3 & _clearOH_T_1 & _T_73; // @[src/main/scala/tilelink/Broadcast.scala 176:84]
  assign TLBroadcastTracker_3_io_d_last = _GEN_24[3] & _T_13 & d_response & d_last; // @[src/main/scala/tilelink/Broadcast.scala 142:65]
  assign TLBroadcastTracker_3_io_e_last = _T[3] & auto_in_e_valid; // @[src/main/scala/tilelink/Broadcast.scala 113:34]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 60:30]
      beatsLeft <= 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
    end else if (latch) begin // @[src/main/scala/tilelink/Arbiter.scala 85:23]
      if (winner__1) begin // @[src/main/scala/tilelink/Arbiter.scala 82:69]
        if (beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          beatsLeft <= beats1_decode;
        end else begin
          beatsLeft <= 2'h0;
        end
      end else begin
        beatsLeft <= 2'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_2;
    end
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_T_13) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (d_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          counter <= beats1_decode;
        end else begin
          counter <= 2'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state__1 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state__1 <= winner__1;
    end
    line_508_valid_reg <= _T_13;
    if (d_first) begin // @[src/main/scala/util/package.scala 80:63]
      d_trackerOH_r <= _d_trackerOH_T_8; // @[src/main/scala/util/package.scala 80:63]
    end
    line_509_valid_reg <= d_first;
    line_510_valid_reg <= _T_20;
    line_511_valid_reg <= _T_21;
    line_512_valid_reg <= d_what[1];
    line_513_valid_reg <= _T_20;
    line_514_valid_reg <= _T_30;
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state__0 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state__0 <= winner__0;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 60:30]
      beatsLeft_1 <= 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
    end else if (latch_1) begin // @[src/main/scala/tilelink/Arbiter.scala 85:23]
      beatsLeft_1 <= initBeats_1;
    end else begin
      beatsLeft_1 <= _beatsLeft_T_6;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1_0 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle_1) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1_0 <= winner_1_0;
    end
    line_515_valid_reg <= _clearOH_T;
    line_516_valid_reg <= _T_20;
    line_517_valid_reg <= _T_122;
    line_518_valid_reg <= _T_20;
    line_519_valid_reg <= _T_129;
    line_520_valid_reg <= _T_20;
    line_521_valid_reg <= _T_156;
    line_522_valid_reg <= _T_20;
    line_523_valid_reg <= _T_169;
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1_1 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle_1) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1_1 <= winner_1_1;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1_2 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle_1) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1_2 <= winner_1_2;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1_3 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle_1) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1_3 <= winner_1_3;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1_4 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle_1) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1_4 <= winner_1_4;
    end
    probe_todo <= _GEN_44[0]; // @[src/main/scala/tilelink/Broadcast.scala 215:{31,31}]
    if (_T_196) begin // @[src/main/scala/tilelink/Broadcast.scala 260:38]
      probe_line <= filter_io_response_bits_address[31:5]; // @[src/main/scala/tilelink/Broadcast.scala 262:21]
    end
    if (_T_196) begin // @[src/main/scala/tilelink/Broadcast.scala 260:38]
      if (filter_io_response_bits_needT) begin // @[src/main/scala/tilelink/Broadcast.scala 263:27]
        probe_perms <= 2'h2;
      end else begin
        probe_perms <= 2'h1;
      end
    end
    line_524_valid_reg <= _T_174;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      a_first_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_a_first_T) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (a_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (a_first_beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 2'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    line_525_valid_reg <= _a_first_T;
    line_526_valid_reg <= _T_196;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~auto_out_d_valid | _d_normal_valid_T_1 | auto_out_d_bits_opcode == 3'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Broadcast.scala:125 assert (!out.d.valid || !d_drop || out.d.bits.opcode === TLMessages.AccessAck)\n"
            ); // @[src/main/scala/tilelink/Broadcast.scala 125:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~d_normal_valid | (|_GEN_24 | d_normal_bits_opcode == 3'h6))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Broadcast.scala:137 assert (!d_normal.valid || (d_trackerOH.orR || d_normal.bits.opcode === TLMessages.ReleaseAck))\n"
            ); // @[src/main/scala/tilelink/Broadcast.scala 137:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~winner__0 | ~winner__1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~(releaseack_valid | d_normal_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~((~winner_1_0 | ~winner_1_1) & (~prefixOR_2 | ~winner_1_2) & (~prefixOR_3 | ~winner_1_3) & (~
          prefixOR_4 | ~winner_1_4))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~(putfull_valid | TLBroadcastTracker_io_out_a_valid | TLBroadcastTracker_1_io_out_a_valid |
          TLBroadcastTracker_2_io_out_a_valid | TLBroadcastTracker_3_io_out_a_valid) | _prefixOR_T_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state__1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_508_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  d_trackerOH_r = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  line_509_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_510_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_511_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_512_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_513_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_514_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state__0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  beatsLeft_1 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  state_1_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_515_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_516_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_517_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_518_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_519_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_520_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_521_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_522_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_523_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  state_1_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  state_1_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  state_1_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_1_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  probe_todo = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  probe_line = _RAND_28[26:0];
  _RAND_29 = {1{`RANDOM}};
  probe_perms = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  line_524_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  a_first_counter = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  line_525_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_526_valid_reg = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~auto_out_d_valid | _d_normal_valid_T_1 | auto_out_d_bits_opcode == 3'h0); // @[src/main/scala/tilelink/Broadcast.scala 125:14]
    end
    //
    if (_T_20) begin
      assert(~d_normal_valid | (|_GEN_24 | d_normal_bits_opcode == 3'h6)); // @[src/main/scala/tilelink/Broadcast.scala 137:14]
    end
    //
    if (_T_20) begin
      assert(~winner__0 | ~winner__1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
    end
    //
    if (_T_20) begin
      assert(~(releaseack_valid | d_normal_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
    end
    //
    if (_T_20) begin
      assert((~winner_1_0 | ~winner_1_1) & (~prefixOR_2 | ~winner_1_2) & (~prefixOR_3 | ~winner_1_3) & (~prefixOR_4 | ~
        winner_1_4)); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
    end
    //
    if (_T_20) begin
      assert(~(putfull_valid | TLBroadcastTracker_io_out_a_valid | TLBroadcastTracker_1_io_out_a_valid |
        TLBroadcastTracker_2_io_out_a_valid | TLBroadcastTracker_3_io_out_a_valid) | _prefixOR_T_1); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
    end
  end
endmodule
module TLJbar(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 248:53]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/tilelink/Xbar.scala 163:55]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/tilelink/Xbar.scala 184:55]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 152:69]
endmodule
module BankBinder(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLWidthWidget_6(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLInterconnectCoupler_8(
  input         clock,
  input         reset,
  output        auto_widget_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_widget_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_widget_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_widget_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_widget_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_widget_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_widget_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_widget_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_widget_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_widget_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_widget_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_bus_xing_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_bus_xing_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_bus_xing_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_bus_xing_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_bus_xing_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bus_xing_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_bus_xing_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_bus_xing_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_bus_xing_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bus_xing_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_in_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_in_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_out_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_out_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [3:0] widget_auto_out_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  TLWidthWidget_6 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_auto_out_d_bits_corrupt)
  );
  assign auto_widget_in_a_ready = widget_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_valid = widget_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_size = widget_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_source = widget_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_denied = widget_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_data = widget_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_widget_in_d_bits_corrupt = widget_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bus_xing_out_a_valid = widget_auto_out_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_size = widget_auto_out_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_source = widget_auto_out_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_address = widget_auto_out_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_mask = widget_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_a_bits_data = widget_auto_out_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_bus_xing_out_d_ready = widget_auto_out_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_opcode = auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_size = auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_source = auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_address = auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_mask = auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_a_bits_data = auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_in_d_ready = auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign widget_auto_out_a_ready = auto_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_valid = auto_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_opcode = auto_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_size = auto_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_source = auto_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_denied = auto_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_data = auto_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign widget_auto_out_d_bits_corrupt = auto_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
endmodule
module CoherenceManagerWrapper(
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coherent_jbar_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coherent_jbar_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_coherent_jbar_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_coherent_jbar_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coherent_jbar_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coherent_jbar_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coherent_jbar_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_coherent_jbar_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coherent_jbar_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_coherent_jbar_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coherent_jbar_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_coherent_jbar_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_coherent_jbar_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coherent_jbar_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coherent_jbar_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coherent_jbar_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_coherent_jbar_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coherent_jbar_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_coherent_jbar_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_coherent_jbar_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_coherent_jbar_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_coherent_jbar_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_coherent_jbar_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
  wire  clockGroup_auto_in_member_subsystem_l2_0_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_in_member_subsystem_l2_0_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_clock; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  clockGroup_auto_out_reset; // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
  wire  fixedClockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  fixedClockNode_auto_out_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_1_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_a_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [31:0] broadcast_1_auto_in_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [7:0] broadcast_1_auto_in_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [63:0] broadcast_1_auto_in_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_b_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_b_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_b_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [31:0] broadcast_1_auto_in_b_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_c_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_c_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_c_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_c_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_c_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_c_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [31:0] broadcast_1_auto_in_c_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [63:0] broadcast_1_auto_in_c_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_d_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_in_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_d_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [63:0] broadcast_1_auto_in_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_in_e_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [1:0] broadcast_1_auto_in_e_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_out_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_out_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [3:0] broadcast_1_auto_out_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [31:0] broadcast_1_auto_out_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [7:0] broadcast_1_auto_out_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [63:0] broadcast_1_auto_out_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_out_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [2:0] broadcast_1_auto_out_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [3:0] broadcast_1_auto_out_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire [63:0] broadcast_1_auto_out_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  broadcast_1_auto_out_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
  wire  coherent_jbar_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_a_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_in_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [7:0] coherent_jbar_auto_in_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_in_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_b_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_b_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_b_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_in_b_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_c_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_c_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_c_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_c_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_c_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_c_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_in_c_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_in_c_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_d_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_in_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_d_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_in_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_in_e_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_in_e_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_a_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_out_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [7:0] coherent_jbar_auto_out_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_out_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_b_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_b_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_b_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_out_b_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_c_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_c_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_c_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_c_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_c_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_c_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [31:0] coherent_jbar_auto_out_c_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_out_c_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_d_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [2:0] coherent_jbar_auto_out_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_d_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [63:0] coherent_jbar_auto_out_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  coherent_jbar_auto_out_e_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire [1:0] coherent_jbar_auto_out_e_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
  wire  binder_clock; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_reset; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_a_ready; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_a_valid; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_in_a_bits_size; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [3:0] binder_auto_in_a_bits_source; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [31:0] binder_auto_in_a_bits_address; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [7:0] binder_auto_in_a_bits_mask; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [63:0] binder_auto_in_a_bits_data; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_d_ready; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_d_valid; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_in_d_bits_size; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [3:0] binder_auto_in_d_bits_source; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_d_bits_denied; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [63:0] binder_auto_in_d_bits_data; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_a_ready; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_a_valid; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_out_a_bits_size; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [3:0] binder_auto_out_a_bits_source; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [31:0] binder_auto_out_a_bits_address; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [7:0] binder_auto_out_a_bits_mask; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [63:0] binder_auto_out_a_bits_data; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_d_ready; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_d_valid; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [2:0] binder_auto_out_d_bits_size; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [3:0] binder_auto_out_d_bits_source; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_d_bits_denied; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire [63:0] binder_auto_out_d_bits_data; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  binder_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/BankBinder.scala 68:28]
  wire  coupler_to_bus_named_subsystem_mbus_clock; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_reset; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [31:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [7:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [2:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [3:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire [63:0] coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  wire  coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
  ClockGroupAggregator_5 subsystem_l2_clock_groups ( // @[src/main/scala/tilelink/BusWrapper.scala 39:48]
    .auto_in_member_subsystem_l2_1_clock(subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock),
    .auto_in_member_subsystem_l2_1_reset(subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset),
    .auto_in_member_subsystem_l2_0_clock(subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock),
    .auto_in_member_subsystem_l2_0_reset(subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset),
    .auto_out_1_member_subsystem_mbus_0_clock(subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock),
    .auto_out_1_member_subsystem_mbus_0_reset(subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset),
    .auto_out_0_member_subsystem_l2_0_clock(subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock),
    .auto_out_0_member_subsystem_l2_0_reset(subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset)
  );
  ClockGroup_5 clockGroup ( // @[src/main/scala/tilelink/BusWrapper.scala 40:38]
    .auto_in_member_subsystem_l2_0_clock(clockGroup_auto_in_member_subsystem_l2_0_clock),
    .auto_in_member_subsystem_l2_0_reset(clockGroup_auto_in_member_subsystem_l2_0_reset),
    .auto_out_clock(clockGroup_auto_out_clock),
    .auto_out_reset(clockGroup_auto_out_reset)
  );
  FixedClockBroadcast_5 fixedClockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(fixedClockNode_auto_in_clock),
    .auto_in_reset(fixedClockNode_auto_in_reset),
    .auto_out_clock(fixedClockNode_auto_out_clock),
    .auto_out_reset(fixedClockNode_auto_out_reset)
  );
  BundleBridgeNexus_5 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  TLBroadcast broadcast_1 ( // @[src/main/scala/subsystem/BankedL2Params.scala 82:24]
    .clock(broadcast_1_clock),
    .reset(broadcast_1_reset),
    .auto_in_a_ready(broadcast_1_auto_in_a_ready),
    .auto_in_a_valid(broadcast_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(broadcast_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(broadcast_1_auto_in_a_bits_param),
    .auto_in_a_bits_size(broadcast_1_auto_in_a_bits_size),
    .auto_in_a_bits_source(broadcast_1_auto_in_a_bits_source),
    .auto_in_a_bits_address(broadcast_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(broadcast_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(broadcast_1_auto_in_a_bits_data),
    .auto_in_b_ready(broadcast_1_auto_in_b_ready),
    .auto_in_b_valid(broadcast_1_auto_in_b_valid),
    .auto_in_b_bits_param(broadcast_1_auto_in_b_bits_param),
    .auto_in_b_bits_address(broadcast_1_auto_in_b_bits_address),
    .auto_in_c_ready(broadcast_1_auto_in_c_ready),
    .auto_in_c_valid(broadcast_1_auto_in_c_valid),
    .auto_in_c_bits_opcode(broadcast_1_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(broadcast_1_auto_in_c_bits_param),
    .auto_in_c_bits_size(broadcast_1_auto_in_c_bits_size),
    .auto_in_c_bits_source(broadcast_1_auto_in_c_bits_source),
    .auto_in_c_bits_address(broadcast_1_auto_in_c_bits_address),
    .auto_in_c_bits_data(broadcast_1_auto_in_c_bits_data),
    .auto_in_d_ready(broadcast_1_auto_in_d_ready),
    .auto_in_d_valid(broadcast_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(broadcast_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(broadcast_1_auto_in_d_bits_param),
    .auto_in_d_bits_size(broadcast_1_auto_in_d_bits_size),
    .auto_in_d_bits_source(broadcast_1_auto_in_d_bits_source),
    .auto_in_d_bits_sink(broadcast_1_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(broadcast_1_auto_in_d_bits_denied),
    .auto_in_d_bits_data(broadcast_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(broadcast_1_auto_in_d_bits_corrupt),
    .auto_in_e_valid(broadcast_1_auto_in_e_valid),
    .auto_in_e_bits_sink(broadcast_1_auto_in_e_bits_sink),
    .auto_out_a_ready(broadcast_1_auto_out_a_ready),
    .auto_out_a_valid(broadcast_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(broadcast_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(broadcast_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(broadcast_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(broadcast_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(broadcast_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(broadcast_1_auto_out_a_bits_data),
    .auto_out_d_ready(broadcast_1_auto_out_d_ready),
    .auto_out_d_valid(broadcast_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(broadcast_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(broadcast_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(broadcast_1_auto_out_d_bits_source),
    .auto_out_d_bits_denied(broadcast_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(broadcast_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(broadcast_1_auto_out_d_bits_corrupt)
  );
  TLJbar coherent_jbar ( // @[src/main/scala/subsystem/BankedL2Params.scala 59:41]
    .clock(coherent_jbar_clock),
    .reset(coherent_jbar_reset),
    .auto_in_a_ready(coherent_jbar_auto_in_a_ready),
    .auto_in_a_valid(coherent_jbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(coherent_jbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(coherent_jbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(coherent_jbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(coherent_jbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(coherent_jbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(coherent_jbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(coherent_jbar_auto_in_a_bits_data),
    .auto_in_b_ready(coherent_jbar_auto_in_b_ready),
    .auto_in_b_valid(coherent_jbar_auto_in_b_valid),
    .auto_in_b_bits_param(coherent_jbar_auto_in_b_bits_param),
    .auto_in_b_bits_address(coherent_jbar_auto_in_b_bits_address),
    .auto_in_c_ready(coherent_jbar_auto_in_c_ready),
    .auto_in_c_valid(coherent_jbar_auto_in_c_valid),
    .auto_in_c_bits_opcode(coherent_jbar_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(coherent_jbar_auto_in_c_bits_param),
    .auto_in_c_bits_size(coherent_jbar_auto_in_c_bits_size),
    .auto_in_c_bits_source(coherent_jbar_auto_in_c_bits_source),
    .auto_in_c_bits_address(coherent_jbar_auto_in_c_bits_address),
    .auto_in_c_bits_data(coherent_jbar_auto_in_c_bits_data),
    .auto_in_d_ready(coherent_jbar_auto_in_d_ready),
    .auto_in_d_valid(coherent_jbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(coherent_jbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(coherent_jbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(coherent_jbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(coherent_jbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(coherent_jbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(coherent_jbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(coherent_jbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(coherent_jbar_auto_in_d_bits_corrupt),
    .auto_in_e_valid(coherent_jbar_auto_in_e_valid),
    .auto_in_e_bits_sink(coherent_jbar_auto_in_e_bits_sink),
    .auto_out_a_ready(coherent_jbar_auto_out_a_ready),
    .auto_out_a_valid(coherent_jbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(coherent_jbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(coherent_jbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(coherent_jbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(coherent_jbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(coherent_jbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(coherent_jbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(coherent_jbar_auto_out_a_bits_data),
    .auto_out_b_ready(coherent_jbar_auto_out_b_ready),
    .auto_out_b_valid(coherent_jbar_auto_out_b_valid),
    .auto_out_b_bits_param(coherent_jbar_auto_out_b_bits_param),
    .auto_out_b_bits_address(coherent_jbar_auto_out_b_bits_address),
    .auto_out_c_ready(coherent_jbar_auto_out_c_ready),
    .auto_out_c_valid(coherent_jbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(coherent_jbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(coherent_jbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(coherent_jbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(coherent_jbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(coherent_jbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(coherent_jbar_auto_out_c_bits_data),
    .auto_out_d_ready(coherent_jbar_auto_out_d_ready),
    .auto_out_d_valid(coherent_jbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(coherent_jbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(coherent_jbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(coherent_jbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(coherent_jbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(coherent_jbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(coherent_jbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(coherent_jbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(coherent_jbar_auto_out_d_bits_corrupt),
    .auto_out_e_valid(coherent_jbar_auto_out_e_valid),
    .auto_out_e_bits_sink(coherent_jbar_auto_out_e_bits_sink)
  );
  BankBinder binder ( // @[src/main/scala/tilelink/BankBinder.scala 68:28]
    .clock(binder_clock),
    .reset(binder_reset),
    .auto_in_a_ready(binder_auto_in_a_ready),
    .auto_in_a_valid(binder_auto_in_a_valid),
    .auto_in_a_bits_opcode(binder_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(binder_auto_in_a_bits_size),
    .auto_in_a_bits_source(binder_auto_in_a_bits_source),
    .auto_in_a_bits_address(binder_auto_in_a_bits_address),
    .auto_in_a_bits_mask(binder_auto_in_a_bits_mask),
    .auto_in_a_bits_data(binder_auto_in_a_bits_data),
    .auto_in_d_ready(binder_auto_in_d_ready),
    .auto_in_d_valid(binder_auto_in_d_valid),
    .auto_in_d_bits_opcode(binder_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(binder_auto_in_d_bits_size),
    .auto_in_d_bits_source(binder_auto_in_d_bits_source),
    .auto_in_d_bits_denied(binder_auto_in_d_bits_denied),
    .auto_in_d_bits_data(binder_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(binder_auto_in_d_bits_corrupt),
    .auto_out_a_ready(binder_auto_out_a_ready),
    .auto_out_a_valid(binder_auto_out_a_valid),
    .auto_out_a_bits_opcode(binder_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(binder_auto_out_a_bits_size),
    .auto_out_a_bits_source(binder_auto_out_a_bits_source),
    .auto_out_a_bits_address(binder_auto_out_a_bits_address),
    .auto_out_a_bits_mask(binder_auto_out_a_bits_mask),
    .auto_out_a_bits_data(binder_auto_out_a_bits_data),
    .auto_out_d_ready(binder_auto_out_d_ready),
    .auto_out_d_valid(binder_auto_out_d_valid),
    .auto_out_d_bits_opcode(binder_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(binder_auto_out_d_bits_size),
    .auto_out_d_bits_source(binder_auto_out_d_bits_source),
    .auto_out_d_bits_denied(binder_auto_out_d_bits_denied),
    .auto_out_d_bits_data(binder_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(binder_auto_out_d_bits_corrupt)
  );
  TLInterconnectCoupler_8 coupler_to_bus_named_subsystem_mbus ( // @[src/main/scala/diplomacy/LazyModule.scala 493:27]
    .clock(coupler_to_bus_named_subsystem_mbus_clock),
    .reset(coupler_to_bus_named_subsystem_mbus_reset),
    .auto_widget_in_a_ready(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready),
    .auto_widget_in_a_valid(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid),
    .auto_widget_in_a_bits_opcode(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode),
    .auto_widget_in_a_bits_size(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size),
    .auto_widget_in_a_bits_source(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source),
    .auto_widget_in_a_bits_address(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address),
    .auto_widget_in_a_bits_mask(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask),
    .auto_widget_in_a_bits_data(coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data),
    .auto_widget_in_d_ready(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready),
    .auto_widget_in_d_valid(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid),
    .auto_widget_in_d_bits_opcode(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode),
    .auto_widget_in_d_bits_size(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size),
    .auto_widget_in_d_bits_source(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source),
    .auto_widget_in_d_bits_denied(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied),
    .auto_widget_in_d_bits_data(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data),
    .auto_widget_in_d_bits_corrupt(coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt),
    .auto_bus_xing_out_a_ready(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready),
    .auto_bus_xing_out_a_valid(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid),
    .auto_bus_xing_out_a_bits_opcode(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode),
    .auto_bus_xing_out_a_bits_size(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size),
    .auto_bus_xing_out_a_bits_source(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source),
    .auto_bus_xing_out_a_bits_address(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address),
    .auto_bus_xing_out_a_bits_mask(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask),
    .auto_bus_xing_out_a_bits_data(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data),
    .auto_bus_xing_out_d_ready(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready),
    .auto_bus_xing_out_d_valid(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid),
    .auto_bus_xing_out_d_bits_opcode(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode),
    .auto_bus_xing_out_d_bits_size(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size),
    .auto_bus_xing_out_d_bits_source(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source),
    .auto_bus_xing_out_d_bits_denied(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied),
    .auto_bus_xing_out_d_bits_data(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data),
    .auto_bus_xing_out_d_bits_corrupt(coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt)
  );
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready =
    coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_coherent_jbar_in_a_ready = coherent_jbar_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_b_valid = coherent_jbar_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_b_bits_param = coherent_jbar_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_b_bits_address = coherent_jbar_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_c_ready = coherent_jbar_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_valid = coherent_jbar_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_opcode = coherent_jbar_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_param = coherent_jbar_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_size = coherent_jbar_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_source = coherent_jbar_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_sink = coherent_jbar_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_denied = coherent_jbar_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_data = coherent_jbar_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_coherent_jbar_in_d_bits_corrupt = coherent_jbar_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock =
    subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset =
    subsystem_l2_clock_groups_auto_out_1_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_clock =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_1_reset =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_clock =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign subsystem_l2_clock_groups_auto_in_member_subsystem_l2_0_reset =
    auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockGroup_auto_in_member_subsystem_l2_0_clock =
    subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign clockGroup_auto_in_member_subsystem_l2_0_reset =
    subsystem_l2_clock_groups_auto_out_0_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_clock = clockGroup_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign fixedClockNode_auto_in_reset = clockGroup_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_valid = coherent_jbar_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_opcode = coherent_jbar_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_param = coherent_jbar_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_size = coherent_jbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_source = coherent_jbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_address = coherent_jbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_mask = coherent_jbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_a_bits_data = coherent_jbar_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_b_ready = coherent_jbar_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_valid = coherent_jbar_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_opcode = coherent_jbar_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_param = coherent_jbar_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_size = coherent_jbar_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_source = coherent_jbar_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_address = coherent_jbar_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_c_bits_data = coherent_jbar_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_d_ready = coherent_jbar_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_e_valid = coherent_jbar_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_in_e_bits_sink = coherent_jbar_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign broadcast_1_auto_out_a_ready = binder_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_valid = binder_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_opcode = binder_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_size = binder_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_source = binder_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_denied = binder_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_data = binder_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign broadcast_1_auto_out_d_bits_corrupt = binder_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coherent_jbar_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_in_a_valid = auto_coherent_jbar_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_opcode = auto_coherent_jbar_in_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_param = auto_coherent_jbar_in_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_size = auto_coherent_jbar_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_source = auto_coherent_jbar_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_address = auto_coherent_jbar_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_mask = auto_coherent_jbar_in_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_a_bits_data = auto_coherent_jbar_in_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_b_ready = auto_coherent_jbar_in_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_valid = auto_coherent_jbar_in_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_opcode = auto_coherent_jbar_in_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_param = auto_coherent_jbar_in_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_size = auto_coherent_jbar_in_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_source = auto_coherent_jbar_in_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_address = auto_coherent_jbar_in_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_c_bits_data = auto_coherent_jbar_in_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_d_ready = auto_coherent_jbar_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_e_valid = auto_coherent_jbar_in_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_in_e_bits_sink = auto_coherent_jbar_in_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign coherent_jbar_auto_out_a_ready = broadcast_1_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_b_valid = broadcast_1_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_b_bits_param = broadcast_1_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_b_bits_address = broadcast_1_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_c_ready = broadcast_1_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_valid = broadcast_1_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_opcode = broadcast_1_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_param = broadcast_1_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_size = broadcast_1_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_source = broadcast_1_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_sink = broadcast_1_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_denied = broadcast_1_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_data = broadcast_1_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coherent_jbar_auto_out_d_bits_corrupt = broadcast_1_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign binder_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign binder_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign binder_auto_in_a_valid = broadcast_1_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_opcode = broadcast_1_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_size = broadcast_1_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_source = broadcast_1_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_address = broadcast_1_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_mask = broadcast_1_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_a_bits_data = broadcast_1_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_in_d_ready = broadcast_1_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_a_ready = coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_valid = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_opcode = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_size = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_source = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_denied = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_data = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign binder_auto_out_d_bits_corrupt = coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_clock = fixedClockNode_auto_out_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_mbus_reset = fixedClockNode_auto_out_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_valid = binder_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_opcode = binder_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_size = binder_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_source = binder_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_address = binder_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_mask = binder_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_a_bits_data = binder_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_widget_in_d_ready = binder_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_a_ready =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_valid =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_opcode =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_size =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_source =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_denied =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_data =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign coupler_to_bus_named_subsystem_mbus_auto_bus_xing_out_d_bits_corrupt =
    auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
endmodule
module TLXbar_8(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_1_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_1_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_1_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_1_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_1_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_1_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_1_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_0_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_0_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_0_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_0_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_0_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_0_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_0_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_0_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_0_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_0_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_0_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_0_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_0_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_0_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_0_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_0_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_0_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  requestBOI_0_0 = ~auto_out_b_bits_source[1]; // @[src/main/scala/diplomacy/Parameters.scala 54:32]
  wire  requestDOI_0_0 = ~auto_out_d_bits_source[1]; // @[src/main/scala/diplomacy/Parameters.scala 54:32]
  wire  requestDOI_0_1 = auto_out_d_bits_source == 2'h2; // @[src/main/scala/diplomacy/Parameters.scala 46:9]
  wire [11:0] _beatsAI_decode_T_1 = 12'h1f << auto_in_0_a_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beatsAI_decode_T_3 = ~_beatsAI_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beatsAI_decode = _beatsAI_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  beatsAI_opdata = ~auto_in_0_a_bits_opcode[2]; // @[src/main/scala/tilelink/Edges.scala 92:28]
  reg [1:0] beatsLeft; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
  wire  idle = beatsLeft == 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 61:28]
  wire  latch = idle & auto_out_a_ready; // @[src/main/scala/tilelink/Arbiter.scala 62:24]
  wire [1:0] readys_valid = {auto_in_1_a_valid,auto_in_0_a_valid}; // @[src/main/scala/tilelink/Arbiter.scala 68:51]
  wire  _readys_T_3 = ~reset; // @[src/main/scala/tilelink/Arbiter.scala 22:12]
  wire  line_527_clock;
  wire  line_527_reset;
  wire  line_527_valid;
  reg  line_527_valid_reg;
  reg [1:0] readys_mask; // @[src/main/scala/tilelink/Arbiter.scala 23:23]
  wire [1:0] _readys_filter_T = ~readys_mask; // @[src/main/scala/tilelink/Arbiter.scala 24:30]
  wire [1:0] _readys_filter_T_1 = readys_valid & _readys_filter_T; // @[src/main/scala/tilelink/Arbiter.scala 24:28]
  wire [3:0] readys_filter = {_readys_filter_T_1,auto_in_1_a_valid,auto_in_0_a_valid}; // @[src/main/scala/tilelink/Arbiter.scala 24:21]
  wire [3:0] _GEN_8 = {{1'd0}, readys_filter[3:1]}; // @[src/main/scala/util/package.scala 254:43]
  wire [3:0] _readys_unready_T_1 = readys_filter | _GEN_8; // @[src/main/scala/util/package.scala 254:43]
  wire [3:0] _readys_unready_T_4 = {readys_mask, 2'h0}; // @[src/main/scala/tilelink/Arbiter.scala 25:66]
  wire [3:0] _GEN_9 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[src/main/scala/tilelink/Arbiter.scala 25:58]
  wire [3:0] readys_unready = _GEN_9 | _readys_unready_T_4; // @[src/main/scala/tilelink/Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[src/main/scala/tilelink/Arbiter.scala 26:39]
  wire [1:0] readys_readys = ~_readys_readys_T_2; // @[src/main/scala/tilelink/Arbiter.scala 26:18]
  wire  _readys_T_6 = latch & |readys_valid; // @[src/main/scala/tilelink/Arbiter.scala 27:18]
  wire  line_528_clock;
  wire  line_528_reset;
  wire  line_528_valid;
  reg  line_528_valid_reg;
  wire [1:0] _readys_mask_T = readys_readys & readys_valid; // @[src/main/scala/tilelink/Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[src/main/scala/util/package.scala 245:48]
  wire [1:0] _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[src/main/scala/util/package.scala 245:43]
  wire  readys_0 = readys_readys[0]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  readys_1 = readys_readys[1]; // @[src/main/scala/tilelink/Arbiter.scala 68:76]
  wire  winner_0 = readys_0 & auto_in_0_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  winner_1 = readys_1 & auto_in_1_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 71:69]
  wire  _prefixOR_T = winner_0 | winner_1; // @[src/main/scala/tilelink/Arbiter.scala 76:48]
  wire  line_529_clock;
  wire  line_529_reset;
  wire  line_529_valid;
  reg  line_529_valid_reg;
  wire  _T_9 = ~(~winner_0 | ~winner_1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
  wire  line_530_clock;
  wire  line_530_reset;
  wire  line_530_valid;
  reg  line_530_valid_reg;
  wire  _T_10 = auto_in_0_a_valid | auto_in_1_a_valid; // @[src/main/scala/tilelink/Arbiter.scala 79:31]
  wire  line_531_clock;
  wire  line_531_reset;
  wire  line_531_valid;
  reg  line_531_valid_reg;
  wire  _T_16 = ~(~(auto_in_0_a_valid | auto_in_1_a_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
  wire  line_532_clock;
  wire  line_532_reset;
  wire  line_532_valid;
  reg  line_532_valid_reg;
  reg  state_0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  reg  state_1; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
  wire  _out_0_a_valid_T_3 = state_0 & auto_in_0_a_valid | state_1 & auto_in_1_a_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  out_0_a_valid = idle ? _T_10 : _out_0_a_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  wire  _beatsLeft_T = auto_out_a_ready & out_0_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_10 = {{1'd0}, _beatsLeft_T}; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire [1:0] _beatsLeft_T_2 = beatsLeft - _GEN_10; // @[src/main/scala/tilelink/Arbiter.scala 85:52]
  wire  muxState_0 = idle ? winner_0 : state_0; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  muxState_1 = idle ? winner_1 : state_1; // @[src/main/scala/tilelink/Arbiter.scala 89:25]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[src/main/scala/tilelink/Arbiter.scala 92:24]
  wire [7:0] _out_0_a_bits_T_6 = muxState_0 ? auto_in_0_a_bits_mask : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _out_0_a_bits_T_7 = muxState_1 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _out_0_a_bits_T_9 = muxState_0 ? auto_in_0_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _out_0_a_bits_T_10 = muxState_1 ? auto_in_1_a_bits_address : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] in_0_a_bits_source = {{1'd0}, auto_in_0_a_bits_source}; // @[src/main/scala/tilelink/Xbar.scala 155:18 163:29]
  wire [1:0] _out_0_a_bits_T_12 = muxState_0 ? in_0_a_bits_source : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _out_0_a_bits_T_13 = muxState_1 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _out_0_a_bits_T_15 = muxState_0 ? auto_in_0_a_bits_size : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _out_0_a_bits_T_16 = muxState_1 ? 3'h5 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _out_0_a_bits_T_21 = muxState_0 ? auto_in_0_a_bits_opcode : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [2:0] _out_0_a_bits_T_22 = muxState_1 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  GEN_w1_line #(.COVER_INDEX(527)) line_527 (
    .clock(line_527_clock),
    .reset(line_527_reset),
    .valid(line_527_valid)
  );
  GEN_w1_line #(.COVER_INDEX(528)) line_528 (
    .clock(line_528_clock),
    .reset(line_528_reset),
    .valid(line_528_valid)
  );
  GEN_w1_line #(.COVER_INDEX(529)) line_529 (
    .clock(line_529_clock),
    .reset(line_529_reset),
    .valid(line_529_valid)
  );
  GEN_w1_line #(.COVER_INDEX(530)) line_530 (
    .clock(line_530_clock),
    .reset(line_530_reset),
    .valid(line_530_valid)
  );
  GEN_w1_line #(.COVER_INDEX(531)) line_531 (
    .clock(line_531_clock),
    .reset(line_531_reset),
    .valid(line_531_valid)
  );
  GEN_w1_line #(.COVER_INDEX(532)) line_532 (
    .clock(line_532_clock),
    .reset(line_532_reset),
    .valid(line_532_valid)
  );
  assign line_527_clock = clock;
  assign line_527_reset = reset;
  assign line_527_valid = _readys_T_3 ^ line_527_valid_reg;
  assign line_528_clock = clock;
  assign line_528_reset = reset;
  assign line_528_valid = _readys_T_6 ^ line_528_valid_reg;
  assign line_529_clock = clock;
  assign line_529_reset = reset;
  assign line_529_valid = _readys_T_3 ^ line_529_valid_reg;
  assign line_530_clock = clock;
  assign line_530_reset = reset;
  assign line_530_valid = _T_9 ^ line_530_valid_reg;
  assign line_531_clock = clock;
  assign line_531_reset = reset;
  assign line_531_valid = _readys_T_3 ^ line_531_valid_reg;
  assign line_532_clock = clock;
  assign line_532_reset = reset;
  assign line_532_valid = _T_16 ^ line_532_valid_reg;
  assign auto_in_1_a_ready = auto_out_a_ready & allowed_1; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_a_ready = auto_out_a_ready & allowed_0; // @[src/main/scala/tilelink/Arbiter.scala 94:31]
  assign auto_in_0_b_valid = auto_out_b_valid & requestBOI_0_0; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_0_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_b_bits_size = auto_out_b_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_b_bits_source = auto_out_b_bits_source[0]; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_0_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  assign auto_in_0_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 248:53]
  assign auto_in_0_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_0_e_ready = auto_out_e_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = idle ? _T_10 : _out_0_a_valid_T_3; // @[src/main/scala/tilelink/Arbiter.scala 96:24]
  assign auto_out_a_bits_opcode = _out_0_a_bits_T_21 | _out_0_a_bits_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_param = muxState_0 ? auto_in_0_a_bits_param : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_size = _out_0_a_bits_T_15 | _out_0_a_bits_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_source = _out_0_a_bits_T_12 | _out_0_a_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_address = _out_0_a_bits_T_9 | _out_0_a_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_mask = _out_0_a_bits_T_6 | _out_0_a_bits_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_a_bits_data = muxState_0 ? auto_in_0_a_bits_data : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_b_ready = requestBOI_0_0 & auto_in_0_b_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_c_valid = auto_in_0_c_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_c_bits_opcode = auto_in_0_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_0_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_0_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = {{1'd0}, auto_in_0_c_bits_source}; // @[src/main/scala/tilelink/Xbar.scala 155:18 184:29]
  assign auto_out_c_bits_address = auto_in_0_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_0_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = requestDOI_0_0 & auto_in_0_d_ready | requestDOI_0_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign auto_out_e_valid = auto_in_0_e_valid; // @[src/main/scala/tilelink/Xbar.scala 352:40]
  assign auto_out_e_bits_sink = auto_in_0_e_bits_sink; // @[src/main/scala/tilelink/Xbar.scala 152:69]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 60:30]
      beatsLeft <= 2'h0; // @[src/main/scala/tilelink/Arbiter.scala 60:30]
    end else if (latch) begin // @[src/main/scala/tilelink/Arbiter.scala 85:23]
      if (winner_0) begin // @[src/main/scala/tilelink/Arbiter.scala 82:69]
        if (beatsAI_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          beatsLeft <= beatsAI_decode;
        end else begin
          beatsLeft <= 2'h0;
        end
      end else begin
        beatsLeft <= 2'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_2;
    end
    line_527_valid_reg <= _readys_T_3;
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 23:23]
      readys_mask <= 2'h3; // @[src/main/scala/tilelink/Arbiter.scala 23:23]
    end else if (latch & |readys_valid) begin // @[src/main/scala/tilelink/Arbiter.scala 27:32]
      readys_mask <= _readys_mask_T_3; // @[src/main/scala/tilelink/Arbiter.scala 28:12]
    end
    line_528_valid_reg <= _readys_T_6;
    line_529_valid_reg <= _readys_T_3;
    line_530_valid_reg <= _T_9;
    line_531_valid_reg <= _readys_T_3;
    line_532_valid_reg <= _T_16;
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_0 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_0 <= winner_0;
    end
    if (reset) begin // @[src/main/scala/tilelink/Arbiter.scala 88:26]
      state_1 <= 1'h0; // @[src/main/scala/tilelink/Arbiter.scala 88:26]
    end else if (idle) begin // @[src/main/scala/tilelink/Arbiter.scala 89:25]
      state_1 <= winner_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~winner_0 | ~winner_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_readys_T_3 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n"); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  line_527_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  readys_mask = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  line_528_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_529_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_530_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_531_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_532_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/tilelink/Arbiter.scala 22:12]
    end
    //
    if (_readys_T_3) begin
      assert(~winner_0 | ~winner_1); // @[src/main/scala/tilelink/Arbiter.scala 77:13]
    end
    //
    if (_readys_T_3) begin
      assert(~(auto_in_0_a_valid | auto_in_1_a_valid) | _prefixOR_T); // @[src/main/scala/tilelink/Arbiter.scala 79:14]
    end
  end
endmodule
module TLXbar_9(
  input   clock,
  input   reset
);
endmodule
module IntXbar_1(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_6(
  input   clock,
  input   reset,
  input   auto_in, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out = auto_in; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module BundleBridgeNexus_7(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_8(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_9(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_10(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_11(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_12(
  input   clock,
  input   reset
);
endmodule
module TLWidthWidget_7(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_size = auto_out_b_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_source = auto_out_b_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_e_ready = auto_out_e_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module OptimizationBarrier(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
endmodule
module PMPChecker(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_1(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ppp, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pal, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_paa, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_eff, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ppp, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pal, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_paa, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_eff, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sw = io_x_sw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sr = io_x_sr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pw = io_x_pw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pr = io_x_pr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ppp = io_x_ppp; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pal = io_x_pal; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_paa = io_x_paa; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_eff = io_x_eff; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_2(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ppp, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pal, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_paa, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_eff, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ppp, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pal, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_paa, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_eff, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sw = io_x_sw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sr = io_x_sr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pw = io_x_pw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pr = io_x_pr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ppp = io_x_ppp; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pal = io_x_pal; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_paa = io_x_paa; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_eff = io_x_eff; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_3(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ppp, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pal, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_paa, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_eff, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ppp, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pal, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_paa, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_eff, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sw = io_x_sw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sr = io_x_sr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pw = io_x_pw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pr = io_x_pr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ppp = io_x_ppp; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pal = io_x_pal; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_paa = io_x_paa; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_eff = io_x_eff; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_4(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pr, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ppp, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pal, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_paa, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_eff, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pr, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ppp, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pal, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_paa, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_eff, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sw = io_x_sw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sr = io_x_sr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pw = io_x_pw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pr = io_x_pr; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ppp = io_x_ppp; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pal = io_x_pal; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_paa = io_x_paa; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_eff = io_x_eff; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_5(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sr, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sr // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sw = io_x_sw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sr = io_x_sr; // @[src/main/scala/util/package.scala 264:12]
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_req_ready, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_req_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [39:0] io_req_bits_vaddr, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_req_bits_passthrough, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [1:0]  io_req_bits_size, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [4:0]  io_req_bits_cmd, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [1:0]  io_req_bits_prv, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_miss, // @[src/main/scala/rocket/TLB.scala 309:14]
  output [31:0] io_resp_paddr, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_pf_ld, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_pf_st, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_ae_ld, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_ae_st, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_ma_ld, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_ma_st, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_cacheable, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_bits_rs1, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_bits_rs2, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [38:0] io_sfence_bits_addr, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_req_ready, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_bits_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  output [26:0] io_ptw_req_bits_bits_addr, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_bits_bits_need_gpa, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_ae_ptw, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_ae_final, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pf, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [43:0] io_ptw_resp_bits_pte_ppn, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_d, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_a, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_g, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_u, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_x, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_w, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_r, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_v, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [1:0]  io_ptw_resp_bits_level, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_homogeneous, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [3:0]  io_ptw_ptbr_mode, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_status_mxr, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_status_sum // @[src/main/scala/rocket/TLB.scala 309:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
`endif // RANDOMIZE_REG_INIT
  wire  mpu_ppn_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  mpu_ppn_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] mpu_ppn_barrier_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] mpu_ppn_barrier_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  pmp_clock; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  pmp_reset; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  entries_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_1_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_1_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_2_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_2_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_3_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_3_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_sr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_pw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_pr; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_ppp; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_pal; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_paa; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_eff; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_4_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_sr; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_4_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_sw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_sr; // @[src/main/scala/util/package.scala 259:25]
  wire [26:0] vpn = io_req_bits_vaddr[38:12]; // @[src/main/scala/rocket/TLB.scala 324:30]
  reg [26:0] sectored_entries_0_0_tag_vpn; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [26:0] sectored_entries_0_1_tag_vpn; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [1:0] superpage_entries_0_level; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [26:0] superpage_entries_0_tag_vpn; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [41:0] superpage_entries_0_data_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg  superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [1:0] superpage_entries_1_level; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [26:0] superpage_entries_1_tag_vpn; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [41:0] superpage_entries_1_data_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg  superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [1:0] special_entry_level; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [26:0] special_entry_tag_vpn; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [41:0] special_entry_data_0; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg  special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [1:0] state; // @[src/main/scala/rocket/TLB.scala 341:22]
  reg [26:0] r_refill_tag; // @[src/main/scala/rocket/TLB.scala 343:25]
  reg  r_superpage_repl_addr; // @[src/main/scala/rocket/TLB.scala 344:34]
  reg  r_sectored_repl_addr; // @[src/main/scala/rocket/TLB.scala 345:33]
  reg  r_sectored_hit_valid; // @[src/main/scala/rocket/TLB.scala 346:27]
  reg  r_sectored_hit_bits; // @[src/main/scala/rocket/TLB.scala 346:27]
  reg  r_need_gpa; // @[src/main/scala/rocket/TLB.scala 350:23]
  wire  priv_s = io_req_bits_prv[0]; // @[src/main/scala/rocket/TLB.scala 359:20]
  wire  priv_uses_vm = io_req_bits_prv <= 2'h1; // @[src/main/scala/rocket/TLB.scala 361:27]
  wire  stage1_en = io_ptw_ptbr_mode[3]; // @[src/main/scala/rocket/TLB.scala 363:41]
  wire  vm_enabled = stage1_en & priv_uses_vm & ~io_req_bits_passthrough; // @[src/main/scala/rocket/TLB.scala 388:61]
  wire [19:0] refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[src/main/scala/rocket/TLB.scala 395:44]
  wire  _invalidate_refill_T = state == 2'h1; // @[src/main/scala/util/package.scala 16:47]
  wire  _invalidate_refill_T_1 = state == 2'h3; // @[src/main/scala/util/package.scala 16:47]
  wire  _invalidate_refill_T_2 = _invalidate_refill_T | _invalidate_refill_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  invalidate_refill = _invalidate_refill_T_2 | io_sfence_valid; // @[src/main/scala/rocket/TLB.scala 399:88]
  wire [1:0] mpu_ppn_res = mpu_ppn_barrier_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire  mpu_ppn_ignore = special_entry_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 187:28]
  wire [26:0] _mpu_ppn_T_24 = mpu_ppn_ignore ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_488 = {{7'd0}, mpu_ppn_barrier_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _mpu_ppn_T_25 = _mpu_ppn_T_24 | _GEN_488; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire  mpu_ppn_ignore_1 = special_entry_level < 2'h2; // @[src/main/scala/rocket/TLB.scala 187:28]
  wire [26:0] _mpu_ppn_T_28 = mpu_ppn_ignore_1 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _mpu_ppn_T_29 = _mpu_ppn_T_28 | _GEN_488; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _mpu_ppn_T_31 = {mpu_ppn_res,_mpu_ppn_T_25[17:9],_mpu_ppn_T_29[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [27:0] _mpu_ppn_T_33 = vm_enabled ? {{8'd0}, _mpu_ppn_T_31} : io_req_bits_vaddr[39:12]; // @[src/main/scala/rocket/TLB.scala 402:20]
  wire [27:0] mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _mpu_ppn_T_33; // @[src/main/scala/rocket/TLB.scala 401:20]
  wire [39:0] mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[src/main/scala/rocket/TLB.scala 403:25]
  wire [39:0] _legal_address_T = mpu_physaddr ^ 40'h10000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [40:0] _legal_address_T_1 = {1'b0,$signed(_legal_address_T)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [40:0] _legal_address_T_3 = $signed(_legal_address_T_1) & -41'sh10000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _legal_address_T_4 = $signed(_legal_address_T_3) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire [39:0] _legal_address_T_5 = mpu_physaddr ^ 40'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [40:0] _legal_address_T_6 = {1'b0,$signed(_legal_address_T_5)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [40:0] _legal_address_T_8 = $signed(_legal_address_T_6) & -41'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _legal_address_T_9 = $signed(_legal_address_T_8) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire  legal_address = _legal_address_T_4 | _legal_address_T_9; // @[src/main/scala/rocket/TLB.scala 412:67]
  wire [40:0] _cacheable_T_8 = $signed(_legal_address_T_6) & 41'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _cacheable_T_9 = $signed(_cacheable_T_8) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire  cacheable = legal_address & _cacheable_T_9; // @[src/main/scala/rocket/TLB.scala 415:19]
  wire  _sector_hits_T_2 = sectored_entries_0_0_valid_0 | sectored_entries_0_0_valid_1 | sectored_entries_0_0_valid_2 |
    sectored_entries_0_0_valid_3; // @[src/main/scala/util/package.scala 73:59]
  wire [26:0] _sector_hits_T_3 = sectored_entries_0_0_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 164:61]
  wire  _sector_hits_T_5 = _sector_hits_T_3[26:2] == 25'h0; // @[src/main/scala/rocket/TLB.scala 164:86]
  wire  sector_hits_0 = _sector_hits_T_2 & _sector_hits_T_5; // @[src/main/scala/rocket/TLB.scala 162:55]
  wire  _sector_hits_T_10 = sectored_entries_0_1_valid_0 | sectored_entries_0_1_valid_1 | sectored_entries_0_1_valid_2
     | sectored_entries_0_1_valid_3; // @[src/main/scala/util/package.scala 73:59]
  wire [26:0] _sector_hits_T_11 = sectored_entries_0_1_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 164:61]
  wire  _sector_hits_T_13 = _sector_hits_T_11[26:2] == 25'h0; // @[src/main/scala/rocket/TLB.scala 164:86]
  wire  sector_hits_1 = _sector_hits_T_10 & _sector_hits_T_13; // @[src/main/scala/rocket/TLB.scala 162:55]
  wire [26:0] _superpage_hits_T = superpage_entries_0_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  superpage_hits_ignore_1 = superpage_entries_0_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 172:28]
  wire  superpage_hits_0 = superpage_entries_0_valid_0 & _superpage_hits_T[26:18] == 9'h0 & (superpage_hits_ignore_1 |
    _superpage_hits_T[17:9] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire [26:0] _superpage_hits_T_14 = superpage_entries_1_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  superpage_hits_ignore_4 = superpage_entries_1_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 172:28]
  wire  superpage_hits_1 = superpage_entries_1_valid_0 & _superpage_hits_T_14[26:18] == 9'h0 & (superpage_hits_ignore_4
     | _superpage_hits_T_14[17:9] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire [1:0] hitsVec_idx = vpn[1:0]; // @[src/main/scala/util/package.scala 155:13]
  wire  _GEN_0 = 2'h0 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_533_clock;
  wire  line_533_reset;
  wire  line_533_valid;
  reg  line_533_valid_reg;
  wire  _GEN_1 = 2'h1 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_534_clock;
  wire  line_534_reset;
  wire  line_534_valid;
  reg  line_534_valid_reg;
  wire  _GEN_146 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_valid_1 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _GEN_2 = 2'h2 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_535_clock;
  wire  line_535_reset;
  wire  line_535_valid;
  reg  line_535_valid_reg;
  wire  _GEN_147 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_valid_2 : _GEN_146; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _GEN_3 = 2'h3 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_536_clock;
  wire  line_536_reset;
  wire  line_536_valid;
  reg  line_536_valid_reg;
  wire  _GEN_148 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_valid_3 : _GEN_147; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _hitsVec_T_5 = _GEN_148 & _sector_hits_T_5; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  hitsVec_0 = vm_enabled & _hitsVec_T_5; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  line_537_clock;
  wire  line_537_reset;
  wire  line_537_valid;
  reg  line_537_valid_reg;
  wire  line_538_clock;
  wire  line_538_reset;
  wire  line_538_valid;
  reg  line_538_valid_reg;
  wire  _GEN_150 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_valid_1 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  line_539_clock;
  wire  line_539_reset;
  wire  line_539_valid;
  reg  line_539_valid_reg;
  wire  _GEN_151 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_valid_2 : _GEN_150; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  line_540_clock;
  wire  line_540_reset;
  wire  line_540_valid;
  reg  line_540_valid_reg;
  wire  _GEN_152 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_valid_3 : _GEN_151; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _hitsVec_T_11 = _GEN_152 & _sector_hits_T_13; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  hitsVec_1 = vm_enabled & _hitsVec_T_11; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  hitsVec_2 = vm_enabled & superpage_hits_0; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  hitsVec_3 = vm_enabled & superpage_hits_1; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire [26:0] _hitsVec_T_42 = special_entry_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  _hitsVec_T_56 = special_entry_valid_0 & _hitsVec_T_42[26:18] == 9'h0 & (mpu_ppn_ignore | _hitsVec_T_42[17:9] == 9'h0
    ) & (mpu_ppn_ignore_1 | _hitsVec_T_42[8:0] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire  hitsVec_4 = vm_enabled & _hitsVec_T_56; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire [4:0] real_hits = {hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[src/main/scala/util/package.scala 37:27]
  wire  _hits_T = ~vm_enabled; // @[src/main/scala/rocket/TLB.scala 434:18]
  wire [5:0] hits = {_hits_T,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[src/main/scala/rocket/TLB.scala 434:17]
  wire  line_541_clock;
  wire  line_541_reset;
  wire  line_541_valid;
  reg  line_541_valid_reg;
  wire  newEntry_g = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/TLB.scala 445:25]
  wire  _newEntry_sr_T_4 = io_ptw_resp_bits_pte_v & (io_ptw_resp_bits_pte_r | io_ptw_resp_bits_pte_x & ~
    io_ptw_resp_bits_pte_w) & io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/PTW.scala 141:52]
  wire  newEntry_sr = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/PTW.scala 149:35]
  wire  newEntry_sw = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_w & io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/PTW.scala 151:40]
  wire  newEntry_sx = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/PTW.scala 153:35]
  wire  _T = ~io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/TLB.scala 466:39]
  wire  line_542_clock;
  wire  line_542_reset;
  wire  line_542_valid;
  reg  line_542_valid_reg;
  wire [10:0] special_entry_data_0_lo = {2'h3,cacheable,legal_address,legal_address,cacheable,3'h0,cacheable,1'h0}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire [5:0] special_entry_data_0_hi_lo = {io_ptw_resp_bits_pf,1'h0,newEntry_sw,newEntry_sx,newEntry_sr,1'h1}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire [41:0] _special_entry_data_0_T = {refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae_ptw,
    io_ptw_resp_bits_ae_final,1'h0,special_entry_data_0_hi_lo,special_entry_data_0_lo}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire  line_543_clock;
  wire  line_543_reset;
  wire  line_543_valid;
  reg  line_543_valid_reg;
  wire  _T_2 = io_ptw_resp_bits_level < 2'h2; // @[src/main/scala/rocket/TLB.scala 468:40]
  wire  line_544_clock;
  wire  line_544_reset;
  wire  line_544_valid;
  reg  line_544_valid_reg;
  wire  _T_3 = ~r_superpage_repl_addr; // @[src/main/scala/rocket/TLB.scala 470:82]
  wire  line_545_clock;
  wire  line_545_reset;
  wire  line_545_valid;
  reg  line_545_valid_reg;
  wire  line_546_clock;
  wire  line_546_reset;
  wire  line_546_valid;
  reg  line_546_valid_reg;
  wire  _GEN_153 = invalidate_refill ? 1'h0 : 1'h1; // @[src/main/scala/rocket/TLB.scala 206:16 472:34 210:46]
  wire  _GEN_157 = ~r_superpage_repl_addr ? _GEN_153 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 470:91]
  wire  line_547_clock;
  wire  line_547_reset;
  wire  line_547_valid;
  reg  line_547_valid_reg;
  wire  line_548_clock;
  wire  line_548_reset;
  wire  line_548_valid;
  reg  line_548_valid_reg;
  wire  _GEN_162 = r_superpage_repl_addr ? _GEN_153 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 470:91]
  wire  line_549_clock;
  wire  line_549_reset;
  wire  line_549_valid;
  reg  line_549_valid_reg;
  wire  waddr_1 = r_sectored_hit_valid ? r_sectored_hit_bits : r_sectored_repl_addr; // @[src/main/scala/rocket/TLB.scala 477:22]
  wire  _T_5 = ~waddr_1; // @[src/main/scala/rocket/TLB.scala 478:75]
  wire  line_550_clock;
  wire  line_550_reset;
  wire  line_550_valid;
  reg  line_550_valid_reg;
  wire  _T_6 = ~r_sectored_hit_valid; // @[src/main/scala/rocket/TLB.scala 479:15]
  wire  line_551_clock;
  wire  line_551_reset;
  wire  line_551_valid;
  reg  line_551_valid_reg;
  wire  _GEN_164 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_165 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_166 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_167 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire [1:0] idx = r_refill_tag[1:0]; // @[src/main/scala/util/package.scala 155:13]
  wire  line_552_clock;
  wire  line_552_reset;
  wire  line_552_valid;
  reg  line_552_valid_reg;
  wire  _GEN_168 = 2'h0 == idx | _GEN_164; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_553_clock;
  wire  line_553_reset;
  wire  line_553_valid;
  reg  line_553_valid_reg;
  wire  _GEN_169 = 2'h1 == idx | _GEN_165; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_554_clock;
  wire  line_554_reset;
  wire  line_554_valid;
  reg  line_554_valid_reg;
  wire  _GEN_170 = 2'h2 == idx | _GEN_166; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_555_clock;
  wire  line_555_reset;
  wire  line_555_valid;
  reg  line_555_valid_reg;
  wire  _GEN_171 = 2'h3 == idx | _GEN_167; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_556_clock;
  wire  line_556_reset;
  wire  line_556_valid;
  reg  line_556_valid_reg;
  wire [41:0] _GEN_172 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_557_clock;
  wire  line_557_reset;
  wire  line_557_valid;
  reg  line_557_valid_reg;
  wire [41:0] _GEN_173 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_1; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_558_clock;
  wire  line_558_reset;
  wire  line_558_valid;
  reg  line_558_valid_reg;
  wire [41:0] _GEN_174 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_2; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_559_clock;
  wire  line_559_reset;
  wire  line_559_valid;
  reg  line_559_valid_reg;
  wire [41:0] _GEN_175 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_3; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_560_clock;
  wire  line_560_reset;
  wire  line_560_valid;
  reg  line_560_valid_reg;
  wire  _GEN_176 = invalidate_refill ? 1'h0 : _GEN_168; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_177 = invalidate_refill ? 1'h0 : _GEN_169; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_178 = invalidate_refill ? 1'h0 : _GEN_170; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_179 = invalidate_refill ? 1'h0 : _GEN_171; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_180 = ~waddr_1 ? _GEN_176 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_181 = ~waddr_1 ? _GEN_177 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_182 = ~waddr_1 ? _GEN_178 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_183 = ~waddr_1 ? _GEN_179 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  line_561_clock;
  wire  line_561_reset;
  wire  line_561_valid;
  reg  line_561_valid_reg;
  wire  line_562_clock;
  wire  line_562_reset;
  wire  line_562_valid;
  reg  line_562_valid_reg;
  wire  _GEN_191 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_192 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_193 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_194 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  line_563_clock;
  wire  line_563_reset;
  wire  line_563_valid;
  reg  line_563_valid_reg;
  wire  _GEN_195 = 2'h0 == idx | _GEN_191; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_564_clock;
  wire  line_564_reset;
  wire  line_564_valid;
  reg  line_564_valid_reg;
  wire  _GEN_196 = 2'h1 == idx | _GEN_192; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_565_clock;
  wire  line_565_reset;
  wire  line_565_valid;
  reg  line_565_valid_reg;
  wire  _GEN_197 = 2'h2 == idx | _GEN_193; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_566_clock;
  wire  line_566_reset;
  wire  line_566_valid;
  reg  line_566_valid_reg;
  wire  _GEN_198 = 2'h3 == idx | _GEN_194; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_567_clock;
  wire  line_567_reset;
  wire  line_567_valid;
  reg  line_567_valid_reg;
  wire [41:0] _GEN_199 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_568_clock;
  wire  line_568_reset;
  wire  line_568_valid;
  reg  line_568_valid_reg;
  wire [41:0] _GEN_200 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_1; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_569_clock;
  wire  line_569_reset;
  wire  line_569_valid;
  reg  line_569_valid_reg;
  wire [41:0] _GEN_201 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_2; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_570_clock;
  wire  line_570_reset;
  wire  line_570_valid;
  reg  line_570_valid_reg;
  wire [41:0] _GEN_202 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_3; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_571_clock;
  wire  line_571_reset;
  wire  line_571_valid;
  reg  line_571_valid_reg;
  wire  _GEN_203 = invalidate_refill ? 1'h0 : _GEN_195; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_204 = invalidate_refill ? 1'h0 : _GEN_196; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_205 = invalidate_refill ? 1'h0 : _GEN_197; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_206 = invalidate_refill ? 1'h0 : _GEN_198; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_207 = waddr_1 ? _GEN_203 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_208 = waddr_1 ? _GEN_204 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_209 = waddr_1 ? _GEN_205 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_210 = waddr_1 ? _GEN_206 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_221 = io_ptw_resp_bits_level < 2'h2 ? _GEN_157 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 468:58]
  wire  _GEN_226 = io_ptw_resp_bits_level < 2'h2 ? _GEN_162 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 468:58]
  wire  _GEN_228 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_0 : _GEN_180; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_229 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_1 : _GEN_181; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_230 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_2 : _GEN_182; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_231 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_3 : _GEN_183; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_239 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_0 : _GEN_207; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_240 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_1 : _GEN_208; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_241 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_2 : _GEN_209; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_242 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_3 : _GEN_210; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_253 = ~io_ptw_resp_bits_homogeneous | special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 206:16 335:56 466:70]
  wire  _GEN_258 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_0_valid_0 : _GEN_221; // @[src/main/scala/rocket/TLB.scala 330:30 466:70]
  wire  _GEN_263 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_1_valid_0 : _GEN_226; // @[src/main/scala/rocket/TLB.scala 330:30 466:70]
  wire  _GEN_265 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_0 : _GEN_228; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_266 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_1 : _GEN_229; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_267 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_2 : _GEN_230; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_268 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_3 : _GEN_231; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_276 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_0 : _GEN_239; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_277 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_1 : _GEN_240; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_278 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_2 : _GEN_241; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_279 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_3 : _GEN_242; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_290 = io_ptw_resp_valid ? _GEN_253 : special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 335:56]
  wire  _GEN_295 = io_ptw_resp_valid ? _GEN_258 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 330:30]
  wire  _GEN_300 = io_ptw_resp_valid ? _GEN_263 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 330:30]
  wire  _GEN_302 = io_ptw_resp_valid ? _GEN_265 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_303 = io_ptw_resp_valid ? _GEN_266 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_304 = io_ptw_resp_valid ? _GEN_267 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_305 = io_ptw_resp_valid ? _GEN_268 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_313 = io_ptw_resp_valid ? _GEN_276 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_314 = io_ptw_resp_valid ? _GEN_277 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_315 = io_ptw_resp_valid ? _GEN_278 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_316 = io_ptw_resp_valid ? _GEN_279 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  line_572_clock;
  wire  line_572_reset;
  wire  line_572_valid;
  reg  line_572_valid_reg;
  wire  line_573_clock;
  wire  line_573_reset;
  wire  line_573_valid;
  reg  line_573_valid_reg;
  wire [41:0] _GEN_328 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_data_1 : sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_574_clock;
  wire  line_574_reset;
  wire  line_574_valid;
  reg  line_574_valid_reg;
  wire [41:0] _GEN_329 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_data_2 : _GEN_328; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_575_clock;
  wire  line_575_reset;
  wire  line_575_valid;
  reg  line_575_valid_reg;
  wire [41:0] _GEN_330 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_data_3 : _GEN_329; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_576_clock;
  wire  line_576_reset;
  wire  line_576_valid;
  reg  line_576_valid_reg;
  wire  line_577_clock;
  wire  line_577_reset;
  wire  line_577_valid;
  reg  line_577_valid_reg;
  wire [41:0] _GEN_332 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_data_1 : sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_578_clock;
  wire  line_578_reset;
  wire  line_578_valid;
  reg  line_578_valid_reg;
  wire [41:0] _GEN_333 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_data_2 : _GEN_332; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_579_clock;
  wire  line_579_reset;
  wire  line_579_valid;
  reg  line_579_valid_reg;
  wire [41:0] _GEN_334 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_data_3 : _GEN_333; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire [1:0] ppn_res = entries_barrier_2_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _ppn_T_1 = superpage_hits_ignore_1 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_498 = {{7'd0}, entries_barrier_2_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_2 = _ppn_T_1 | _GEN_498; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_6 = vpn | _GEN_498; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_8 = {ppn_res,_ppn_T_2[17:9],_ppn_T_6[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [1:0] ppn_res_1 = entries_barrier_3_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _ppn_T_9 = superpage_hits_ignore_4 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_500 = {{7'd0}, entries_barrier_3_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_10 = _ppn_T_9 | _GEN_500; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_14 = vpn | _GEN_500; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_16 = {ppn_res_1,_ppn_T_10[17:9],_ppn_T_14[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [1:0] ppn_res_2 = entries_barrier_4_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _GEN_502 = {{7'd0}, entries_barrier_4_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_18 = _mpu_ppn_T_24 | _GEN_502; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_22 = _mpu_ppn_T_28 | _GEN_502; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_24 = {ppn_res_2,_ppn_T_18[17:9],_ppn_T_22[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [19:0] _ppn_T_26 = hitsVec_0 ? entries_barrier_io_y_ppn : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_27 = hitsVec_1 ? entries_barrier_1_io_y_ppn : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_28 = hitsVec_2 ? _ppn_T_8 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_29 = hitsVec_3 ? _ppn_T_16 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_30 = hitsVec_4 ? _ppn_T_24 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_31 = _hits_T ? vpn[19:0] : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_32 = _ppn_T_26 | _ppn_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_33 = _ppn_T_32 | _ppn_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_34 = _ppn_T_33 | _ppn_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_35 = _ppn_T_34 | _ppn_T_30; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] ppn = _ppn_T_35 | _ppn_T_31; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [5:0] ptw_ae_array = {1'h0,entries_barrier_4_io_y_ae_ptw,entries_barrier_3_io_y_ae_ptw,
    entries_barrier_2_io_y_ae_ptw,entries_barrier_1_io_y_ae_ptw,entries_barrier_io_y_ae_ptw}; // @[src/main/scala/rocket/TLB.scala 498:25]
  wire [5:0] final_ae_array = {1'h0,entries_barrier_4_io_y_ae_final,entries_barrier_3_io_y_ae_final,
    entries_barrier_2_io_y_ae_final,entries_barrier_1_io_y_ae_final,entries_barrier_io_y_ae_final}; // @[src/main/scala/rocket/TLB.scala 499:27]
  wire [5:0] ptw_pf_array = {1'h0,entries_barrier_4_io_y_pf,entries_barrier_3_io_y_pf,entries_barrier_2_io_y_pf,
    entries_barrier_1_io_y_pf,entries_barrier_io_y_pf}; // @[src/main/scala/rocket/TLB.scala 500:25]
  wire [5:0] ptw_gf_array = {1'h0,entries_barrier_4_io_y_gf,entries_barrier_3_io_y_gf,entries_barrier_2_io_y_gf,
    entries_barrier_1_io_y_gf,entries_barrier_io_y_gf}; // @[src/main/scala/rocket/TLB.scala 501:25]
  wire [4:0] _priv_rw_ok_T_2 = {entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,
    entries_barrier_1_io_y_u,entries_barrier_io_y_u}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _priv_rw_ok_T_3 = ~priv_s | io_ptw_status_sum ? _priv_rw_ok_T_2 : 5'h0; // @[src/main/scala/rocket/TLB.scala 505:23]
  wire [4:0] _priv_rw_ok_T_5 = ~_priv_rw_ok_T_2; // @[src/main/scala/rocket/TLB.scala 505:84]
  wire [4:0] _priv_rw_ok_T_6 = priv_s ? _priv_rw_ok_T_5 : 5'h0; // @[src/main/scala/rocket/TLB.scala 505:75]
  wire [4:0] priv_rw_ok = _priv_rw_ok_T_3 | _priv_rw_ok_T_6; // @[src/main/scala/rocket/TLB.scala 505:70]
  wire [4:0] _r_array_T = {entries_barrier_4_io_y_sr,entries_barrier_3_io_y_sr,entries_barrier_2_io_y_sr,
    entries_barrier_1_io_y_sr,entries_barrier_io_y_sr}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _r_array_T_1 = {entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,
    entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _r_array_T_2 = io_ptw_status_mxr ? _r_array_T_1 : 5'h0; // @[src/main/scala/rocket/TLB.scala 512:74]
  wire [4:0] _r_array_T_3 = _r_array_T | _r_array_T_2; // @[src/main/scala/rocket/TLB.scala 512:69]
  wire [4:0] _r_array_T_4 = priv_rw_ok & _r_array_T_3; // @[src/main/scala/rocket/TLB.scala 512:41]
  wire [5:0] r_array = {1'h1,_r_array_T_4}; // @[src/main/scala/rocket/TLB.scala 512:20]
  wire [4:0] _w_array_T = {entries_barrier_4_io_y_sw,entries_barrier_3_io_y_sw,entries_barrier_2_io_y_sw,
    entries_barrier_1_io_y_sw,entries_barrier_io_y_sw}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _w_array_T_1 = priv_rw_ok & _w_array_T; // @[src/main/scala/rocket/TLB.scala 513:41]
  wire [5:0] w_array = {1'h1,_w_array_T_1}; // @[src/main/scala/rocket/TLB.scala 513:20]
  wire [1:0] _pr_array_T = legal_address ? 2'h3 : 2'h0; // @[src/main/scala/rocket/TLB.scala 521:26]
  wire [5:0] _pr_array_T_2 = {_pr_array_T,entries_barrier_3_io_y_pr,entries_barrier_2_io_y_pr,entries_barrier_1_io_y_pr,
    entries_barrier_io_y_pr}; // @[src/main/scala/rocket/TLB.scala 521:21]
  wire [5:0] _pr_array_T_3 = ptw_ae_array | final_ae_array; // @[src/main/scala/rocket/TLB.scala 521:104]
  wire [5:0] _pr_array_T_4 = ~_pr_array_T_3; // @[src/main/scala/rocket/TLB.scala 521:89]
  wire [5:0] pr_array = _pr_array_T_2 & _pr_array_T_4; // @[src/main/scala/rocket/TLB.scala 521:87]
  wire [1:0] _pw_array_T = cacheable ? 2'h3 : 2'h0; // @[src/main/scala/rocket/TLB.scala 523:26]
  wire [5:0] _pw_array_T_2 = {_pw_array_T,entries_barrier_3_io_y_pw,entries_barrier_2_io_y_pw,entries_barrier_1_io_y_pw,
    entries_barrier_io_y_pw}; // @[src/main/scala/rocket/TLB.scala 523:21]
  wire [5:0] pw_array = _pw_array_T_2 & _pr_array_T_4; // @[src/main/scala/rocket/TLB.scala 523:87]
  wire [5:0] eff_array = {2'h0,entries_barrier_3_io_y_eff,entries_barrier_2_io_y_eff,entries_barrier_1_io_y_eff,
    entries_barrier_io_y_eff}; // @[src/main/scala/rocket/TLB.scala 527:22]
  wire [5:0] c_array = {_pw_array_T,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,
    entries_barrier_io_y_c}; // @[src/main/scala/rocket/TLB.scala 529:20]
  wire [5:0] ppp_array = {_pw_array_T,entries_barrier_3_io_y_ppp,entries_barrier_2_io_y_ppp,entries_barrier_1_io_y_ppp,
    entries_barrier_io_y_ppp}; // @[src/main/scala/rocket/TLB.scala 531:22]
  wire [5:0] paa_array = {2'h0,entries_barrier_3_io_y_paa,entries_barrier_2_io_y_paa,entries_barrier_1_io_y_paa,
    entries_barrier_io_y_paa}; // @[src/main/scala/rocket/TLB.scala 533:22]
  wire [5:0] pal_array = {2'h0,entries_barrier_3_io_y_pal,entries_barrier_2_io_y_pal,entries_barrier_1_io_y_pal,
    entries_barrier_io_y_pal}; // @[src/main/scala/rocket/TLB.scala 535:22]
  wire [5:0] ppp_array_if_cached = ppp_array | c_array; // @[src/main/scala/rocket/TLB.scala 536:39]
  wire [5:0] paa_array_if_cached = paa_array | c_array; // @[src/main/scala/rocket/TLB.scala 537:39]
  wire [5:0] pal_array_if_cached = pal_array | c_array; // @[src/main/scala/rocket/TLB.scala 538:39]
  wire [3:0] _misaligned_T = 4'h1 << io_req_bits_size; // @[src/main/scala/chisel3/util/OneHot.scala 58:35]
  wire [3:0] _misaligned_T_2 = _misaligned_T - 4'h1; // @[src/main/scala/rocket/TLB.scala 542:69]
  wire [39:0] _GEN_504 = {{36'd0}, _misaligned_T_2}; // @[src/main/scala/rocket/TLB.scala 542:39]
  wire [39:0] _misaligned_T_3 = io_req_bits_vaddr & _GEN_504; // @[src/main/scala/rocket/TLB.scala 542:39]
  wire  misaligned = |_misaligned_T_3; // @[src/main/scala/rocket/TLB.scala 542:77]
  wire [39:0] bad_va_maskedVAddr = io_req_bits_vaddr & 40'hc000000000; // @[src/main/scala/rocket/TLB.scala 551:43]
  wire  _bad_va_T_6 = ~(bad_va_maskedVAddr == 40'h0 | bad_va_maskedVAddr == 40'hc000000000); // @[src/main/scala/rocket/TLB.scala 552:37]
  wire  bad_va = vm_enabled & stage1_en & _bad_va_T_6; // @[src/main/scala/rocket/TLB.scala 560:34]
  wire  _cmd_lrsc_T = io_req_bits_cmd == 5'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_lrsc_T_1 = io_req_bits_cmd == 5'h7; // @[src/main/scala/util/package.scala 16:47]
  wire  cmd_lrsc = _cmd_lrsc_T | _cmd_lrsc_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  _cmd_amo_logical_T = io_req_bits_cmd == 5'h4; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_logical_T_1 = io_req_bits_cmd == 5'h9; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_logical_T_2 = io_req_bits_cmd == 5'ha; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_logical_T_3 = io_req_bits_cmd == 5'hb; // @[src/main/scala/util/package.scala 16:47]
  wire  cmd_amo_logical = _cmd_amo_logical_T | _cmd_amo_logical_T_1 | _cmd_amo_logical_T_2 | _cmd_amo_logical_T_3; // @[src/main/scala/util/package.scala 73:59]
  wire  _cmd_amo_arithmetic_T = io_req_bits_cmd == 5'h8; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_arithmetic_T_1 = io_req_bits_cmd == 5'hc; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_arithmetic_T_2 = io_req_bits_cmd == 5'hd; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_arithmetic_T_3 = io_req_bits_cmd == 5'he; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_amo_arithmetic_T_4 = io_req_bits_cmd == 5'hf; // @[src/main/scala/util/package.scala 16:47]
  wire  cmd_amo_arithmetic = _cmd_amo_arithmetic_T | _cmd_amo_arithmetic_T_1 | _cmd_amo_arithmetic_T_2 |
    _cmd_amo_arithmetic_T_3 | _cmd_amo_arithmetic_T_4; // @[src/main/scala/util/package.scala 73:59]
  wire  cmd_put_partial = io_req_bits_cmd == 5'h11; // @[src/main/scala/rocket/TLB.scala 565:41]
  wire  _cmd_read_T = io_req_bits_cmd == 5'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_read_T_1 = io_req_bits_cmd == 5'h10; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_read_T_6 = _cmd_read_T | _cmd_read_T_1 | _cmd_lrsc_T | _cmd_lrsc_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  _cmd_read_T_23 = cmd_amo_logical | cmd_amo_arithmetic; // @[src/main/scala/rocket/Consts.scala 83:44]
  wire  cmd_read = _cmd_read_T_6 | _cmd_read_T_23; // @[src/main/scala/rocket/Consts.scala 85:68]
  wire  cmd_write = io_req_bits_cmd == 5'h1 | cmd_put_partial | _cmd_lrsc_T_1 | _cmd_read_T_23; // @[src/main/scala/rocket/Consts.scala 86:76]
  wire  _cmd_write_perms_T = io_req_bits_cmd == 5'h5; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_write_perms_T_1 = io_req_bits_cmd == 5'h17; // @[src/main/scala/util/package.scala 16:47]
  wire  _cmd_write_perms_T_2 = _cmd_write_perms_T | _cmd_write_perms_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  cmd_write_perms = cmd_write | _cmd_write_perms_T_2; // @[src/main/scala/rocket/TLB.scala 569:35]
  wire [5:0] _ae_array_T = misaligned ? eff_array : 6'h0; // @[src/main/scala/rocket/TLB.scala 574:8]
  wire [5:0] _ae_array_T_1 = ~c_array; // @[src/main/scala/rocket/TLB.scala 575:19]
  wire [5:0] _ae_array_T_2 = cmd_lrsc ? _ae_array_T_1 : 6'h0; // @[src/main/scala/rocket/TLB.scala 575:8]
  wire [5:0] ae_array = _ae_array_T | _ae_array_T_2; // @[src/main/scala/rocket/TLB.scala 574:37]
  wire [5:0] _ae_ld_array_T = ~pr_array; // @[src/main/scala/rocket/TLB.scala 578:46]
  wire [5:0] _ae_ld_array_T_1 = ae_array | _ae_ld_array_T; // @[src/main/scala/rocket/TLB.scala 578:44]
  wire [5:0] ae_ld_array = cmd_read ? _ae_ld_array_T_1 : 6'h0; // @[src/main/scala/rocket/TLB.scala 578:24]
  wire [5:0] _ae_st_array_T = ~pw_array; // @[src/main/scala/rocket/TLB.scala 580:37]
  wire [5:0] _ae_st_array_T_1 = ae_array | _ae_st_array_T; // @[src/main/scala/rocket/TLB.scala 580:35]
  wire [5:0] _ae_st_array_T_2 = cmd_write_perms ? _ae_st_array_T_1 : 6'h0; // @[src/main/scala/rocket/TLB.scala 580:8]
  wire [5:0] _ae_st_array_T_3 = ~ppp_array_if_cached; // @[src/main/scala/rocket/TLB.scala 581:26]
  wire [5:0] _ae_st_array_T_4 = cmd_put_partial ? _ae_st_array_T_3 : 6'h0; // @[src/main/scala/rocket/TLB.scala 581:8]
  wire [5:0] _ae_st_array_T_5 = _ae_st_array_T_2 | _ae_st_array_T_4; // @[src/main/scala/rocket/TLB.scala 580:53]
  wire [5:0] _ae_st_array_T_6 = ~pal_array_if_cached; // @[src/main/scala/rocket/TLB.scala 582:26]
  wire [5:0] _ae_st_array_T_7 = cmd_amo_logical ? _ae_st_array_T_6 : 6'h0; // @[src/main/scala/rocket/TLB.scala 582:8]
  wire [5:0] _ae_st_array_T_8 = _ae_st_array_T_5 | _ae_st_array_T_7; // @[src/main/scala/rocket/TLB.scala 581:53]
  wire [5:0] _ae_st_array_T_9 = ~paa_array_if_cached; // @[src/main/scala/rocket/TLB.scala 583:29]
  wire [5:0] _ae_st_array_T_10 = cmd_amo_arithmetic ? _ae_st_array_T_9 : 6'h0; // @[src/main/scala/rocket/TLB.scala 583:8]
  wire [5:0] ae_st_array = _ae_st_array_T_8 | _ae_st_array_T_10; // @[src/main/scala/rocket/TLB.scala 582:53]
  wire [5:0] _pf_ld_array_T_1 = ~r_array; // @[src/main/scala/rocket/TLB.scala 589:37]
  wire [5:0] _pf_ld_array_T_2 = ~ptw_ae_array; // @[src/main/scala/rocket/TLB.scala 589:73]
  wire [5:0] _pf_ld_array_T_3 = _pf_ld_array_T_1 & _pf_ld_array_T_2; // @[src/main/scala/rocket/TLB.scala 589:71]
  wire [5:0] _pf_ld_array_T_4 = _pf_ld_array_T_3 | ptw_pf_array; // @[src/main/scala/rocket/TLB.scala 589:88]
  wire [5:0] _pf_ld_array_T_5 = ~ptw_gf_array; // @[src/main/scala/rocket/TLB.scala 589:106]
  wire [5:0] _pf_ld_array_T_6 = _pf_ld_array_T_4 & _pf_ld_array_T_5; // @[src/main/scala/rocket/TLB.scala 589:104]
  wire [5:0] pf_ld_array = cmd_read ? _pf_ld_array_T_6 : 6'h0; // @[src/main/scala/rocket/TLB.scala 589:24]
  wire [5:0] _pf_st_array_T = ~w_array; // @[src/main/scala/rocket/TLB.scala 590:44]
  wire [5:0] _pf_st_array_T_2 = _pf_st_array_T & _pf_ld_array_T_2; // @[src/main/scala/rocket/TLB.scala 590:53]
  wire [5:0] _pf_st_array_T_3 = _pf_st_array_T_2 | ptw_pf_array; // @[src/main/scala/rocket/TLB.scala 590:70]
  wire [5:0] _pf_st_array_T_5 = _pf_st_array_T_3 & _pf_ld_array_T_5; // @[src/main/scala/rocket/TLB.scala 590:86]
  wire [5:0] pf_st_array = cmd_write_perms ? _pf_st_array_T_5 : 6'h0; // @[src/main/scala/rocket/TLB.scala 590:24]
  wire  tlb_hit_if_not_gpa_miss = |real_hits; // @[src/main/scala/rocket/TLB.scala 602:43]
  wire  tlb_miss = vm_enabled & ~bad_va & ~tlb_hit_if_not_gpa_miss; // @[src/main/scala/rocket/TLB.scala 605:64]
  reg  state_vec_0; // @[src/main/scala/util/Replacement.scala 374:17]
  reg  state_reg_1; // @[src/main/scala/util/Replacement.scala 168:72]
  wire  _T_9 = io_req_valid & vm_enabled; // @[src/main/scala/rocket/TLB.scala 609:22]
  wire  line_580_clock;
  wire  line_580_reset;
  wire  line_580_valid;
  reg  line_580_valid_reg;
  wire  _T_10 = sector_hits_0 | sector_hits_1; // @[src/main/scala/util/package.scala 73:59]
  wire  line_581_clock;
  wire  line_581_reset;
  wire  line_581_valid;
  reg  line_581_valid_reg;
  wire [1:0] _T_11 = {sector_hits_1,sector_hits_0}; // @[src/main/scala/chisel3/util/OneHot.scala 21:45]
  wire  state_vec_0_touch_way_sized = _T_11[1]; // @[src/main/scala/chisel3/util/CircuitMath.scala 28:8]
  wire  _state_vec_0_T_1 = ~state_vec_0_touch_way_sized; // @[src/main/scala/util/Replacement.scala 218:7]
  wire  _T_13 = superpage_hits_0 | superpage_hits_1; // @[src/main/scala/util/package.scala 73:59]
  wire  line_582_clock;
  wire  line_582_reset;
  wire  line_582_valid;
  reg  line_582_valid_reg;
  wire [1:0] _T_14 = {superpage_hits_1,superpage_hits_0}; // @[src/main/scala/chisel3/util/OneHot.scala 21:45]
  wire  state_reg_touch_way_sized = _T_14[1]; // @[src/main/scala/chisel3/util/CircuitMath.scala 28:8]
  wire  _state_reg_T_1 = ~state_reg_touch_way_sized; // @[src/main/scala/util/Replacement.scala 218:7]
  wire  multipleHits_leftOne = real_hits[0]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_rightOne = real_hits[1]; // @[src/main/scala/util/Misc.scala 182:39]
  wire  multipleHits_leftOne_1 = multipleHits_leftOne | multipleHits_rightOne; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_leftTwo = multipleHits_leftOne & multipleHits_rightOne; // @[src/main/scala/util/Misc.scala 183:61]
  wire  multipleHits_leftOne_2 = real_hits[2]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_leftOne_3 = real_hits[3]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_rightOne_1 = real_hits[4]; // @[src/main/scala/util/Misc.scala 182:39]
  wire  multipleHits_rightOne_2 = multipleHits_leftOne_3 | multipleHits_rightOne_1; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_rightTwo = multipleHits_leftOne_3 & multipleHits_rightOne_1; // @[src/main/scala/util/Misc.scala 183:61]
  wire  multipleHits_rightOne_3 = multipleHits_leftOne_2 | multipleHits_rightOne_2; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_rightTwo_1 = multipleHits_rightTwo | multipleHits_leftOne_2 & multipleHits_rightOne_2; // @[src/main/scala/util/Misc.scala 183:49]
  wire  multipleHits = multipleHits_leftTwo | multipleHits_rightTwo_1 | multipleHits_leftOne_1 & multipleHits_rightOne_3
    ; // @[src/main/scala/util/Misc.scala 183:49]
  wire [5:0] _io_resp_pf_ld_T_1 = pf_ld_array & hits; // @[src/main/scala/rocket/TLB.scala 625:57]
  wire [5:0] _io_resp_pf_st_T_1 = pf_st_array & hits; // @[src/main/scala/rocket/TLB.scala 626:64]
  wire [5:0] _io_resp_ae_ld_T = ae_ld_array & hits; // @[src/main/scala/rocket/TLB.scala 633:33]
  wire [5:0] _io_resp_ae_st_T = ae_st_array & hits; // @[src/main/scala/rocket/TLB.scala 634:33]
  wire [5:0] _io_resp_cacheable_T = c_array & hits; // @[src/main/scala/rocket/TLB.scala 640:33]
  wire  _T_16 = io_ptw_req_ready & io_ptw_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_17 = _T_16 & io_ptw_req_bits_valid; // @[src/main/scala/rocket/TLB.scala 660:26]
  wire  line_583_clock;
  wire  line_583_reset;
  wire  line_583_valid;
  reg  line_583_valid_reg;
  wire  _T_18 = io_req_ready & io_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_19 = _T_18 & tlb_miss; // @[src/main/scala/rocket/TLB.scala 669:23]
  wire  line_584_clock;
  wire  line_584_reset;
  wire  line_584_valid;
  reg  line_584_valid_reg;
  wire [1:0] r_superpage_repl_addr_valids = {superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[src/main/scala/util/package.scala 37:27]
  wire [1:0] _r_superpage_repl_addr_T_2 = ~r_superpage_repl_addr_valids; // @[src/main/scala/rocket/TLB.scala 747:43]
  wire [1:0] r_sectored_repl_addr_valids = {_sector_hits_T_10,_sector_hits_T_2}; // @[src/main/scala/util/package.scala 37:27]
  wire [1:0] _r_sectored_repl_addr_T_2 = ~r_sectored_repl_addr_valids; // @[src/main/scala/rocket/TLB.scala 747:43]
  wire [1:0] _GEN_341 = _T_18 & tlb_miss ? 2'h1 : state; // @[src/main/scala/rocket/TLB.scala 669:36 670:13 341:22]
  wire  line_585_clock;
  wire  line_585_reset;
  wire  line_585_valid;
  reg  line_585_valid_reg;
  wire  line_586_clock;
  wire  line_586_reset;
  wire  line_586_valid;
  reg  line_586_valid_reg;
  wire [1:0] _GEN_352 = io_sfence_valid ? 2'h0 : _GEN_341; // @[src/main/scala/rocket/TLB.scala 691:{21,29}]
  wire  line_587_clock;
  wire  line_587_reset;
  wire  line_587_valid;
  reg  line_587_valid_reg;
  wire [1:0] _state_T = io_sfence_valid ? 2'h3 : 2'h2; // @[src/main/scala/rocket/TLB.scala 694:45]
  wire [1:0] _GEN_353 = io_ptw_req_ready ? _state_T : _GEN_352; // @[src/main/scala/rocket/TLB.scala 694:{31,39}]
  wire  _T_22 = state == 2'h2 & io_sfence_valid; // @[src/main/scala/rocket/TLB.scala 699:28]
  wire  line_588_clock;
  wire  line_588_reset;
  wire  line_588_valid;
  reg  line_588_valid_reg;
  wire  line_589_clock;
  wire  line_589_reset;
  wire  line_589_valid;
  reg  line_589_valid_reg;
  wire  line_590_clock;
  wire  line_590_reset;
  wire  line_590_valid;
  reg  line_590_valid_reg;
  wire  _T_28 = ~reset; // @[src/main/scala/rocket/TLB.scala 709:13]
  wire  line_591_clock;
  wire  line_591_reset;
  wire  line_591_valid;
  reg  line_591_valid_reg;
  wire  _T_29 = ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn); // @[src/main/scala/rocket/TLB.scala 709:13]
  wire  line_592_clock;
  wire  line_592_reset;
  wire  line_592_valid;
  reg  line_592_valid_reg;
  wire  line_593_clock;
  wire  line_593_reset;
  wire  line_593_valid;
  reg  line_593_valid_reg;
  wire  line_594_clock;
  wire  line_594_reset;
  wire  line_594_valid;
  reg  line_594_valid_reg;
  wire  line_595_clock;
  wire  line_595_reset;
  wire  line_595_valid;
  reg  line_595_valid_reg;
  wire  _GEN_358 = _GEN_0 ? 1'h0 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_596_clock;
  wire  line_596_reset;
  wire  line_596_valid;
  reg  line_596_valid_reg;
  wire  _GEN_359 = _GEN_1 ? 1'h0 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_597_clock;
  wire  line_597_reset;
  wire  line_597_valid;
  reg  line_597_valid_reg;
  wire  _GEN_360 = _GEN_2 ? 1'h0 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_598_clock;
  wire  line_598_reset;
  wire  line_598_valid;
  reg  line_598_valid_reg;
  wire  _GEN_361 = _GEN_3 ? 1'h0 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  _GEN_362 = _sector_hits_T_5 ? _GEN_358 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_363 = _sector_hits_T_5 ? _GEN_359 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_364 = _sector_hits_T_5 ? _GEN_360 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_365 = _sector_hits_T_5 ? _GEN_361 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _T_147 = _sector_hits_T_3[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_599_clock;
  wire  line_599_reset;
  wire  line_599_valid;
  reg  line_599_valid_reg;
  wire  line_600_clock;
  wire  line_600_reset;
  wire  line_600_valid;
  reg  line_600_valid_reg;
  wire  _GEN_366 = sectored_entries_0_0_data_0[0] ? 1'h0 : _GEN_362; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_601_clock;
  wire  line_601_reset;
  wire  line_601_valid;
  reg  line_601_valid_reg;
  wire  _GEN_367 = sectored_entries_0_0_data_1[0] ? 1'h0 : _GEN_363; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_602_clock;
  wire  line_602_reset;
  wire  line_602_valid;
  reg  line_602_valid_reg;
  wire  _GEN_368 = sectored_entries_0_0_data_2[0] ? 1'h0 : _GEN_364; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_603_clock;
  wire  line_603_reset;
  wire  line_603_valid;
  reg  line_603_valid_reg;
  wire  _GEN_369 = sectored_entries_0_0_data_3[0] ? 1'h0 : _GEN_365; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_604_clock;
  wire  line_604_reset;
  wire  line_604_valid;
  reg  line_604_valid_reg;
  wire  line_605_clock;
  wire  line_605_reset;
  wire  line_605_valid;
  reg  line_605_valid_reg;
  wire  _T_343 = ~sectored_entries_0_0_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_606_clock;
  wire  line_606_reset;
  wire  line_606_valid;
  reg  line_606_valid_reg;
  wire  _GEN_374 = ~sectored_entries_0_0_data_0[20] ? 1'h0 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_346 = ~sectored_entries_0_0_data_1[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_607_clock;
  wire  line_607_reset;
  wire  line_607_valid;
  reg  line_607_valid_reg;
  wire  _GEN_375 = ~sectored_entries_0_0_data_1[20] ? 1'h0 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_349 = ~sectored_entries_0_0_data_2[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_608_clock;
  wire  line_608_reset;
  wire  line_608_valid;
  reg  line_608_valid_reg;
  wire  _GEN_376 = ~sectored_entries_0_0_data_2[20] ? 1'h0 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_352 = ~sectored_entries_0_0_data_3[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_609_clock;
  wire  line_609_reset;
  wire  line_609_valid;
  reg  line_609_valid_reg;
  wire  _GEN_377 = ~sectored_entries_0_0_data_3[20] ? 1'h0 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_610_clock;
  wire  line_610_reset;
  wire  line_610_valid;
  reg  line_610_valid_reg;
  wire  _GEN_382 = io_sfence_bits_rs2 & _GEN_374; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_383 = io_sfence_bits_rs2 & _GEN_375; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_384 = io_sfence_bits_rs2 & _GEN_376; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_385 = io_sfence_bits_rs2 & _GEN_377; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_611_clock;
  wire  line_611_reset;
  wire  line_611_valid;
  reg  line_611_valid_reg;
  wire  line_612_clock;
  wire  line_612_reset;
  wire  line_612_valid;
  reg  line_612_valid_reg;
  wire  line_613_clock;
  wire  line_613_reset;
  wire  line_613_valid;
  reg  line_613_valid_reg;
  wire  _GEN_390 = _GEN_0 ? 1'h0 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_614_clock;
  wire  line_614_reset;
  wire  line_614_valid;
  reg  line_614_valid_reg;
  wire  _GEN_391 = _GEN_1 ? 1'h0 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_615_clock;
  wire  line_615_reset;
  wire  line_615_valid;
  reg  line_615_valid_reg;
  wire  _GEN_392 = _GEN_2 ? 1'h0 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_616_clock;
  wire  line_616_reset;
  wire  line_616_valid;
  reg  line_616_valid_reg;
  wire  _GEN_393 = _GEN_3 ? 1'h0 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  _GEN_394 = _sector_hits_T_13 ? _GEN_390 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_395 = _sector_hits_T_13 ? _GEN_391 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_396 = _sector_hits_T_13 ? _GEN_392 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_397 = _sector_hits_T_13 ? _GEN_393 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _T_568 = _sector_hits_T_11[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_617_clock;
  wire  line_617_reset;
  wire  line_617_valid;
  reg  line_617_valid_reg;
  wire  line_618_clock;
  wire  line_618_reset;
  wire  line_618_valid;
  reg  line_618_valid_reg;
  wire  _GEN_398 = sectored_entries_0_1_data_0[0] ? 1'h0 : _GEN_394; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_619_clock;
  wire  line_619_reset;
  wire  line_619_valid;
  reg  line_619_valid_reg;
  wire  _GEN_399 = sectored_entries_0_1_data_1[0] ? 1'h0 : _GEN_395; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_620_clock;
  wire  line_620_reset;
  wire  line_620_valid;
  reg  line_620_valid_reg;
  wire  _GEN_400 = sectored_entries_0_1_data_2[0] ? 1'h0 : _GEN_396; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_621_clock;
  wire  line_621_reset;
  wire  line_621_valid;
  reg  line_621_valid_reg;
  wire  _GEN_401 = sectored_entries_0_1_data_3[0] ? 1'h0 : _GEN_397; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_622_clock;
  wire  line_622_reset;
  wire  line_622_valid;
  reg  line_622_valid_reg;
  wire  line_623_clock;
  wire  line_623_reset;
  wire  line_623_valid;
  reg  line_623_valid_reg;
  wire  _T_764 = ~sectored_entries_0_1_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_624_clock;
  wire  line_624_reset;
  wire  line_624_valid;
  reg  line_624_valid_reg;
  wire  _GEN_406 = ~sectored_entries_0_1_data_0[20] ? 1'h0 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_767 = ~sectored_entries_0_1_data_1[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_625_clock;
  wire  line_625_reset;
  wire  line_625_valid;
  reg  line_625_valid_reg;
  wire  _GEN_407 = ~sectored_entries_0_1_data_1[20] ? 1'h0 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_770 = ~sectored_entries_0_1_data_2[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_626_clock;
  wire  line_626_reset;
  wire  line_626_valid;
  reg  line_626_valid_reg;
  wire  _GEN_408 = ~sectored_entries_0_1_data_2[20] ? 1'h0 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_773 = ~sectored_entries_0_1_data_3[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_627_clock;
  wire  line_627_reset;
  wire  line_627_valid;
  reg  line_627_valid_reg;
  wire  _GEN_409 = ~sectored_entries_0_1_data_3[20] ? 1'h0 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_628_clock;
  wire  line_628_reset;
  wire  line_628_valid;
  reg  line_628_valid_reg;
  wire  _GEN_414 = io_sfence_bits_rs2 & _GEN_406; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_415 = io_sfence_bits_rs2 & _GEN_407; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_416 = io_sfence_bits_rs2 & _GEN_408; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_417 = io_sfence_bits_rs2 & _GEN_409; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_629_clock;
  wire  line_629_reset;
  wire  line_629_valid;
  reg  line_629_valid_reg;
  wire  line_630_clock;
  wire  line_630_reset;
  wire  line_630_valid;
  reg  line_630_valid_reg;
  wire  _GEN_422 = superpage_hits_0 ? 1'h0 : _GEN_295; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_891 = _superpage_hits_T[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_631_clock;
  wire  line_631_reset;
  wire  line_631_valid;
  reg  line_631_valid_reg;
  wire  line_632_clock;
  wire  line_632_reset;
  wire  line_632_valid;
  reg  line_632_valid_reg;
  wire  _GEN_423 = superpage_entries_0_data_0[0] ? 1'h0 : _GEN_422; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_633_clock;
  wire  line_633_reset;
  wire  line_633_valid;
  reg  line_633_valid_reg;
  wire  line_634_clock;
  wire  line_634_reset;
  wire  line_634_valid;
  reg  line_634_valid_reg;
  wire  _T_943 = ~superpage_entries_0_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_635_clock;
  wire  line_635_reset;
  wire  line_635_valid;
  reg  line_635_valid_reg;
  wire  _GEN_425 = ~superpage_entries_0_data_0[20] ? 1'h0 : _GEN_295; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_636_clock;
  wire  line_636_reset;
  wire  line_636_valid;
  reg  line_636_valid_reg;
  wire  _GEN_427 = io_sfence_bits_rs2 & _GEN_425; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_637_clock;
  wire  line_637_reset;
  wire  line_637_valid;
  reg  line_637_valid_reg;
  wire  line_638_clock;
  wire  line_638_reset;
  wire  line_638_valid;
  reg  line_638_valid_reg;
  wire  _GEN_429 = superpage_hits_1 ? 1'h0 : _GEN_300; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_989 = _superpage_hits_T_14[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_639_clock;
  wire  line_639_reset;
  wire  line_639_valid;
  reg  line_639_valid_reg;
  wire  line_640_clock;
  wire  line_640_reset;
  wire  line_640_valid;
  reg  line_640_valid_reg;
  wire  _GEN_430 = superpage_entries_1_data_0[0] ? 1'h0 : _GEN_429; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_641_clock;
  wire  line_641_reset;
  wire  line_641_valid;
  reg  line_641_valid_reg;
  wire  line_642_clock;
  wire  line_642_reset;
  wire  line_642_valid;
  reg  line_642_valid_reg;
  wire  _T_1041 = ~superpage_entries_1_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_643_clock;
  wire  line_643_reset;
  wire  line_643_valid;
  reg  line_643_valid_reg;
  wire  _GEN_432 = ~superpage_entries_1_data_0[20] ? 1'h0 : _GEN_300; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_644_clock;
  wire  line_644_reset;
  wire  line_644_valid;
  reg  line_644_valid_reg;
  wire  _GEN_434 = io_sfence_bits_rs2 & _GEN_432; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_645_clock;
  wire  line_645_reset;
  wire  line_645_valid;
  reg  line_645_valid_reg;
  wire  line_646_clock;
  wire  line_646_reset;
  wire  line_646_valid;
  reg  line_646_valid_reg;
  wire  _GEN_436 = _hitsVec_T_56 ? 1'h0 : _GEN_290; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_1087 = _hitsVec_T_42[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_647_clock;
  wire  line_647_reset;
  wire  line_647_valid;
  reg  line_647_valid_reg;
  wire  line_648_clock;
  wire  line_648_reset;
  wire  line_648_valid;
  reg  line_648_valid_reg;
  wire  _GEN_437 = special_entry_data_0[0] ? 1'h0 : _GEN_436; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_649_clock;
  wire  line_649_reset;
  wire  line_649_valid;
  reg  line_649_valid_reg;
  wire  line_650_clock;
  wire  line_650_reset;
  wire  line_650_valid;
  reg  line_650_valid_reg;
  wire  _T_1139 = ~special_entry_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_651_clock;
  wire  line_651_reset;
  wire  line_651_valid;
  reg  line_651_valid_reg;
  wire  _GEN_439 = ~special_entry_data_0[20] ? 1'h0 : _GEN_290; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_652_clock;
  wire  line_652_reset;
  wire  line_652_valid;
  reg  line_652_valid_reg;
  wire  _GEN_441 = io_sfence_bits_rs2 & _GEN_439; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _T_1433 = multipleHits | reset; // @[src/main/scala/rocket/TLB.scala 722:24]
  wire  line_653_clock;
  wire  line_653_reset;
  wire  line_653_valid;
  reg  line_653_valid_reg;
  OptimizationBarrier mpu_ppn_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(mpu_ppn_barrier_clock),
    .reset(mpu_ppn_barrier_reset),
    .io_x_ppn(mpu_ppn_barrier_io_x_ppn),
    .io_y_ppn(mpu_ppn_barrier_io_y_ppn)
  );
  PMPChecker pmp ( // @[src/main/scala/rocket/TLB.scala 405:19]
    .clock(pmp_clock),
    .reset(pmp_reset)
  );
  OptimizationBarrier_1 entries_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_clock),
    .reset(entries_barrier_reset),
    .io_x_ppn(entries_barrier_io_x_ppn),
    .io_x_u(entries_barrier_io_x_u),
    .io_x_ae_ptw(entries_barrier_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_io_x_ae_final),
    .io_x_pf(entries_barrier_io_x_pf),
    .io_x_gf(entries_barrier_io_x_gf),
    .io_x_sw(entries_barrier_io_x_sw),
    .io_x_sx(entries_barrier_io_x_sx),
    .io_x_sr(entries_barrier_io_x_sr),
    .io_x_pw(entries_barrier_io_x_pw),
    .io_x_pr(entries_barrier_io_x_pr),
    .io_x_ppp(entries_barrier_io_x_ppp),
    .io_x_pal(entries_barrier_io_x_pal),
    .io_x_paa(entries_barrier_io_x_paa),
    .io_x_eff(entries_barrier_io_x_eff),
    .io_x_c(entries_barrier_io_x_c),
    .io_y_ppn(entries_barrier_io_y_ppn),
    .io_y_u(entries_barrier_io_y_u),
    .io_y_ae_ptw(entries_barrier_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_io_y_ae_final),
    .io_y_pf(entries_barrier_io_y_pf),
    .io_y_gf(entries_barrier_io_y_gf),
    .io_y_sw(entries_barrier_io_y_sw),
    .io_y_sx(entries_barrier_io_y_sx),
    .io_y_sr(entries_barrier_io_y_sr),
    .io_y_pw(entries_barrier_io_y_pw),
    .io_y_pr(entries_barrier_io_y_pr),
    .io_y_ppp(entries_barrier_io_y_ppp),
    .io_y_pal(entries_barrier_io_y_pal),
    .io_y_paa(entries_barrier_io_y_paa),
    .io_y_eff(entries_barrier_io_y_eff),
    .io_y_c(entries_barrier_io_y_c)
  );
  OptimizationBarrier_2 entries_barrier_1 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_1_clock),
    .reset(entries_barrier_1_reset),
    .io_x_ppn(entries_barrier_1_io_x_ppn),
    .io_x_u(entries_barrier_1_io_x_u),
    .io_x_ae_ptw(entries_barrier_1_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_1_io_x_ae_final),
    .io_x_pf(entries_barrier_1_io_x_pf),
    .io_x_gf(entries_barrier_1_io_x_gf),
    .io_x_sw(entries_barrier_1_io_x_sw),
    .io_x_sx(entries_barrier_1_io_x_sx),
    .io_x_sr(entries_barrier_1_io_x_sr),
    .io_x_pw(entries_barrier_1_io_x_pw),
    .io_x_pr(entries_barrier_1_io_x_pr),
    .io_x_ppp(entries_barrier_1_io_x_ppp),
    .io_x_pal(entries_barrier_1_io_x_pal),
    .io_x_paa(entries_barrier_1_io_x_paa),
    .io_x_eff(entries_barrier_1_io_x_eff),
    .io_x_c(entries_barrier_1_io_x_c),
    .io_y_ppn(entries_barrier_1_io_y_ppn),
    .io_y_u(entries_barrier_1_io_y_u),
    .io_y_ae_ptw(entries_barrier_1_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_1_io_y_ae_final),
    .io_y_pf(entries_barrier_1_io_y_pf),
    .io_y_gf(entries_barrier_1_io_y_gf),
    .io_y_sw(entries_barrier_1_io_y_sw),
    .io_y_sx(entries_barrier_1_io_y_sx),
    .io_y_sr(entries_barrier_1_io_y_sr),
    .io_y_pw(entries_barrier_1_io_y_pw),
    .io_y_pr(entries_barrier_1_io_y_pr),
    .io_y_ppp(entries_barrier_1_io_y_ppp),
    .io_y_pal(entries_barrier_1_io_y_pal),
    .io_y_paa(entries_barrier_1_io_y_paa),
    .io_y_eff(entries_barrier_1_io_y_eff),
    .io_y_c(entries_barrier_1_io_y_c)
  );
  OptimizationBarrier_3 entries_barrier_2 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_2_clock),
    .reset(entries_barrier_2_reset),
    .io_x_ppn(entries_barrier_2_io_x_ppn),
    .io_x_u(entries_barrier_2_io_x_u),
    .io_x_ae_ptw(entries_barrier_2_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_2_io_x_ae_final),
    .io_x_pf(entries_barrier_2_io_x_pf),
    .io_x_gf(entries_barrier_2_io_x_gf),
    .io_x_sw(entries_barrier_2_io_x_sw),
    .io_x_sx(entries_barrier_2_io_x_sx),
    .io_x_sr(entries_barrier_2_io_x_sr),
    .io_x_pw(entries_barrier_2_io_x_pw),
    .io_x_pr(entries_barrier_2_io_x_pr),
    .io_x_ppp(entries_barrier_2_io_x_ppp),
    .io_x_pal(entries_barrier_2_io_x_pal),
    .io_x_paa(entries_barrier_2_io_x_paa),
    .io_x_eff(entries_barrier_2_io_x_eff),
    .io_x_c(entries_barrier_2_io_x_c),
    .io_y_ppn(entries_barrier_2_io_y_ppn),
    .io_y_u(entries_barrier_2_io_y_u),
    .io_y_ae_ptw(entries_barrier_2_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_2_io_y_ae_final),
    .io_y_pf(entries_barrier_2_io_y_pf),
    .io_y_gf(entries_barrier_2_io_y_gf),
    .io_y_sw(entries_barrier_2_io_y_sw),
    .io_y_sx(entries_barrier_2_io_y_sx),
    .io_y_sr(entries_barrier_2_io_y_sr),
    .io_y_pw(entries_barrier_2_io_y_pw),
    .io_y_pr(entries_barrier_2_io_y_pr),
    .io_y_ppp(entries_barrier_2_io_y_ppp),
    .io_y_pal(entries_barrier_2_io_y_pal),
    .io_y_paa(entries_barrier_2_io_y_paa),
    .io_y_eff(entries_barrier_2_io_y_eff),
    .io_y_c(entries_barrier_2_io_y_c)
  );
  OptimizationBarrier_4 entries_barrier_3 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_3_clock),
    .reset(entries_barrier_3_reset),
    .io_x_ppn(entries_barrier_3_io_x_ppn),
    .io_x_u(entries_barrier_3_io_x_u),
    .io_x_ae_ptw(entries_barrier_3_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_3_io_x_ae_final),
    .io_x_pf(entries_barrier_3_io_x_pf),
    .io_x_gf(entries_barrier_3_io_x_gf),
    .io_x_sw(entries_barrier_3_io_x_sw),
    .io_x_sx(entries_barrier_3_io_x_sx),
    .io_x_sr(entries_barrier_3_io_x_sr),
    .io_x_pw(entries_barrier_3_io_x_pw),
    .io_x_pr(entries_barrier_3_io_x_pr),
    .io_x_ppp(entries_barrier_3_io_x_ppp),
    .io_x_pal(entries_barrier_3_io_x_pal),
    .io_x_paa(entries_barrier_3_io_x_paa),
    .io_x_eff(entries_barrier_3_io_x_eff),
    .io_x_c(entries_barrier_3_io_x_c),
    .io_y_ppn(entries_barrier_3_io_y_ppn),
    .io_y_u(entries_barrier_3_io_y_u),
    .io_y_ae_ptw(entries_barrier_3_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_3_io_y_ae_final),
    .io_y_pf(entries_barrier_3_io_y_pf),
    .io_y_gf(entries_barrier_3_io_y_gf),
    .io_y_sw(entries_barrier_3_io_y_sw),
    .io_y_sx(entries_barrier_3_io_y_sx),
    .io_y_sr(entries_barrier_3_io_y_sr),
    .io_y_pw(entries_barrier_3_io_y_pw),
    .io_y_pr(entries_barrier_3_io_y_pr),
    .io_y_ppp(entries_barrier_3_io_y_ppp),
    .io_y_pal(entries_barrier_3_io_y_pal),
    .io_y_paa(entries_barrier_3_io_y_paa),
    .io_y_eff(entries_barrier_3_io_y_eff),
    .io_y_c(entries_barrier_3_io_y_c)
  );
  OptimizationBarrier_5 entries_barrier_4 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_4_clock),
    .reset(entries_barrier_4_reset),
    .io_x_ppn(entries_barrier_4_io_x_ppn),
    .io_x_u(entries_barrier_4_io_x_u),
    .io_x_ae_ptw(entries_barrier_4_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_4_io_x_ae_final),
    .io_x_pf(entries_barrier_4_io_x_pf),
    .io_x_gf(entries_barrier_4_io_x_gf),
    .io_x_sw(entries_barrier_4_io_x_sw),
    .io_x_sx(entries_barrier_4_io_x_sx),
    .io_x_sr(entries_barrier_4_io_x_sr),
    .io_y_ppn(entries_barrier_4_io_y_ppn),
    .io_y_u(entries_barrier_4_io_y_u),
    .io_y_ae_ptw(entries_barrier_4_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_4_io_y_ae_final),
    .io_y_pf(entries_barrier_4_io_y_pf),
    .io_y_gf(entries_barrier_4_io_y_gf),
    .io_y_sw(entries_barrier_4_io_y_sw),
    .io_y_sx(entries_barrier_4_io_y_sx),
    .io_y_sr(entries_barrier_4_io_y_sr)
  );
  GEN_w1_line #(.COVER_INDEX(533)) line_533 (
    .clock(line_533_clock),
    .reset(line_533_reset),
    .valid(line_533_valid)
  );
  GEN_w1_line #(.COVER_INDEX(534)) line_534 (
    .clock(line_534_clock),
    .reset(line_534_reset),
    .valid(line_534_valid)
  );
  GEN_w1_line #(.COVER_INDEX(535)) line_535 (
    .clock(line_535_clock),
    .reset(line_535_reset),
    .valid(line_535_valid)
  );
  GEN_w1_line #(.COVER_INDEX(536)) line_536 (
    .clock(line_536_clock),
    .reset(line_536_reset),
    .valid(line_536_valid)
  );
  GEN_w1_line #(.COVER_INDEX(537)) line_537 (
    .clock(line_537_clock),
    .reset(line_537_reset),
    .valid(line_537_valid)
  );
  GEN_w1_line #(.COVER_INDEX(538)) line_538 (
    .clock(line_538_clock),
    .reset(line_538_reset),
    .valid(line_538_valid)
  );
  GEN_w1_line #(.COVER_INDEX(539)) line_539 (
    .clock(line_539_clock),
    .reset(line_539_reset),
    .valid(line_539_valid)
  );
  GEN_w1_line #(.COVER_INDEX(540)) line_540 (
    .clock(line_540_clock),
    .reset(line_540_reset),
    .valid(line_540_valid)
  );
  GEN_w1_line #(.COVER_INDEX(541)) line_541 (
    .clock(line_541_clock),
    .reset(line_541_reset),
    .valid(line_541_valid)
  );
  GEN_w1_line #(.COVER_INDEX(542)) line_542 (
    .clock(line_542_clock),
    .reset(line_542_reset),
    .valid(line_542_valid)
  );
  GEN_w1_line #(.COVER_INDEX(543)) line_543 (
    .clock(line_543_clock),
    .reset(line_543_reset),
    .valid(line_543_valid)
  );
  GEN_w1_line #(.COVER_INDEX(544)) line_544 (
    .clock(line_544_clock),
    .reset(line_544_reset),
    .valid(line_544_valid)
  );
  GEN_w1_line #(.COVER_INDEX(545)) line_545 (
    .clock(line_545_clock),
    .reset(line_545_reset),
    .valid(line_545_valid)
  );
  GEN_w1_line #(.COVER_INDEX(546)) line_546 (
    .clock(line_546_clock),
    .reset(line_546_reset),
    .valid(line_546_valid)
  );
  GEN_w1_line #(.COVER_INDEX(547)) line_547 (
    .clock(line_547_clock),
    .reset(line_547_reset),
    .valid(line_547_valid)
  );
  GEN_w1_line #(.COVER_INDEX(548)) line_548 (
    .clock(line_548_clock),
    .reset(line_548_reset),
    .valid(line_548_valid)
  );
  GEN_w1_line #(.COVER_INDEX(549)) line_549 (
    .clock(line_549_clock),
    .reset(line_549_reset),
    .valid(line_549_valid)
  );
  GEN_w1_line #(.COVER_INDEX(550)) line_550 (
    .clock(line_550_clock),
    .reset(line_550_reset),
    .valid(line_550_valid)
  );
  GEN_w1_line #(.COVER_INDEX(551)) line_551 (
    .clock(line_551_clock),
    .reset(line_551_reset),
    .valid(line_551_valid)
  );
  GEN_w1_line #(.COVER_INDEX(552)) line_552 (
    .clock(line_552_clock),
    .reset(line_552_reset),
    .valid(line_552_valid)
  );
  GEN_w1_line #(.COVER_INDEX(553)) line_553 (
    .clock(line_553_clock),
    .reset(line_553_reset),
    .valid(line_553_valid)
  );
  GEN_w1_line #(.COVER_INDEX(554)) line_554 (
    .clock(line_554_clock),
    .reset(line_554_reset),
    .valid(line_554_valid)
  );
  GEN_w1_line #(.COVER_INDEX(555)) line_555 (
    .clock(line_555_clock),
    .reset(line_555_reset),
    .valid(line_555_valid)
  );
  GEN_w1_line #(.COVER_INDEX(556)) line_556 (
    .clock(line_556_clock),
    .reset(line_556_reset),
    .valid(line_556_valid)
  );
  GEN_w1_line #(.COVER_INDEX(557)) line_557 (
    .clock(line_557_clock),
    .reset(line_557_reset),
    .valid(line_557_valid)
  );
  GEN_w1_line #(.COVER_INDEX(558)) line_558 (
    .clock(line_558_clock),
    .reset(line_558_reset),
    .valid(line_558_valid)
  );
  GEN_w1_line #(.COVER_INDEX(559)) line_559 (
    .clock(line_559_clock),
    .reset(line_559_reset),
    .valid(line_559_valid)
  );
  GEN_w1_line #(.COVER_INDEX(560)) line_560 (
    .clock(line_560_clock),
    .reset(line_560_reset),
    .valid(line_560_valid)
  );
  GEN_w1_line #(.COVER_INDEX(561)) line_561 (
    .clock(line_561_clock),
    .reset(line_561_reset),
    .valid(line_561_valid)
  );
  GEN_w1_line #(.COVER_INDEX(562)) line_562 (
    .clock(line_562_clock),
    .reset(line_562_reset),
    .valid(line_562_valid)
  );
  GEN_w1_line #(.COVER_INDEX(563)) line_563 (
    .clock(line_563_clock),
    .reset(line_563_reset),
    .valid(line_563_valid)
  );
  GEN_w1_line #(.COVER_INDEX(564)) line_564 (
    .clock(line_564_clock),
    .reset(line_564_reset),
    .valid(line_564_valid)
  );
  GEN_w1_line #(.COVER_INDEX(565)) line_565 (
    .clock(line_565_clock),
    .reset(line_565_reset),
    .valid(line_565_valid)
  );
  GEN_w1_line #(.COVER_INDEX(566)) line_566 (
    .clock(line_566_clock),
    .reset(line_566_reset),
    .valid(line_566_valid)
  );
  GEN_w1_line #(.COVER_INDEX(567)) line_567 (
    .clock(line_567_clock),
    .reset(line_567_reset),
    .valid(line_567_valid)
  );
  GEN_w1_line #(.COVER_INDEX(568)) line_568 (
    .clock(line_568_clock),
    .reset(line_568_reset),
    .valid(line_568_valid)
  );
  GEN_w1_line #(.COVER_INDEX(569)) line_569 (
    .clock(line_569_clock),
    .reset(line_569_reset),
    .valid(line_569_valid)
  );
  GEN_w1_line #(.COVER_INDEX(570)) line_570 (
    .clock(line_570_clock),
    .reset(line_570_reset),
    .valid(line_570_valid)
  );
  GEN_w1_line #(.COVER_INDEX(571)) line_571 (
    .clock(line_571_clock),
    .reset(line_571_reset),
    .valid(line_571_valid)
  );
  GEN_w1_line #(.COVER_INDEX(572)) line_572 (
    .clock(line_572_clock),
    .reset(line_572_reset),
    .valid(line_572_valid)
  );
  GEN_w1_line #(.COVER_INDEX(573)) line_573 (
    .clock(line_573_clock),
    .reset(line_573_reset),
    .valid(line_573_valid)
  );
  GEN_w1_line #(.COVER_INDEX(574)) line_574 (
    .clock(line_574_clock),
    .reset(line_574_reset),
    .valid(line_574_valid)
  );
  GEN_w1_line #(.COVER_INDEX(575)) line_575 (
    .clock(line_575_clock),
    .reset(line_575_reset),
    .valid(line_575_valid)
  );
  GEN_w1_line #(.COVER_INDEX(576)) line_576 (
    .clock(line_576_clock),
    .reset(line_576_reset),
    .valid(line_576_valid)
  );
  GEN_w1_line #(.COVER_INDEX(577)) line_577 (
    .clock(line_577_clock),
    .reset(line_577_reset),
    .valid(line_577_valid)
  );
  GEN_w1_line #(.COVER_INDEX(578)) line_578 (
    .clock(line_578_clock),
    .reset(line_578_reset),
    .valid(line_578_valid)
  );
  GEN_w1_line #(.COVER_INDEX(579)) line_579 (
    .clock(line_579_clock),
    .reset(line_579_reset),
    .valid(line_579_valid)
  );
  GEN_w1_line #(.COVER_INDEX(580)) line_580 (
    .clock(line_580_clock),
    .reset(line_580_reset),
    .valid(line_580_valid)
  );
  GEN_w1_line #(.COVER_INDEX(581)) line_581 (
    .clock(line_581_clock),
    .reset(line_581_reset),
    .valid(line_581_valid)
  );
  GEN_w1_line #(.COVER_INDEX(582)) line_582 (
    .clock(line_582_clock),
    .reset(line_582_reset),
    .valid(line_582_valid)
  );
  GEN_w1_line #(.COVER_INDEX(583)) line_583 (
    .clock(line_583_clock),
    .reset(line_583_reset),
    .valid(line_583_valid)
  );
  GEN_w1_line #(.COVER_INDEX(584)) line_584 (
    .clock(line_584_clock),
    .reset(line_584_reset),
    .valid(line_584_valid)
  );
  GEN_w1_line #(.COVER_INDEX(585)) line_585 (
    .clock(line_585_clock),
    .reset(line_585_reset),
    .valid(line_585_valid)
  );
  GEN_w1_line #(.COVER_INDEX(586)) line_586 (
    .clock(line_586_clock),
    .reset(line_586_reset),
    .valid(line_586_valid)
  );
  GEN_w1_line #(.COVER_INDEX(587)) line_587 (
    .clock(line_587_clock),
    .reset(line_587_reset),
    .valid(line_587_valid)
  );
  GEN_w1_line #(.COVER_INDEX(588)) line_588 (
    .clock(line_588_clock),
    .reset(line_588_reset),
    .valid(line_588_valid)
  );
  GEN_w1_line #(.COVER_INDEX(589)) line_589 (
    .clock(line_589_clock),
    .reset(line_589_reset),
    .valid(line_589_valid)
  );
  GEN_w1_line #(.COVER_INDEX(590)) line_590 (
    .clock(line_590_clock),
    .reset(line_590_reset),
    .valid(line_590_valid)
  );
  GEN_w1_line #(.COVER_INDEX(591)) line_591 (
    .clock(line_591_clock),
    .reset(line_591_reset),
    .valid(line_591_valid)
  );
  GEN_w1_line #(.COVER_INDEX(592)) line_592 (
    .clock(line_592_clock),
    .reset(line_592_reset),
    .valid(line_592_valid)
  );
  GEN_w1_line #(.COVER_INDEX(593)) line_593 (
    .clock(line_593_clock),
    .reset(line_593_reset),
    .valid(line_593_valid)
  );
  GEN_w1_line #(.COVER_INDEX(594)) line_594 (
    .clock(line_594_clock),
    .reset(line_594_reset),
    .valid(line_594_valid)
  );
  GEN_w1_line #(.COVER_INDEX(595)) line_595 (
    .clock(line_595_clock),
    .reset(line_595_reset),
    .valid(line_595_valid)
  );
  GEN_w1_line #(.COVER_INDEX(596)) line_596 (
    .clock(line_596_clock),
    .reset(line_596_reset),
    .valid(line_596_valid)
  );
  GEN_w1_line #(.COVER_INDEX(597)) line_597 (
    .clock(line_597_clock),
    .reset(line_597_reset),
    .valid(line_597_valid)
  );
  GEN_w1_line #(.COVER_INDEX(598)) line_598 (
    .clock(line_598_clock),
    .reset(line_598_reset),
    .valid(line_598_valid)
  );
  GEN_w1_line #(.COVER_INDEX(599)) line_599 (
    .clock(line_599_clock),
    .reset(line_599_reset),
    .valid(line_599_valid)
  );
  GEN_w1_line #(.COVER_INDEX(600)) line_600 (
    .clock(line_600_clock),
    .reset(line_600_reset),
    .valid(line_600_valid)
  );
  GEN_w1_line #(.COVER_INDEX(601)) line_601 (
    .clock(line_601_clock),
    .reset(line_601_reset),
    .valid(line_601_valid)
  );
  GEN_w1_line #(.COVER_INDEX(602)) line_602 (
    .clock(line_602_clock),
    .reset(line_602_reset),
    .valid(line_602_valid)
  );
  GEN_w1_line #(.COVER_INDEX(603)) line_603 (
    .clock(line_603_clock),
    .reset(line_603_reset),
    .valid(line_603_valid)
  );
  GEN_w1_line #(.COVER_INDEX(604)) line_604 (
    .clock(line_604_clock),
    .reset(line_604_reset),
    .valid(line_604_valid)
  );
  GEN_w1_line #(.COVER_INDEX(605)) line_605 (
    .clock(line_605_clock),
    .reset(line_605_reset),
    .valid(line_605_valid)
  );
  GEN_w1_line #(.COVER_INDEX(606)) line_606 (
    .clock(line_606_clock),
    .reset(line_606_reset),
    .valid(line_606_valid)
  );
  GEN_w1_line #(.COVER_INDEX(607)) line_607 (
    .clock(line_607_clock),
    .reset(line_607_reset),
    .valid(line_607_valid)
  );
  GEN_w1_line #(.COVER_INDEX(608)) line_608 (
    .clock(line_608_clock),
    .reset(line_608_reset),
    .valid(line_608_valid)
  );
  GEN_w1_line #(.COVER_INDEX(609)) line_609 (
    .clock(line_609_clock),
    .reset(line_609_reset),
    .valid(line_609_valid)
  );
  GEN_w1_line #(.COVER_INDEX(610)) line_610 (
    .clock(line_610_clock),
    .reset(line_610_reset),
    .valid(line_610_valid)
  );
  GEN_w1_line #(.COVER_INDEX(611)) line_611 (
    .clock(line_611_clock),
    .reset(line_611_reset),
    .valid(line_611_valid)
  );
  GEN_w1_line #(.COVER_INDEX(612)) line_612 (
    .clock(line_612_clock),
    .reset(line_612_reset),
    .valid(line_612_valid)
  );
  GEN_w1_line #(.COVER_INDEX(613)) line_613 (
    .clock(line_613_clock),
    .reset(line_613_reset),
    .valid(line_613_valid)
  );
  GEN_w1_line #(.COVER_INDEX(614)) line_614 (
    .clock(line_614_clock),
    .reset(line_614_reset),
    .valid(line_614_valid)
  );
  GEN_w1_line #(.COVER_INDEX(615)) line_615 (
    .clock(line_615_clock),
    .reset(line_615_reset),
    .valid(line_615_valid)
  );
  GEN_w1_line #(.COVER_INDEX(616)) line_616 (
    .clock(line_616_clock),
    .reset(line_616_reset),
    .valid(line_616_valid)
  );
  GEN_w1_line #(.COVER_INDEX(617)) line_617 (
    .clock(line_617_clock),
    .reset(line_617_reset),
    .valid(line_617_valid)
  );
  GEN_w1_line #(.COVER_INDEX(618)) line_618 (
    .clock(line_618_clock),
    .reset(line_618_reset),
    .valid(line_618_valid)
  );
  GEN_w1_line #(.COVER_INDEX(619)) line_619 (
    .clock(line_619_clock),
    .reset(line_619_reset),
    .valid(line_619_valid)
  );
  GEN_w1_line #(.COVER_INDEX(620)) line_620 (
    .clock(line_620_clock),
    .reset(line_620_reset),
    .valid(line_620_valid)
  );
  GEN_w1_line #(.COVER_INDEX(621)) line_621 (
    .clock(line_621_clock),
    .reset(line_621_reset),
    .valid(line_621_valid)
  );
  GEN_w1_line #(.COVER_INDEX(622)) line_622 (
    .clock(line_622_clock),
    .reset(line_622_reset),
    .valid(line_622_valid)
  );
  GEN_w1_line #(.COVER_INDEX(623)) line_623 (
    .clock(line_623_clock),
    .reset(line_623_reset),
    .valid(line_623_valid)
  );
  GEN_w1_line #(.COVER_INDEX(624)) line_624 (
    .clock(line_624_clock),
    .reset(line_624_reset),
    .valid(line_624_valid)
  );
  GEN_w1_line #(.COVER_INDEX(625)) line_625 (
    .clock(line_625_clock),
    .reset(line_625_reset),
    .valid(line_625_valid)
  );
  GEN_w1_line #(.COVER_INDEX(626)) line_626 (
    .clock(line_626_clock),
    .reset(line_626_reset),
    .valid(line_626_valid)
  );
  GEN_w1_line #(.COVER_INDEX(627)) line_627 (
    .clock(line_627_clock),
    .reset(line_627_reset),
    .valid(line_627_valid)
  );
  GEN_w1_line #(.COVER_INDEX(628)) line_628 (
    .clock(line_628_clock),
    .reset(line_628_reset),
    .valid(line_628_valid)
  );
  GEN_w1_line #(.COVER_INDEX(629)) line_629 (
    .clock(line_629_clock),
    .reset(line_629_reset),
    .valid(line_629_valid)
  );
  GEN_w1_line #(.COVER_INDEX(630)) line_630 (
    .clock(line_630_clock),
    .reset(line_630_reset),
    .valid(line_630_valid)
  );
  GEN_w1_line #(.COVER_INDEX(631)) line_631 (
    .clock(line_631_clock),
    .reset(line_631_reset),
    .valid(line_631_valid)
  );
  GEN_w1_line #(.COVER_INDEX(632)) line_632 (
    .clock(line_632_clock),
    .reset(line_632_reset),
    .valid(line_632_valid)
  );
  GEN_w1_line #(.COVER_INDEX(633)) line_633 (
    .clock(line_633_clock),
    .reset(line_633_reset),
    .valid(line_633_valid)
  );
  GEN_w1_line #(.COVER_INDEX(634)) line_634 (
    .clock(line_634_clock),
    .reset(line_634_reset),
    .valid(line_634_valid)
  );
  GEN_w1_line #(.COVER_INDEX(635)) line_635 (
    .clock(line_635_clock),
    .reset(line_635_reset),
    .valid(line_635_valid)
  );
  GEN_w1_line #(.COVER_INDEX(636)) line_636 (
    .clock(line_636_clock),
    .reset(line_636_reset),
    .valid(line_636_valid)
  );
  GEN_w1_line #(.COVER_INDEX(637)) line_637 (
    .clock(line_637_clock),
    .reset(line_637_reset),
    .valid(line_637_valid)
  );
  GEN_w1_line #(.COVER_INDEX(638)) line_638 (
    .clock(line_638_clock),
    .reset(line_638_reset),
    .valid(line_638_valid)
  );
  GEN_w1_line #(.COVER_INDEX(639)) line_639 (
    .clock(line_639_clock),
    .reset(line_639_reset),
    .valid(line_639_valid)
  );
  GEN_w1_line #(.COVER_INDEX(640)) line_640 (
    .clock(line_640_clock),
    .reset(line_640_reset),
    .valid(line_640_valid)
  );
  GEN_w1_line #(.COVER_INDEX(641)) line_641 (
    .clock(line_641_clock),
    .reset(line_641_reset),
    .valid(line_641_valid)
  );
  GEN_w1_line #(.COVER_INDEX(642)) line_642 (
    .clock(line_642_clock),
    .reset(line_642_reset),
    .valid(line_642_valid)
  );
  GEN_w1_line #(.COVER_INDEX(643)) line_643 (
    .clock(line_643_clock),
    .reset(line_643_reset),
    .valid(line_643_valid)
  );
  GEN_w1_line #(.COVER_INDEX(644)) line_644 (
    .clock(line_644_clock),
    .reset(line_644_reset),
    .valid(line_644_valid)
  );
  GEN_w1_line #(.COVER_INDEX(645)) line_645 (
    .clock(line_645_clock),
    .reset(line_645_reset),
    .valid(line_645_valid)
  );
  GEN_w1_line #(.COVER_INDEX(646)) line_646 (
    .clock(line_646_clock),
    .reset(line_646_reset),
    .valid(line_646_valid)
  );
  GEN_w1_line #(.COVER_INDEX(647)) line_647 (
    .clock(line_647_clock),
    .reset(line_647_reset),
    .valid(line_647_valid)
  );
  GEN_w1_line #(.COVER_INDEX(648)) line_648 (
    .clock(line_648_clock),
    .reset(line_648_reset),
    .valid(line_648_valid)
  );
  GEN_w1_line #(.COVER_INDEX(649)) line_649 (
    .clock(line_649_clock),
    .reset(line_649_reset),
    .valid(line_649_valid)
  );
  GEN_w1_line #(.COVER_INDEX(650)) line_650 (
    .clock(line_650_clock),
    .reset(line_650_reset),
    .valid(line_650_valid)
  );
  GEN_w1_line #(.COVER_INDEX(651)) line_651 (
    .clock(line_651_clock),
    .reset(line_651_reset),
    .valid(line_651_valid)
  );
  GEN_w1_line #(.COVER_INDEX(652)) line_652 (
    .clock(line_652_clock),
    .reset(line_652_reset),
    .valid(line_652_valid)
  );
  GEN_w1_line #(.COVER_INDEX(653)) line_653 (
    .clock(line_653_clock),
    .reset(line_653_reset),
    .valid(line_653_valid)
  );
  assign line_533_clock = clock;
  assign line_533_reset = reset;
  assign line_533_valid = 2'h0 == hitsVec_idx ^ line_533_valid_reg;
  assign line_534_clock = clock;
  assign line_534_reset = reset;
  assign line_534_valid = 2'h1 == hitsVec_idx ^ line_534_valid_reg;
  assign line_535_clock = clock;
  assign line_535_reset = reset;
  assign line_535_valid = 2'h2 == hitsVec_idx ^ line_535_valid_reg;
  assign line_536_clock = clock;
  assign line_536_reset = reset;
  assign line_536_valid = 2'h3 == hitsVec_idx ^ line_536_valid_reg;
  assign line_537_clock = clock;
  assign line_537_reset = reset;
  assign line_537_valid = 2'h0 == hitsVec_idx ^ line_537_valid_reg;
  assign line_538_clock = clock;
  assign line_538_reset = reset;
  assign line_538_valid = 2'h1 == hitsVec_idx ^ line_538_valid_reg;
  assign line_539_clock = clock;
  assign line_539_reset = reset;
  assign line_539_valid = 2'h2 == hitsVec_idx ^ line_539_valid_reg;
  assign line_540_clock = clock;
  assign line_540_reset = reset;
  assign line_540_valid = 2'h3 == hitsVec_idx ^ line_540_valid_reg;
  assign line_541_clock = clock;
  assign line_541_reset = reset;
  assign line_541_valid = io_ptw_resp_valid ^ line_541_valid_reg;
  assign line_542_clock = clock;
  assign line_542_reset = reset;
  assign line_542_valid = _T ^ line_542_valid_reg;
  assign line_543_clock = clock;
  assign line_543_reset = reset;
  assign line_543_valid = _T ^ line_543_valid_reg;
  assign line_544_clock = clock;
  assign line_544_reset = reset;
  assign line_544_valid = _T_2 ^ line_544_valid_reg;
  assign line_545_clock = clock;
  assign line_545_reset = reset;
  assign line_545_valid = _T_3 ^ line_545_valid_reg;
  assign line_546_clock = clock;
  assign line_546_reset = reset;
  assign line_546_valid = invalidate_refill ^ line_546_valid_reg;
  assign line_547_clock = clock;
  assign line_547_reset = reset;
  assign line_547_valid = r_superpage_repl_addr ^ line_547_valid_reg;
  assign line_548_clock = clock;
  assign line_548_reset = reset;
  assign line_548_valid = invalidate_refill ^ line_548_valid_reg;
  assign line_549_clock = clock;
  assign line_549_reset = reset;
  assign line_549_valid = _T_2 ^ line_549_valid_reg;
  assign line_550_clock = clock;
  assign line_550_reset = reset;
  assign line_550_valid = _T_5 ^ line_550_valid_reg;
  assign line_551_clock = clock;
  assign line_551_reset = reset;
  assign line_551_valid = _T_6 ^ line_551_valid_reg;
  assign line_552_clock = clock;
  assign line_552_reset = reset;
  assign line_552_valid = 2'h0 == idx ^ line_552_valid_reg;
  assign line_553_clock = clock;
  assign line_553_reset = reset;
  assign line_553_valid = 2'h1 == idx ^ line_553_valid_reg;
  assign line_554_clock = clock;
  assign line_554_reset = reset;
  assign line_554_valid = 2'h2 == idx ^ line_554_valid_reg;
  assign line_555_clock = clock;
  assign line_555_reset = reset;
  assign line_555_valid = 2'h3 == idx ^ line_555_valid_reg;
  assign line_556_clock = clock;
  assign line_556_reset = reset;
  assign line_556_valid = 2'h0 == idx ^ line_556_valid_reg;
  assign line_557_clock = clock;
  assign line_557_reset = reset;
  assign line_557_valid = 2'h1 == idx ^ line_557_valid_reg;
  assign line_558_clock = clock;
  assign line_558_reset = reset;
  assign line_558_valid = 2'h2 == idx ^ line_558_valid_reg;
  assign line_559_clock = clock;
  assign line_559_reset = reset;
  assign line_559_valid = 2'h3 == idx ^ line_559_valid_reg;
  assign line_560_clock = clock;
  assign line_560_reset = reset;
  assign line_560_valid = invalidate_refill ^ line_560_valid_reg;
  assign line_561_clock = clock;
  assign line_561_reset = reset;
  assign line_561_valid = waddr_1 ^ line_561_valid_reg;
  assign line_562_clock = clock;
  assign line_562_reset = reset;
  assign line_562_valid = _T_6 ^ line_562_valid_reg;
  assign line_563_clock = clock;
  assign line_563_reset = reset;
  assign line_563_valid = 2'h0 == idx ^ line_563_valid_reg;
  assign line_564_clock = clock;
  assign line_564_reset = reset;
  assign line_564_valid = 2'h1 == idx ^ line_564_valid_reg;
  assign line_565_clock = clock;
  assign line_565_reset = reset;
  assign line_565_valid = 2'h2 == idx ^ line_565_valid_reg;
  assign line_566_clock = clock;
  assign line_566_reset = reset;
  assign line_566_valid = 2'h3 == idx ^ line_566_valid_reg;
  assign line_567_clock = clock;
  assign line_567_reset = reset;
  assign line_567_valid = 2'h0 == idx ^ line_567_valid_reg;
  assign line_568_clock = clock;
  assign line_568_reset = reset;
  assign line_568_valid = 2'h1 == idx ^ line_568_valid_reg;
  assign line_569_clock = clock;
  assign line_569_reset = reset;
  assign line_569_valid = 2'h2 == idx ^ line_569_valid_reg;
  assign line_570_clock = clock;
  assign line_570_reset = reset;
  assign line_570_valid = 2'h3 == idx ^ line_570_valid_reg;
  assign line_571_clock = clock;
  assign line_571_reset = reset;
  assign line_571_valid = invalidate_refill ^ line_571_valid_reg;
  assign line_572_clock = clock;
  assign line_572_reset = reset;
  assign line_572_valid = 2'h0 == hitsVec_idx ^ line_572_valid_reg;
  assign line_573_clock = clock;
  assign line_573_reset = reset;
  assign line_573_valid = 2'h1 == hitsVec_idx ^ line_573_valid_reg;
  assign line_574_clock = clock;
  assign line_574_reset = reset;
  assign line_574_valid = 2'h2 == hitsVec_idx ^ line_574_valid_reg;
  assign line_575_clock = clock;
  assign line_575_reset = reset;
  assign line_575_valid = 2'h3 == hitsVec_idx ^ line_575_valid_reg;
  assign line_576_clock = clock;
  assign line_576_reset = reset;
  assign line_576_valid = 2'h0 == hitsVec_idx ^ line_576_valid_reg;
  assign line_577_clock = clock;
  assign line_577_reset = reset;
  assign line_577_valid = 2'h1 == hitsVec_idx ^ line_577_valid_reg;
  assign line_578_clock = clock;
  assign line_578_reset = reset;
  assign line_578_valid = 2'h2 == hitsVec_idx ^ line_578_valid_reg;
  assign line_579_clock = clock;
  assign line_579_reset = reset;
  assign line_579_valid = 2'h3 == hitsVec_idx ^ line_579_valid_reg;
  assign line_580_clock = clock;
  assign line_580_reset = reset;
  assign line_580_valid = _T_9 ^ line_580_valid_reg;
  assign line_581_clock = clock;
  assign line_581_reset = reset;
  assign line_581_valid = _T_10 ^ line_581_valid_reg;
  assign line_582_clock = clock;
  assign line_582_reset = reset;
  assign line_582_valid = _T_13 ^ line_582_valid_reg;
  assign line_583_clock = clock;
  assign line_583_reset = reset;
  assign line_583_valid = _T_17 ^ line_583_valid_reg;
  assign line_584_clock = clock;
  assign line_584_reset = reset;
  assign line_584_valid = _T_19 ^ line_584_valid_reg;
  assign line_585_clock = clock;
  assign line_585_reset = reset;
  assign line_585_valid = _invalidate_refill_T ^ line_585_valid_reg;
  assign line_586_clock = clock;
  assign line_586_reset = reset;
  assign line_586_valid = io_sfence_valid ^ line_586_valid_reg;
  assign line_587_clock = clock;
  assign line_587_reset = reset;
  assign line_587_valid = io_ptw_req_ready ^ line_587_valid_reg;
  assign line_588_clock = clock;
  assign line_588_reset = reset;
  assign line_588_valid = _T_22 ^ line_588_valid_reg;
  assign line_589_clock = clock;
  assign line_589_reset = reset;
  assign line_589_valid = io_ptw_resp_valid ^ line_589_valid_reg;
  assign line_590_clock = clock;
  assign line_590_reset = reset;
  assign line_590_valid = io_sfence_valid ^ line_590_valid_reg;
  assign line_591_clock = clock;
  assign line_591_reset = reset;
  assign line_591_valid = _T_28 ^ line_591_valid_reg;
  assign line_592_clock = clock;
  assign line_592_reset = reset;
  assign line_592_valid = _T_29 ^ line_592_valid_reg;
  assign line_593_clock = clock;
  assign line_593_reset = reset;
  assign line_593_valid = io_sfence_bits_rs1 ^ line_593_valid_reg;
  assign line_594_clock = clock;
  assign line_594_reset = reset;
  assign line_594_valid = _sector_hits_T_5 ^ line_594_valid_reg;
  assign line_595_clock = clock;
  assign line_595_reset = reset;
  assign line_595_valid = _GEN_0 ^ line_595_valid_reg;
  assign line_596_clock = clock;
  assign line_596_reset = reset;
  assign line_596_valid = _GEN_1 ^ line_596_valid_reg;
  assign line_597_clock = clock;
  assign line_597_reset = reset;
  assign line_597_valid = _GEN_2 ^ line_597_valid_reg;
  assign line_598_clock = clock;
  assign line_598_reset = reset;
  assign line_598_valid = _GEN_3 ^ line_598_valid_reg;
  assign line_599_clock = clock;
  assign line_599_reset = reset;
  assign line_599_valid = _T_147 ^ line_599_valid_reg;
  assign line_600_clock = clock;
  assign line_600_reset = reset;
  assign line_600_valid = sectored_entries_0_0_data_0[0] ^ line_600_valid_reg;
  assign line_601_clock = clock;
  assign line_601_reset = reset;
  assign line_601_valid = sectored_entries_0_0_data_1[0] ^ line_601_valid_reg;
  assign line_602_clock = clock;
  assign line_602_reset = reset;
  assign line_602_valid = sectored_entries_0_0_data_2[0] ^ line_602_valid_reg;
  assign line_603_clock = clock;
  assign line_603_reset = reset;
  assign line_603_valid = sectored_entries_0_0_data_3[0] ^ line_603_valid_reg;
  assign line_604_clock = clock;
  assign line_604_reset = reset;
  assign line_604_valid = io_sfence_bits_rs1 ^ line_604_valid_reg;
  assign line_605_clock = clock;
  assign line_605_reset = reset;
  assign line_605_valid = io_sfence_bits_rs2 ^ line_605_valid_reg;
  assign line_606_clock = clock;
  assign line_606_reset = reset;
  assign line_606_valid = _T_343 ^ line_606_valid_reg;
  assign line_607_clock = clock;
  assign line_607_reset = reset;
  assign line_607_valid = _T_346 ^ line_607_valid_reg;
  assign line_608_clock = clock;
  assign line_608_reset = reset;
  assign line_608_valid = _T_349 ^ line_608_valid_reg;
  assign line_609_clock = clock;
  assign line_609_reset = reset;
  assign line_609_valid = _T_352 ^ line_609_valid_reg;
  assign line_610_clock = clock;
  assign line_610_reset = reset;
  assign line_610_valid = io_sfence_bits_rs2 ^ line_610_valid_reg;
  assign line_611_clock = clock;
  assign line_611_reset = reset;
  assign line_611_valid = io_sfence_bits_rs1 ^ line_611_valid_reg;
  assign line_612_clock = clock;
  assign line_612_reset = reset;
  assign line_612_valid = _sector_hits_T_13 ^ line_612_valid_reg;
  assign line_613_clock = clock;
  assign line_613_reset = reset;
  assign line_613_valid = _GEN_0 ^ line_613_valid_reg;
  assign line_614_clock = clock;
  assign line_614_reset = reset;
  assign line_614_valid = _GEN_1 ^ line_614_valid_reg;
  assign line_615_clock = clock;
  assign line_615_reset = reset;
  assign line_615_valid = _GEN_2 ^ line_615_valid_reg;
  assign line_616_clock = clock;
  assign line_616_reset = reset;
  assign line_616_valid = _GEN_3 ^ line_616_valid_reg;
  assign line_617_clock = clock;
  assign line_617_reset = reset;
  assign line_617_valid = _T_568 ^ line_617_valid_reg;
  assign line_618_clock = clock;
  assign line_618_reset = reset;
  assign line_618_valid = sectored_entries_0_1_data_0[0] ^ line_618_valid_reg;
  assign line_619_clock = clock;
  assign line_619_reset = reset;
  assign line_619_valid = sectored_entries_0_1_data_1[0] ^ line_619_valid_reg;
  assign line_620_clock = clock;
  assign line_620_reset = reset;
  assign line_620_valid = sectored_entries_0_1_data_2[0] ^ line_620_valid_reg;
  assign line_621_clock = clock;
  assign line_621_reset = reset;
  assign line_621_valid = sectored_entries_0_1_data_3[0] ^ line_621_valid_reg;
  assign line_622_clock = clock;
  assign line_622_reset = reset;
  assign line_622_valid = io_sfence_bits_rs1 ^ line_622_valid_reg;
  assign line_623_clock = clock;
  assign line_623_reset = reset;
  assign line_623_valid = io_sfence_bits_rs2 ^ line_623_valid_reg;
  assign line_624_clock = clock;
  assign line_624_reset = reset;
  assign line_624_valid = _T_764 ^ line_624_valid_reg;
  assign line_625_clock = clock;
  assign line_625_reset = reset;
  assign line_625_valid = _T_767 ^ line_625_valid_reg;
  assign line_626_clock = clock;
  assign line_626_reset = reset;
  assign line_626_valid = _T_770 ^ line_626_valid_reg;
  assign line_627_clock = clock;
  assign line_627_reset = reset;
  assign line_627_valid = _T_773 ^ line_627_valid_reg;
  assign line_628_clock = clock;
  assign line_628_reset = reset;
  assign line_628_valid = io_sfence_bits_rs2 ^ line_628_valid_reg;
  assign line_629_clock = clock;
  assign line_629_reset = reset;
  assign line_629_valid = io_sfence_bits_rs1 ^ line_629_valid_reg;
  assign line_630_clock = clock;
  assign line_630_reset = reset;
  assign line_630_valid = superpage_hits_0 ^ line_630_valid_reg;
  assign line_631_clock = clock;
  assign line_631_reset = reset;
  assign line_631_valid = _T_891 ^ line_631_valid_reg;
  assign line_632_clock = clock;
  assign line_632_reset = reset;
  assign line_632_valid = superpage_entries_0_data_0[0] ^ line_632_valid_reg;
  assign line_633_clock = clock;
  assign line_633_reset = reset;
  assign line_633_valid = io_sfence_bits_rs1 ^ line_633_valid_reg;
  assign line_634_clock = clock;
  assign line_634_reset = reset;
  assign line_634_valid = io_sfence_bits_rs2 ^ line_634_valid_reg;
  assign line_635_clock = clock;
  assign line_635_reset = reset;
  assign line_635_valid = _T_943 ^ line_635_valid_reg;
  assign line_636_clock = clock;
  assign line_636_reset = reset;
  assign line_636_valid = io_sfence_bits_rs2 ^ line_636_valid_reg;
  assign line_637_clock = clock;
  assign line_637_reset = reset;
  assign line_637_valid = io_sfence_bits_rs1 ^ line_637_valid_reg;
  assign line_638_clock = clock;
  assign line_638_reset = reset;
  assign line_638_valid = superpage_hits_1 ^ line_638_valid_reg;
  assign line_639_clock = clock;
  assign line_639_reset = reset;
  assign line_639_valid = _T_989 ^ line_639_valid_reg;
  assign line_640_clock = clock;
  assign line_640_reset = reset;
  assign line_640_valid = superpage_entries_1_data_0[0] ^ line_640_valid_reg;
  assign line_641_clock = clock;
  assign line_641_reset = reset;
  assign line_641_valid = io_sfence_bits_rs1 ^ line_641_valid_reg;
  assign line_642_clock = clock;
  assign line_642_reset = reset;
  assign line_642_valid = io_sfence_bits_rs2 ^ line_642_valid_reg;
  assign line_643_clock = clock;
  assign line_643_reset = reset;
  assign line_643_valid = _T_1041 ^ line_643_valid_reg;
  assign line_644_clock = clock;
  assign line_644_reset = reset;
  assign line_644_valid = io_sfence_bits_rs2 ^ line_644_valid_reg;
  assign line_645_clock = clock;
  assign line_645_reset = reset;
  assign line_645_valid = io_sfence_bits_rs1 ^ line_645_valid_reg;
  assign line_646_clock = clock;
  assign line_646_reset = reset;
  assign line_646_valid = _hitsVec_T_56 ^ line_646_valid_reg;
  assign line_647_clock = clock;
  assign line_647_reset = reset;
  assign line_647_valid = _T_1087 ^ line_647_valid_reg;
  assign line_648_clock = clock;
  assign line_648_reset = reset;
  assign line_648_valid = special_entry_data_0[0] ^ line_648_valid_reg;
  assign line_649_clock = clock;
  assign line_649_reset = reset;
  assign line_649_valid = io_sfence_bits_rs1 ^ line_649_valid_reg;
  assign line_650_clock = clock;
  assign line_650_reset = reset;
  assign line_650_valid = io_sfence_bits_rs2 ^ line_650_valid_reg;
  assign line_651_clock = clock;
  assign line_651_reset = reset;
  assign line_651_valid = _T_1139 ^ line_651_valid_reg;
  assign line_652_clock = clock;
  assign line_652_reset = reset;
  assign line_652_valid = io_sfence_bits_rs2 ^ line_652_valid_reg;
  assign line_653_clock = clock;
  assign line_653_reset = reset;
  assign line_653_valid = _T_1433 ^ line_653_valid_reg;
  assign io_req_ready = state == 2'h0; // @[src/main/scala/rocket/TLB.scala 623:25]
  assign io_resp_miss = io_ptw_resp_valid | tlb_miss | multipleHits; // @[src/main/scala/rocket/TLB.scala 643:64]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[src/main/scala/rocket/TLB.scala 644:23]
  assign io_resp_pf_ld = bad_va & cmd_read | |_io_resp_pf_ld_T_1; // @[src/main/scala/rocket/TLB.scala 625:41]
  assign io_resp_pf_st = bad_va & cmd_write_perms | |_io_resp_pf_st_T_1; // @[src/main/scala/rocket/TLB.scala 626:48]
  assign io_resp_ae_ld = |_io_resp_ae_ld_T; // @[src/main/scala/rocket/TLB.scala 633:41]
  assign io_resp_ae_st = |_io_resp_ae_st_T; // @[src/main/scala/rocket/TLB.scala 634:41]
  assign io_resp_ma_ld = misaligned & cmd_read; // @[src/main/scala/rocket/TLB.scala 637:31]
  assign io_resp_ma_st = misaligned & cmd_write; // @[src/main/scala/rocket/TLB.scala 638:31]
  assign io_resp_cacheable = |_io_resp_cacheable_T; // @[src/main/scala/rocket/TLB.scala 640:41]
  assign io_ptw_req_valid = state == 2'h1; // @[src/main/scala/rocket/TLB.scala 652:29]
  assign io_ptw_req_bits_valid = 1'h1; // @[src/main/scala/rocket/TLB.scala 653:28]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[src/main/scala/rocket/TLB.scala 654:29]
  assign io_ptw_req_bits_bits_need_gpa = r_need_gpa; // @[src/main/scala/rocket/TLB.scala 657:33]
  assign mpu_ppn_barrier_clock = clock;
  assign mpu_ppn_barrier_reset = reset;
  assign mpu_ppn_barrier_io_x_ppn = special_entry_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign entries_barrier_clock = clock;
  assign entries_barrier_reset = reset;
  assign entries_barrier_io_x_ppn = _GEN_330[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_u = _GEN_330[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_ae_ptw = _GEN_330[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_ae_final = _GEN_330[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_pf = _GEN_330[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_gf = _GEN_330[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_sw = _GEN_330[14]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_sx = _GEN_330[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_sr = _GEN_330[12]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_pw = _GEN_330[8]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_pr = _GEN_330[6]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_ppp = _GEN_330[5]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_pal = _GEN_330[4]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_paa = _GEN_330[3]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_eff = _GEN_330[2]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_c = _GEN_330[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_clock = clock;
  assign entries_barrier_1_reset = reset;
  assign entries_barrier_1_io_x_ppn = _GEN_334[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_u = _GEN_334[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_ae_ptw = _GEN_334[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_ae_final = _GEN_334[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_pf = _GEN_334[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_gf = _GEN_334[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_sw = _GEN_334[14]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_sx = _GEN_334[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_sr = _GEN_334[12]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_pw = _GEN_334[8]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_pr = _GEN_334[6]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_ppp = _GEN_334[5]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_pal = _GEN_334[4]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_paa = _GEN_334[3]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_eff = _GEN_334[2]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_c = _GEN_334[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_clock = clock;
  assign entries_barrier_2_reset = reset;
  assign entries_barrier_2_io_x_ppn = superpage_entries_0_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_u = superpage_entries_0_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_ae_ptw = superpage_entries_0_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_ae_final = superpage_entries_0_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_pf = superpage_entries_0_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_gf = superpage_entries_0_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_sw = superpage_entries_0_data_0[14]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_sx = superpage_entries_0_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_sr = superpage_entries_0_data_0[12]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_pw = superpage_entries_0_data_0[8]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_pr = superpage_entries_0_data_0[6]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_ppp = superpage_entries_0_data_0[5]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_pal = superpage_entries_0_data_0[4]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_paa = superpage_entries_0_data_0[3]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_eff = superpage_entries_0_data_0[2]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_c = superpage_entries_0_data_0[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_clock = clock;
  assign entries_barrier_3_reset = reset;
  assign entries_barrier_3_io_x_ppn = superpage_entries_1_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_u = superpage_entries_1_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_ae_ptw = superpage_entries_1_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_ae_final = superpage_entries_1_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_pf = superpage_entries_1_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_gf = superpage_entries_1_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_sw = superpage_entries_1_data_0[14]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_sx = superpage_entries_1_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_sr = superpage_entries_1_data_0[12]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_pw = superpage_entries_1_data_0[8]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_pr = superpage_entries_1_data_0[6]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_ppp = superpage_entries_1_data_0[5]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_pal = superpage_entries_1_data_0[4]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_paa = superpage_entries_1_data_0[3]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_eff = superpage_entries_1_data_0[2]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_c = superpage_entries_1_data_0[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_clock = clock;
  assign entries_barrier_4_reset = reset;
  assign entries_barrier_4_io_x_ppn = special_entry_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_u = special_entry_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_ae_ptw = special_entry_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_ae_final = special_entry_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_pf = special_entry_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_gf = special_entry_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_sw = special_entry_data_0[14]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_sx = special_entry_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_sr = special_entry_data_0[12]; // @[src/main/scala/rocket/TLB.scala 160:77]
  always @(posedge clock) begin
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_0 <= _GEN_172;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_1 <= _GEN_173;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_2 <= _GEN_174;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_3 <= _GEN_175;
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_0 <= _GEN_366;
        end else begin
          sectored_entries_0_0_valid_0 <= _GEN_362;
        end
      end else begin
        sectored_entries_0_0_valid_0 <= _GEN_382;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_0 <= _GEN_228;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_1 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_1 <= _GEN_367;
        end else begin
          sectored_entries_0_0_valid_1 <= _GEN_363;
        end
      end else begin
        sectored_entries_0_0_valid_1 <= _GEN_383;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_1 <= _GEN_229;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_2 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_2 <= _GEN_368;
        end else begin
          sectored_entries_0_0_valid_2 <= _GEN_364;
        end
      end else begin
        sectored_entries_0_0_valid_2 <= _GEN_384;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_2 <= _GEN_230;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_3 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_3 <= _GEN_369;
        end else begin
          sectored_entries_0_0_valid_3 <= _GEN_365;
        end
      end else begin
        sectored_entries_0_0_valid_3 <= _GEN_385;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_3 <= _GEN_231;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_0 <= _GEN_199;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_1 <= _GEN_200;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_2 <= _GEN_201;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_3 <= _GEN_202;
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_0 <= _GEN_398;
        end else begin
          sectored_entries_0_1_valid_0 <= _GEN_394;
        end
      end else begin
        sectored_entries_0_1_valid_0 <= _GEN_414;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_0 <= _GEN_239;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_1 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_1 <= _GEN_399;
        end else begin
          sectored_entries_0_1_valid_1 <= _GEN_395;
        end
      end else begin
        sectored_entries_0_1_valid_1 <= _GEN_415;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_1 <= _GEN_240;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_2 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_2 <= _GEN_400;
        end else begin
          sectored_entries_0_1_valid_2 <= _GEN_396;
        end
      end else begin
        sectored_entries_0_1_valid_2 <= _GEN_416;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_2 <= _GEN_241;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_3 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_3 <= _GEN_401;
        end else begin
          sectored_entries_0_1_valid_3 <= _GEN_397;
        end
      end else begin
        sectored_entries_0_1_valid_3 <= _GEN_417;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_3 <= _GEN_242;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[src/main/scala/rocket/TLB.scala 203:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      superpage_entries_0_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_superpage_hits_T[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          superpage_entries_0_valid_0 <= _GEN_423;
        end else begin
          superpage_entries_0_valid_0 <= _GEN_422;
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_427;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        superpage_entries_0_valid_0 <= _GEN_221;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[src/main/scala/rocket/TLB.scala 203:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      superpage_entries_1_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_superpage_hits_T_14[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          superpage_entries_1_valid_0 <= _GEN_430;
        end else begin
          superpage_entries_1_valid_0 <= _GEN_429;
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_434;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        superpage_entries_1_valid_0 <= _GEN_226;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_level <= io_ptw_resp_bits_level; // @[src/main/scala/rocket/TLB.scala 203:16]
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      special_entry_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_hitsVec_T_42[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          special_entry_valid_0 <= _GEN_437;
        end else begin
          special_entry_valid_0 <= _GEN_436;
        end
      end else begin
        special_entry_valid_0 <= _GEN_441;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      special_entry_valid_0 <= _GEN_253;
    end
    if (reset) begin // @[src/main/scala/rocket/TLB.scala 341:22]
      state <= 2'h0; // @[src/main/scala/rocket/TLB.scala 341:22]
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 703:30]
      state <= 2'h0; // @[src/main/scala/rocket/TLB.scala 704:13]
    end else if (state == 2'h2 & io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 699:39]
      state <= 2'h3; // @[src/main/scala/rocket/TLB.scala 700:13]
    end else if (_invalidate_refill_T) begin // @[src/main/scala/rocket/TLB.scala 689:32]
      state <= _GEN_353;
    end else begin
      state <= _GEN_341;
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_refill_tag <= vpn; // @[src/main/scala/rocket/TLB.scala 671:20]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      if (&r_superpage_repl_addr_valids) begin // @[src/main/scala/rocket/TLB.scala 747:8]
        r_superpage_repl_addr <= state_reg_1;
      end else if (_r_superpage_repl_addr_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        r_superpage_repl_addr <= 1'h0;
      end else begin
        r_superpage_repl_addr <= 1'h1;
      end
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      if (&r_sectored_repl_addr_valids) begin // @[src/main/scala/rocket/TLB.scala 747:8]
        r_sectored_repl_addr <= state_vec_0;
      end else if (_r_sectored_repl_addr_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        r_sectored_repl_addr <= 1'h0;
      end else begin
        r_sectored_repl_addr <= 1'h1;
      end
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_sectored_hit_valid <= _T_10; // @[src/main/scala/rocket/TLB.scala 677:28]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_sectored_hit_bits <= state_vec_0_touch_way_sized; // @[src/main/scala/rocket/TLB.scala 678:27]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_need_gpa <= tlb_hit_if_not_gpa_miss; // @[src/main/scala/rocket/TLB.scala 672:18]
    end
    line_533_valid_reg <= 2'h0 == hitsVec_idx;
    line_534_valid_reg <= 2'h1 == hitsVec_idx;
    line_535_valid_reg <= 2'h2 == hitsVec_idx;
    line_536_valid_reg <= 2'h3 == hitsVec_idx;
    line_537_valid_reg <= 2'h0 == hitsVec_idx;
    line_538_valid_reg <= 2'h1 == hitsVec_idx;
    line_539_valid_reg <= 2'h2 == hitsVec_idx;
    line_540_valid_reg <= 2'h3 == hitsVec_idx;
    line_541_valid_reg <= io_ptw_resp_valid;
    line_542_valid_reg <= _T;
    line_543_valid_reg <= _T;
    line_544_valid_reg <= _T_2;
    line_545_valid_reg <= _T_3;
    line_546_valid_reg <= invalidate_refill;
    line_547_valid_reg <= r_superpage_repl_addr;
    line_548_valid_reg <= invalidate_refill;
    line_549_valid_reg <= _T_2;
    line_550_valid_reg <= _T_5;
    line_551_valid_reg <= _T_6;
    line_552_valid_reg <= 2'h0 == idx;
    line_553_valid_reg <= 2'h1 == idx;
    line_554_valid_reg <= 2'h2 == idx;
    line_555_valid_reg <= 2'h3 == idx;
    line_556_valid_reg <= 2'h0 == idx;
    line_557_valid_reg <= 2'h1 == idx;
    line_558_valid_reg <= 2'h2 == idx;
    line_559_valid_reg <= 2'h3 == idx;
    line_560_valid_reg <= invalidate_refill;
    if (r_sectored_hit_valid) begin // @[src/main/scala/rocket/TLB.scala 477:22]
      line_561_valid_reg <= r_sectored_hit_bits;
    end else begin
      line_561_valid_reg <= r_sectored_repl_addr;
    end
    line_562_valid_reg <= _T_6;
    line_563_valid_reg <= 2'h0 == idx;
    line_564_valid_reg <= 2'h1 == idx;
    line_565_valid_reg <= 2'h2 == idx;
    line_566_valid_reg <= 2'h3 == idx;
    line_567_valid_reg <= 2'h0 == idx;
    line_568_valid_reg <= 2'h1 == idx;
    line_569_valid_reg <= 2'h2 == idx;
    line_570_valid_reg <= 2'h3 == idx;
    line_571_valid_reg <= invalidate_refill;
    line_572_valid_reg <= 2'h0 == hitsVec_idx;
    line_573_valid_reg <= 2'h1 == hitsVec_idx;
    line_574_valid_reg <= 2'h2 == hitsVec_idx;
    line_575_valid_reg <= 2'h3 == hitsVec_idx;
    line_576_valid_reg <= 2'h0 == hitsVec_idx;
    line_577_valid_reg <= 2'h1 == hitsVec_idx;
    line_578_valid_reg <= 2'h2 == hitsVec_idx;
    line_579_valid_reg <= 2'h3 == hitsVec_idx;
    if (reset) begin // @[src/main/scala/util/Replacement.scala 374:17]
      state_vec_0 <= 1'h0; // @[src/main/scala/util/Replacement.scala 374:17]
    end else if (io_req_valid & vm_enabled) begin // @[src/main/scala/rocket/TLB.scala 609:37]
      if (_T_10) begin // @[src/main/scala/rocket/TLB.scala 611:28]
        state_vec_0 <= _state_vec_0_T_1; // @[src/main/scala/util/Replacement.scala 377:20]
      end
    end
    if (reset) begin // @[src/main/scala/util/Replacement.scala 168:72]
      state_reg_1 <= 1'h0; // @[src/main/scala/util/Replacement.scala 168:72]
    end else if (io_req_valid & vm_enabled) begin // @[src/main/scala/rocket/TLB.scala 609:37]
      if (_T_13) begin // @[src/main/scala/rocket/TLB.scala 612:31]
        state_reg_1 <= _state_reg_T_1; // @[src/main/scala/util/Replacement.scala 172:15]
      end
    end
    line_580_valid_reg <= _T_9;
    line_581_valid_reg <= _T_10;
    line_582_valid_reg <= _T_13;
    line_583_valid_reg <= _T_17;
    line_584_valid_reg <= _T_19;
    line_585_valid_reg <= _invalidate_refill_T;
    line_586_valid_reg <= io_sfence_valid;
    line_587_valid_reg <= io_ptw_req_ready;
    line_588_valid_reg <= _T_22;
    line_589_valid_reg <= io_ptw_resp_valid;
    line_590_valid_reg <= io_sfence_valid;
    line_591_valid_reg <= _T_28;
    line_592_valid_reg <= _T_29;
    line_593_valid_reg <= io_sfence_bits_rs1;
    line_594_valid_reg <= _sector_hits_T_5;
    line_595_valid_reg <= _GEN_0;
    line_596_valid_reg <= _GEN_1;
    line_597_valid_reg <= _GEN_2;
    line_598_valid_reg <= _GEN_3;
    line_599_valid_reg <= _T_147;
    line_600_valid_reg <= sectored_entries_0_0_data_0[0];
    line_601_valid_reg <= sectored_entries_0_0_data_1[0];
    line_602_valid_reg <= sectored_entries_0_0_data_2[0];
    line_603_valid_reg <= sectored_entries_0_0_data_3[0];
    line_604_valid_reg <= io_sfence_bits_rs1;
    line_605_valid_reg <= io_sfence_bits_rs2;
    line_606_valid_reg <= _T_343;
    line_607_valid_reg <= _T_346;
    line_608_valid_reg <= _T_349;
    line_609_valid_reg <= _T_352;
    line_610_valid_reg <= io_sfence_bits_rs2;
    line_611_valid_reg <= io_sfence_bits_rs1;
    line_612_valid_reg <= _sector_hits_T_13;
    line_613_valid_reg <= _GEN_0;
    line_614_valid_reg <= _GEN_1;
    line_615_valid_reg <= _GEN_2;
    line_616_valid_reg <= _GEN_3;
    line_617_valid_reg <= _T_568;
    line_618_valid_reg <= sectored_entries_0_1_data_0[0];
    line_619_valid_reg <= sectored_entries_0_1_data_1[0];
    line_620_valid_reg <= sectored_entries_0_1_data_2[0];
    line_621_valid_reg <= sectored_entries_0_1_data_3[0];
    line_622_valid_reg <= io_sfence_bits_rs1;
    line_623_valid_reg <= io_sfence_bits_rs2;
    line_624_valid_reg <= _T_764;
    line_625_valid_reg <= _T_767;
    line_626_valid_reg <= _T_770;
    line_627_valid_reg <= _T_773;
    line_628_valid_reg <= io_sfence_bits_rs2;
    line_629_valid_reg <= io_sfence_bits_rs1;
    line_630_valid_reg <= superpage_hits_0;
    line_631_valid_reg <= _T_891;
    line_632_valid_reg <= superpage_entries_0_data_0[0];
    line_633_valid_reg <= io_sfence_bits_rs1;
    line_634_valid_reg <= io_sfence_bits_rs2;
    line_635_valid_reg <= _T_943;
    line_636_valid_reg <= io_sfence_bits_rs2;
    line_637_valid_reg <= io_sfence_bits_rs1;
    line_638_valid_reg <= superpage_hits_1;
    line_639_valid_reg <= _T_989;
    line_640_valid_reg <= superpage_entries_1_data_0[0];
    line_641_valid_reg <= io_sfence_bits_rs1;
    line_642_valid_reg <= io_sfence_bits_rs2;
    line_643_valid_reg <= _T_1041;
    line_644_valid_reg <= io_sfence_bits_rs2;
    line_645_valid_reg <= io_sfence_bits_rs1;
    line_646_valid_reg <= _hitsVec_T_56;
    line_647_valid_reg <= _T_1087;
    line_648_valid_reg <= special_entry_data_0[0];
    line_649_valid_reg <= io_sfence_bits_rs1;
    line_650_valid_reg <= io_sfence_bits_rs2;
    line_651_valid_reg <= _T_1139;
    line_652_valid_reg <= io_sfence_bits_rs2;
    line_653_valid_reg <= _T_1433;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~reset & ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TLB.scala:709 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"
            ); // @[src/main/scala/rocket/TLB.scala 709:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_0_tag_vpn = _RAND_0[26:0];
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_0_data_0 = _RAND_1[41:0];
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_0_data_1 = _RAND_2[41:0];
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_0_data_2 = _RAND_3[41:0];
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_0_data_3 = _RAND_4[41:0];
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_0_1_tag_vpn = _RAND_9[26:0];
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_0_1_data_0 = _RAND_10[41:0];
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_0_1_data_1 = _RAND_11[41:0];
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_0_1_data_2 = _RAND_12[41:0];
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_0_1_data_3 = _RAND_13[41:0];
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_0_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_0_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_0_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_0_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  superpage_entries_0_tag_vpn = _RAND_19[26:0];
  _RAND_20 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_20[41:0];
  _RAND_21 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  superpage_entries_1_tag_vpn = _RAND_23[26:0];
  _RAND_24 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_24[41:0];
  _RAND_25 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  special_entry_level = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  special_entry_tag_vpn = _RAND_27[26:0];
  _RAND_28 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_28[41:0];
  _RAND_29 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  r_refill_tag = _RAND_31[26:0];
  _RAND_32 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_sectored_hit_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_sectored_hit_bits = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_need_gpa = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_533_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_534_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_535_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_536_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_537_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_538_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_539_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_540_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_541_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_542_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_543_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_544_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_545_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_546_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_547_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_548_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_549_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_550_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_551_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_552_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_553_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_554_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_555_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_556_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_557_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_558_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_559_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_560_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_561_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_562_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_563_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_564_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_565_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_566_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_567_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_568_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_569_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_570_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_571_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_572_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_573_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_574_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_575_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_576_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_577_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_578_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_579_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  state_vec_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  state_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_580_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_581_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_582_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_583_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_584_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_585_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_586_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_587_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_588_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_589_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_590_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_591_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_592_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_593_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_594_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_595_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_596_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_597_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_598_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_599_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_600_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_601_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_602_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_603_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_604_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_605_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_606_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_607_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_608_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_609_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_610_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_611_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_612_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_613_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_614_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_615_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_616_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_617_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_618_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_619_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_620_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_621_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_622_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_623_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_624_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_625_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_626_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_627_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_628_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_629_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_630_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_631_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_632_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_633_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_634_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_635_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_636_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_637_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_638_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_639_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_640_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_641_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_642_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_643_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_644_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_645_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_646_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_647_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_648_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_649_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_650_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_651_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_652_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_653_valid_reg = _RAND_159[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (io_sfence_valid & ~reset) begin
      assert(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn); // @[src/main/scala/rocket/TLB.scala 709:13]
    end
  end
endmodule
module OptimizationBarrier_6(
  input   clock,
  input   reset
);
endmodule
module PMPChecker_1(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_7(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_8(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_9(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_10(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_11(
  input   clock,
  input   reset
);
endmodule
module DCacheModuleImpl_Anon(
  input         clock,
  input         reset,
  input  [39:0] io_req_bits_vaddr // @[src/main/scala/rocket/TLB.scala 309:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  mpu_ppn_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  mpu_ppn_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire  pmp_clock; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  pmp_reset; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  entries_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_reset; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_reset; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_reset; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [26:0] vpn = io_req_bits_vaddr[38:12]; // @[src/main/scala/rocket/TLB.scala 324:30]
  wire  _sector_hits_T_5 = vpn[26:2] == 25'h0; // @[src/main/scala/rocket/TLB.scala 164:86]
  wire [1:0] hitsVec_idx = vpn[1:0]; // @[src/main/scala/util/package.scala 155:13]
  wire  _GEN_0 = 2'h0 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_654_clock;
  wire  line_654_reset;
  wire  line_654_valid;
  reg  line_654_valid_reg;
  wire  _GEN_1 = 2'h1 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_655_clock;
  wire  line_655_reset;
  wire  line_655_valid;
  reg  line_655_valid_reg;
  wire  _GEN_2 = 2'h2 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_656_clock;
  wire  line_656_reset;
  wire  line_656_valid;
  reg  line_656_valid_reg;
  wire  _GEN_3 = 2'h3 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_657_clock;
  wire  line_657_reset;
  wire  line_657_valid;
  reg  line_657_valid_reg;
  wire  line_658_clock;
  wire  line_658_reset;
  wire  line_658_valid;
  reg  line_658_valid_reg;
  wire  line_659_clock;
  wire  line_659_reset;
  wire  line_659_valid;
  reg  line_659_valid_reg;
  wire  line_660_clock;
  wire  line_660_reset;
  wire  line_660_valid;
  reg  line_660_valid_reg;
  wire  line_661_clock;
  wire  line_661_reset;
  wire  line_661_valid;
  reg  line_661_valid_reg;
  wire  line_662_clock;
  wire  line_662_reset;
  wire  line_662_valid;
  reg  line_662_valid_reg;
  wire  line_663_clock;
  wire  line_663_reset;
  wire  line_663_valid;
  reg  line_663_valid_reg;
  wire  line_664_clock;
  wire  line_664_reset;
  wire  line_664_valid;
  reg  line_664_valid_reg;
  wire  line_665_clock;
  wire  line_665_reset;
  wire  line_665_valid;
  reg  line_665_valid_reg;
  wire  line_666_clock;
  wire  line_666_reset;
  wire  line_666_valid;
  reg  line_666_valid_reg;
  wire  line_667_clock;
  wire  line_667_reset;
  wire  line_667_valid;
  reg  line_667_valid_reg;
  wire  line_668_clock;
  wire  line_668_reset;
  wire  line_668_valid;
  reg  line_668_valid_reg;
  wire  line_669_clock;
  wire  line_669_reset;
  wire  line_669_valid;
  reg  line_669_valid_reg;
  wire  _T_28 = ~reset; // @[src/main/scala/rocket/TLB.scala 709:13]
  wire  line_670_clock;
  wire  line_670_reset;
  wire  line_670_valid;
  reg  line_670_valid_reg;
  wire  line_671_clock;
  wire  line_671_reset;
  wire  line_671_valid;
  reg  line_671_valid_reg;
  wire  line_672_clock;
  wire  line_672_reset;
  wire  line_672_valid;
  reg  line_672_valid_reg;
  wire  line_673_clock;
  wire  line_673_reset;
  wire  line_673_valid;
  reg  line_673_valid_reg;
  wire  line_674_clock;
  wire  line_674_reset;
  wire  line_674_valid;
  reg  line_674_valid_reg;
  wire  line_675_clock;
  wire  line_675_reset;
  wire  line_675_valid;
  reg  line_675_valid_reg;
  wire  _T_147 = vpn[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_676_clock;
  wire  line_676_reset;
  wire  line_676_valid;
  reg  line_676_valid_reg;
  wire  line_677_clock;
  wire  line_677_reset;
  wire  line_677_valid;
  reg  line_677_valid_reg;
  wire  line_678_clock;
  wire  line_678_reset;
  wire  line_678_valid;
  reg  line_678_valid_reg;
  wire  line_679_clock;
  wire  line_679_reset;
  wire  line_679_valid;
  reg  line_679_valid_reg;
  wire  line_680_clock;
  wire  line_680_reset;
  wire  line_680_valid;
  reg  line_680_valid_reg;
  wire  line_681_clock;
  wire  line_681_reset;
  wire  line_681_valid;
  reg  line_681_valid_reg;
  wire  line_682_clock;
  wire  line_682_reset;
  wire  line_682_valid;
  reg  line_682_valid_reg;
  wire  line_683_clock;
  wire  line_683_reset;
  wire  line_683_valid;
  reg  line_683_valid_reg;
  wire  line_684_clock;
  wire  line_684_reset;
  wire  line_684_valid;
  reg  line_684_valid_reg;
  wire  line_685_clock;
  wire  line_685_reset;
  wire  line_685_valid;
  reg  line_685_valid_reg;
  wire  line_686_clock;
  wire  line_686_reset;
  wire  line_686_valid;
  reg  line_686_valid_reg;
  OptimizationBarrier_6 mpu_ppn_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(mpu_ppn_barrier_clock),
    .reset(mpu_ppn_barrier_reset)
  );
  PMPChecker_1 pmp ( // @[src/main/scala/rocket/TLB.scala 405:19]
    .clock(pmp_clock),
    .reset(pmp_reset)
  );
  OptimizationBarrier_7 entries_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_clock),
    .reset(entries_barrier_reset)
  );
  OptimizationBarrier_8 entries_barrier_1 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_1_clock),
    .reset(entries_barrier_1_reset)
  );
  OptimizationBarrier_9 entries_barrier_2 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_2_clock),
    .reset(entries_barrier_2_reset)
  );
  OptimizationBarrier_10 entries_barrier_3 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_3_clock),
    .reset(entries_barrier_3_reset)
  );
  OptimizationBarrier_11 entries_barrier_4 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_4_clock),
    .reset(entries_barrier_4_reset)
  );
  GEN_w1_line #(.COVER_INDEX(654)) line_654 (
    .clock(line_654_clock),
    .reset(line_654_reset),
    .valid(line_654_valid)
  );
  GEN_w1_line #(.COVER_INDEX(655)) line_655 (
    .clock(line_655_clock),
    .reset(line_655_reset),
    .valid(line_655_valid)
  );
  GEN_w1_line #(.COVER_INDEX(656)) line_656 (
    .clock(line_656_clock),
    .reset(line_656_reset),
    .valid(line_656_valid)
  );
  GEN_w1_line #(.COVER_INDEX(657)) line_657 (
    .clock(line_657_clock),
    .reset(line_657_reset),
    .valid(line_657_valid)
  );
  GEN_w1_line #(.COVER_INDEX(658)) line_658 (
    .clock(line_658_clock),
    .reset(line_658_reset),
    .valid(line_658_valid)
  );
  GEN_w1_line #(.COVER_INDEX(659)) line_659 (
    .clock(line_659_clock),
    .reset(line_659_reset),
    .valid(line_659_valid)
  );
  GEN_w1_line #(.COVER_INDEX(660)) line_660 (
    .clock(line_660_clock),
    .reset(line_660_reset),
    .valid(line_660_valid)
  );
  GEN_w1_line #(.COVER_INDEX(661)) line_661 (
    .clock(line_661_clock),
    .reset(line_661_reset),
    .valid(line_661_valid)
  );
  GEN_w1_line #(.COVER_INDEX(662)) line_662 (
    .clock(line_662_clock),
    .reset(line_662_reset),
    .valid(line_662_valid)
  );
  GEN_w1_line #(.COVER_INDEX(663)) line_663 (
    .clock(line_663_clock),
    .reset(line_663_reset),
    .valid(line_663_valid)
  );
  GEN_w1_line #(.COVER_INDEX(664)) line_664 (
    .clock(line_664_clock),
    .reset(line_664_reset),
    .valid(line_664_valid)
  );
  GEN_w1_line #(.COVER_INDEX(665)) line_665 (
    .clock(line_665_clock),
    .reset(line_665_reset),
    .valid(line_665_valid)
  );
  GEN_w1_line #(.COVER_INDEX(666)) line_666 (
    .clock(line_666_clock),
    .reset(line_666_reset),
    .valid(line_666_valid)
  );
  GEN_w1_line #(.COVER_INDEX(667)) line_667 (
    .clock(line_667_clock),
    .reset(line_667_reset),
    .valid(line_667_valid)
  );
  GEN_w1_line #(.COVER_INDEX(668)) line_668 (
    .clock(line_668_clock),
    .reset(line_668_reset),
    .valid(line_668_valid)
  );
  GEN_w1_line #(.COVER_INDEX(669)) line_669 (
    .clock(line_669_clock),
    .reset(line_669_reset),
    .valid(line_669_valid)
  );
  GEN_w1_line #(.COVER_INDEX(670)) line_670 (
    .clock(line_670_clock),
    .reset(line_670_reset),
    .valid(line_670_valid)
  );
  GEN_w1_line #(.COVER_INDEX(671)) line_671 (
    .clock(line_671_clock),
    .reset(line_671_reset),
    .valid(line_671_valid)
  );
  GEN_w1_line #(.COVER_INDEX(672)) line_672 (
    .clock(line_672_clock),
    .reset(line_672_reset),
    .valid(line_672_valid)
  );
  GEN_w1_line #(.COVER_INDEX(673)) line_673 (
    .clock(line_673_clock),
    .reset(line_673_reset),
    .valid(line_673_valid)
  );
  GEN_w1_line #(.COVER_INDEX(674)) line_674 (
    .clock(line_674_clock),
    .reset(line_674_reset),
    .valid(line_674_valid)
  );
  GEN_w1_line #(.COVER_INDEX(675)) line_675 (
    .clock(line_675_clock),
    .reset(line_675_reset),
    .valid(line_675_valid)
  );
  GEN_w1_line #(.COVER_INDEX(676)) line_676 (
    .clock(line_676_clock),
    .reset(line_676_reset),
    .valid(line_676_valid)
  );
  GEN_w1_line #(.COVER_INDEX(677)) line_677 (
    .clock(line_677_clock),
    .reset(line_677_reset),
    .valid(line_677_valid)
  );
  GEN_w1_line #(.COVER_INDEX(678)) line_678 (
    .clock(line_678_clock),
    .reset(line_678_reset),
    .valid(line_678_valid)
  );
  GEN_w1_line #(.COVER_INDEX(679)) line_679 (
    .clock(line_679_clock),
    .reset(line_679_reset),
    .valid(line_679_valid)
  );
  GEN_w1_line #(.COVER_INDEX(680)) line_680 (
    .clock(line_680_clock),
    .reset(line_680_reset),
    .valid(line_680_valid)
  );
  GEN_w1_line #(.COVER_INDEX(681)) line_681 (
    .clock(line_681_clock),
    .reset(line_681_reset),
    .valid(line_681_valid)
  );
  GEN_w1_line #(.COVER_INDEX(682)) line_682 (
    .clock(line_682_clock),
    .reset(line_682_reset),
    .valid(line_682_valid)
  );
  GEN_w1_line #(.COVER_INDEX(683)) line_683 (
    .clock(line_683_clock),
    .reset(line_683_reset),
    .valid(line_683_valid)
  );
  GEN_w1_line #(.COVER_INDEX(684)) line_684 (
    .clock(line_684_clock),
    .reset(line_684_reset),
    .valid(line_684_valid)
  );
  GEN_w1_line #(.COVER_INDEX(685)) line_685 (
    .clock(line_685_clock),
    .reset(line_685_reset),
    .valid(line_685_valid)
  );
  GEN_w1_line #(.COVER_INDEX(686)) line_686 (
    .clock(line_686_clock),
    .reset(line_686_reset),
    .valid(line_686_valid)
  );
  assign line_654_clock = clock;
  assign line_654_reset = reset;
  assign line_654_valid = 2'h0 == hitsVec_idx ^ line_654_valid_reg;
  assign line_655_clock = clock;
  assign line_655_reset = reset;
  assign line_655_valid = 2'h1 == hitsVec_idx ^ line_655_valid_reg;
  assign line_656_clock = clock;
  assign line_656_reset = reset;
  assign line_656_valid = 2'h2 == hitsVec_idx ^ line_656_valid_reg;
  assign line_657_clock = clock;
  assign line_657_reset = reset;
  assign line_657_valid = 2'h3 == hitsVec_idx ^ line_657_valid_reg;
  assign line_658_clock = clock;
  assign line_658_reset = reset;
  assign line_658_valid = 2'h0 == hitsVec_idx ^ line_658_valid_reg;
  assign line_659_clock = clock;
  assign line_659_reset = reset;
  assign line_659_valid = 2'h1 == hitsVec_idx ^ line_659_valid_reg;
  assign line_660_clock = clock;
  assign line_660_reset = reset;
  assign line_660_valid = 2'h2 == hitsVec_idx ^ line_660_valid_reg;
  assign line_661_clock = clock;
  assign line_661_reset = reset;
  assign line_661_valid = 2'h3 == hitsVec_idx ^ line_661_valid_reg;
  assign line_662_clock = clock;
  assign line_662_reset = reset;
  assign line_662_valid = 2'h0 == hitsVec_idx ^ line_662_valid_reg;
  assign line_663_clock = clock;
  assign line_663_reset = reset;
  assign line_663_valid = 2'h1 == hitsVec_idx ^ line_663_valid_reg;
  assign line_664_clock = clock;
  assign line_664_reset = reset;
  assign line_664_valid = 2'h2 == hitsVec_idx ^ line_664_valid_reg;
  assign line_665_clock = clock;
  assign line_665_reset = reset;
  assign line_665_valid = 2'h3 == hitsVec_idx ^ line_665_valid_reg;
  assign line_666_clock = clock;
  assign line_666_reset = reset;
  assign line_666_valid = 2'h0 == hitsVec_idx ^ line_666_valid_reg;
  assign line_667_clock = clock;
  assign line_667_reset = reset;
  assign line_667_valid = 2'h1 == hitsVec_idx ^ line_667_valid_reg;
  assign line_668_clock = clock;
  assign line_668_reset = reset;
  assign line_668_valid = 2'h2 == hitsVec_idx ^ line_668_valid_reg;
  assign line_669_clock = clock;
  assign line_669_reset = reset;
  assign line_669_valid = 2'h3 == hitsVec_idx ^ line_669_valid_reg;
  assign line_670_clock = clock;
  assign line_670_reset = reset;
  assign line_670_valid = _T_28 ^ line_670_valid_reg;
  assign line_671_clock = clock;
  assign line_671_reset = reset;
  assign line_671_valid = _sector_hits_T_5 ^ line_671_valid_reg;
  assign line_672_clock = clock;
  assign line_672_reset = reset;
  assign line_672_valid = _GEN_0 ^ line_672_valid_reg;
  assign line_673_clock = clock;
  assign line_673_reset = reset;
  assign line_673_valid = _GEN_1 ^ line_673_valid_reg;
  assign line_674_clock = clock;
  assign line_674_reset = reset;
  assign line_674_valid = _GEN_2 ^ line_674_valid_reg;
  assign line_675_clock = clock;
  assign line_675_reset = reset;
  assign line_675_valid = _GEN_3 ^ line_675_valid_reg;
  assign line_676_clock = clock;
  assign line_676_reset = reset;
  assign line_676_valid = _T_147 ^ line_676_valid_reg;
  assign line_677_clock = clock;
  assign line_677_reset = reset;
  assign line_677_valid = _sector_hits_T_5 ^ line_677_valid_reg;
  assign line_678_clock = clock;
  assign line_678_reset = reset;
  assign line_678_valid = _GEN_0 ^ line_678_valid_reg;
  assign line_679_clock = clock;
  assign line_679_reset = reset;
  assign line_679_valid = _GEN_1 ^ line_679_valid_reg;
  assign line_680_clock = clock;
  assign line_680_reset = reset;
  assign line_680_valid = _GEN_2 ^ line_680_valid_reg;
  assign line_681_clock = clock;
  assign line_681_reset = reset;
  assign line_681_valid = _GEN_3 ^ line_681_valid_reg;
  assign line_682_clock = clock;
  assign line_682_reset = reset;
  assign line_682_valid = _T_147 ^ line_682_valid_reg;
  assign line_683_clock = clock;
  assign line_683_reset = reset;
  assign line_683_valid = _T_147 ^ line_683_valid_reg;
  assign line_684_clock = clock;
  assign line_684_reset = reset;
  assign line_684_valid = _T_147 ^ line_684_valid_reg;
  assign line_685_clock = clock;
  assign line_685_reset = reset;
  assign line_685_valid = _T_147 ^ line_685_valid_reg;
  assign line_686_clock = clock;
  assign line_686_reset = reset;
  assign line_686_valid = reset ^ line_686_valid_reg;
  assign mpu_ppn_barrier_clock = clock;
  assign mpu_ppn_barrier_reset = reset;
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign entries_barrier_clock = clock;
  assign entries_barrier_reset = reset;
  assign entries_barrier_1_clock = clock;
  assign entries_barrier_1_reset = reset;
  assign entries_barrier_2_clock = clock;
  assign entries_barrier_2_reset = reset;
  assign entries_barrier_3_clock = clock;
  assign entries_barrier_3_reset = reset;
  assign entries_barrier_4_clock = clock;
  assign entries_barrier_4_reset = reset;
  always @(posedge clock) begin
    line_654_valid_reg <= 2'h0 == hitsVec_idx;
    line_655_valid_reg <= 2'h1 == hitsVec_idx;
    line_656_valid_reg <= 2'h2 == hitsVec_idx;
    line_657_valid_reg <= 2'h3 == hitsVec_idx;
    line_658_valid_reg <= 2'h0 == hitsVec_idx;
    line_659_valid_reg <= 2'h1 == hitsVec_idx;
    line_660_valid_reg <= 2'h2 == hitsVec_idx;
    line_661_valid_reg <= 2'h3 == hitsVec_idx;
    line_662_valid_reg <= 2'h0 == hitsVec_idx;
    line_663_valid_reg <= 2'h1 == hitsVec_idx;
    line_664_valid_reg <= 2'h2 == hitsVec_idx;
    line_665_valid_reg <= 2'h3 == hitsVec_idx;
    line_666_valid_reg <= 2'h0 == hitsVec_idx;
    line_667_valid_reg <= 2'h1 == hitsVec_idx;
    line_668_valid_reg <= 2'h2 == hitsVec_idx;
    line_669_valid_reg <= 2'h3 == hitsVec_idx;
    line_670_valid_reg <= _T_28;
    line_671_valid_reg <= _sector_hits_T_5;
    line_672_valid_reg <= _GEN_0;
    line_673_valid_reg <= _GEN_1;
    line_674_valid_reg <= _GEN_2;
    line_675_valid_reg <= _GEN_3;
    line_676_valid_reg <= _T_147;
    line_677_valid_reg <= _sector_hits_T_5;
    line_678_valid_reg <= _GEN_0;
    line_679_valid_reg <= _GEN_1;
    line_680_valid_reg <= _GEN_2;
    line_681_valid_reg <= _GEN_3;
    line_682_valid_reg <= _T_147;
    line_683_valid_reg <= _T_147;
    line_684_valid_reg <= _T_147;
    line_685_valid_reg <= _T_147;
    line_686_valid_reg <= reset;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_654_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_655_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_656_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_657_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_658_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_659_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_660_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_661_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_662_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_663_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_664_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_665_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_666_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_667_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_668_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_669_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_670_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_671_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_672_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_673_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_674_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  line_675_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_676_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  line_677_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_678_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_679_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_680_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_681_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_682_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_683_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_684_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_685_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_686_valid_reg = _RAND_32[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  input   io_increment // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  line_687_clock;
  wire  line_687_reset;
  wire  line_687_valid;
  reg  line_687_valid_reg;
  GEN_w1_line #(.COVER_INDEX(687)) line_687 (
    .clock(line_687_clock),
    .reset(line_687_reset),
    .valid(line_687_valid)
  );
  assign line_687_clock = clock;
  assign line_687_reset = reset;
  assign line_687_valid = io_increment ^ line_687_valid_reg;
  always @(posedge clock) begin
    line_687_valid_reg <= io_increment;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_687_valid_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheModuleImpl_Anon_1(
  input         clock,
  input         reset,
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_2_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [27:0] io_in_2_bits_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_3_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_3_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_3_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [27:0] io_in_3_bits_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_4_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_4_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_4_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_4_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [27:0] io_in_4_bits_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_5_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_5_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_5_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_5_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_6_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_6_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_6_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_6_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [27:0] io_in_6_bits_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_7_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_7_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [39:0] io_in_7_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_7_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [27:0] io_in_7_bits_data, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_write, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [39:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_idx, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [27:0] io_out_bits_data // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  line_688_clock;
  wire  line_688_reset;
  wire  line_688_valid;
  reg  line_688_valid_reg;
  wire [39:0] _GEN_9 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  wire  _GEN_10 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  wire [27:0] _GEN_12 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  wire  line_689_clock;
  wire  line_689_reset;
  wire  line_689_valid;
  reg  line_689_valid_reg;
  wire [39:0] _GEN_21 = io_in_4_valid ? io_in_4_bits_addr : _GEN_9; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  _GEN_22 = io_in_4_valid ? io_in_4_bits_idx : _GEN_10; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire [27:0] _GEN_24 = io_in_4_valid ? io_in_4_bits_data : _GEN_12; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  line_690_clock;
  wire  line_690_reset;
  wire  line_690_valid;
  reg  line_690_valid_reg;
  wire [39:0] _GEN_27 = io_in_3_valid ? io_in_3_bits_addr : _GEN_21; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  _GEN_28 = io_in_3_valid ? io_in_3_bits_idx : _GEN_22; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire [27:0] _GEN_30 = io_in_3_valid ? io_in_3_bits_data : _GEN_24; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  line_691_clock;
  wire  line_691_reset;
  wire  line_691_valid;
  reg  line_691_valid_reg;
  wire [39:0] _GEN_33 = io_in_2_valid ? io_in_2_bits_addr : _GEN_27; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  _GEN_34 = io_in_2_valid ? io_in_2_bits_idx : _GEN_28; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire [27:0] _GEN_36 = io_in_2_valid ? io_in_2_bits_data : _GEN_30; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  line_692_clock;
  wire  line_692_reset;
  wire  line_692_valid;
  reg  line_692_valid_reg;
  wire  grant_7 = ~(io_in_0_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid | io_in_6_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  GEN_w1_line #(.COVER_INDEX(688)) line_688 (
    .clock(line_688_clock),
    .reset(line_688_reset),
    .valid(line_688_valid)
  );
  GEN_w1_line #(.COVER_INDEX(689)) line_689 (
    .clock(line_689_clock),
    .reset(line_689_reset),
    .valid(line_689_valid)
  );
  GEN_w1_line #(.COVER_INDEX(690)) line_690 (
    .clock(line_690_clock),
    .reset(line_690_reset),
    .valid(line_690_valid)
  );
  GEN_w1_line #(.COVER_INDEX(691)) line_691 (
    .clock(line_691_clock),
    .reset(line_691_reset),
    .valid(line_691_valid)
  );
  GEN_w1_line #(.COVER_INDEX(692)) line_692 (
    .clock(line_692_clock),
    .reset(line_692_reset),
    .valid(line_692_valid)
  );
  assign line_688_clock = clock;
  assign line_688_reset = reset;
  assign line_688_valid = io_in_6_valid ^ line_688_valid_reg;
  assign line_689_clock = clock;
  assign line_689_reset = reset;
  assign line_689_valid = io_in_4_valid ^ line_689_valid_reg;
  assign line_690_clock = clock;
  assign line_690_reset = reset;
  assign line_690_valid = io_in_3_valid ^ line_690_valid_reg;
  assign line_691_clock = clock;
  assign line_691_reset = reset;
  assign line_691_valid = io_in_2_valid ^ line_691_valid_reg;
  assign line_692_clock = clock;
  assign line_692_reset = reset;
  assign line_692_valid = io_in_0_valid ^ line_692_valid_reg;
  assign io_in_4_ready = ~(io_in_0_valid | io_in_2_valid | io_in_3_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_5_ready = ~(io_in_0_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_6_ready = ~(io_in_0_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_7_ready = ~(io_in_0_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid | io_in_6_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_7 | io_in_7_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_write = io_in_0_valid | (io_in_2_valid | (io_in_3_valid | io_in_4_valid)); // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_33; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_idx = io_in_0_valid ? io_in_0_bits_idx : _GEN_34; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_data = io_in_0_valid ? 28'h0 : _GEN_36; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  always @(posedge clock) begin
    line_688_valid_reg <= io_in_6_valid;
    line_689_valid_reg <= io_in_4_valid;
    line_690_valid_reg <= io_in_3_valid;
    line_691_valid_reg <= io_in_2_valid;
    line_692_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_688_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_689_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_690_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_691_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_692_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheDataArray(
  input         clock,
  input         reset,
  input         io_req_valid, // @[src/main/scala/rocket/DCache.scala 43:14]
  input  [5:0]  io_req_bits_addr, // @[src/main/scala/rocket/DCache.scala 43:14]
  input         io_req_bits_write, // @[src/main/scala/rocket/DCache.scala 43:14]
  input  [63:0] io_req_bits_wdata, // @[src/main/scala/rocket/DCache.scala 43:14]
  input  [7:0]  io_req_bits_eccMask, // @[src/main/scala/rocket/DCache.scala 43:14]
  output [63:0] io_resp_0 // @[src/main/scala/rocket/DCache.scala 43:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_arrays_0_0 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_0_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_0_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_0_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_0_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_0_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_0_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_1 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_1_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_1_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_1_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_1_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_1_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_1_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_1_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_1_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_1_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_2 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_2_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_2_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_2_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_2_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_2_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_2_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_2_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_2_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_2_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_3 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_3_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_3_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_3_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_3_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_3_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_3_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_3_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_3_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_3_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_4 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_4_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_4_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_4_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_4_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_4_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_4_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_4_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_4_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_4_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_5 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_5_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_5_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_5_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_5_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_5_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_5_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_5_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_5_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_5_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_6 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_6_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_6_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_6_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_6_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_6_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_6_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_6_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_6_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_6_rdata_data_addr_pipe_0;
  reg [7:0] data_arrays_0_7 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_7_rdata_data_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_7_rdata_data_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_7_rdata_data_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [7:0] data_arrays_0_7_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_7_rdata_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_7_rdata_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_7_rdata_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_7_rdata_data_en_pipe_0;
  reg [2:0] data_arrays_0_7_rdata_data_addr_pipe_0;
  wire  eccMask_0 = io_req_bits_eccMask[0]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_1 = io_req_bits_eccMask[1]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_2 = io_req_bits_eccMask[2]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_3 = io_req_bits_eccMask[3]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_4 = io_req_bits_eccMask[4]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_5 = io_req_bits_eccMask[5]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_6 = io_req_bits_eccMask[6]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  eccMask_7 = io_req_bits_eccMask[7]; // @[src/main/scala/rocket/DCache.scala 49:82]
  wire  _rdata_T = io_req_valid & io_req_bits_write; // @[src/main/scala/rocket/DCache.scala 65:17]
  wire  line_693_clock;
  wire  line_693_reset;
  wire  line_693_valid;
  reg  line_693_valid_reg;
  wire  line_694_clock;
  wire  line_694_reset;
  wire  line_694_valid;
  reg  line_694_valid_reg;
  wire  line_695_clock;
  wire  line_695_reset;
  wire  line_695_valid;
  reg  line_695_valid_reg;
  wire  line_696_clock;
  wire  line_696_reset;
  wire  line_696_valid;
  reg  line_696_valid_reg;
  wire  line_697_clock;
  wire  line_697_reset;
  wire  line_697_valid;
  reg  line_697_valid_reg;
  wire  line_698_clock;
  wire  line_698_reset;
  wire  line_698_valid;
  reg  line_698_valid_reg;
  wire  line_699_clock;
  wire  line_699_reset;
  wire  line_699_valid;
  reg  line_699_valid_reg;
  wire  line_700_clock;
  wire  line_700_reset;
  wire  line_700_valid;
  reg  line_700_valid_reg;
  wire  line_701_clock;
  wire  line_701_reset;
  wire  line_701_valid;
  reg  line_701_valid_reg;
  wire  _rdata_data_T = ~io_req_bits_write; // @[src/main/scala/rocket/DCache.scala 70:42]
  wire  _rdata_data_T_1 = io_req_valid & ~io_req_bits_write; // @[src/main/scala/rocket/DCache.scala 70:39]
  wire  line_702_clock;
  wire  line_702_reset;
  wire  line_702_valid;
  reg  line_702_valid_reg;
  wire [31:0] rdata_lo = {data_arrays_0_3_rdata_data_data,data_arrays_0_2_rdata_data_data,
    data_arrays_0_1_rdata_data_data,data_arrays_0_0_rdata_data_data}; // @[src/main/scala/util/package.scala 37:27]
  wire [31:0] rdata_hi = {data_arrays_0_7_rdata_data_data,data_arrays_0_6_rdata_data_data,
    data_arrays_0_5_rdata_data_data,data_arrays_0_4_rdata_data_data}; // @[src/main/scala/util/package.scala 37:27]
  GEN_w1_line #(.COVER_INDEX(693)) line_693 (
    .clock(line_693_clock),
    .reset(line_693_reset),
    .valid(line_693_valid)
  );
  GEN_w1_line #(.COVER_INDEX(694)) line_694 (
    .clock(line_694_clock),
    .reset(line_694_reset),
    .valid(line_694_valid)
  );
  GEN_w1_line #(.COVER_INDEX(695)) line_695 (
    .clock(line_695_clock),
    .reset(line_695_reset),
    .valid(line_695_valid)
  );
  GEN_w1_line #(.COVER_INDEX(696)) line_696 (
    .clock(line_696_clock),
    .reset(line_696_reset),
    .valid(line_696_valid)
  );
  GEN_w1_line #(.COVER_INDEX(697)) line_697 (
    .clock(line_697_clock),
    .reset(line_697_reset),
    .valid(line_697_valid)
  );
  GEN_w1_line #(.COVER_INDEX(698)) line_698 (
    .clock(line_698_clock),
    .reset(line_698_reset),
    .valid(line_698_valid)
  );
  GEN_w1_line #(.COVER_INDEX(699)) line_699 (
    .clock(line_699_clock),
    .reset(line_699_reset),
    .valid(line_699_valid)
  );
  GEN_w1_line #(.COVER_INDEX(700)) line_700 (
    .clock(line_700_clock),
    .reset(line_700_reset),
    .valid(line_700_valid)
  );
  GEN_w1_line #(.COVER_INDEX(701)) line_701 (
    .clock(line_701_clock),
    .reset(line_701_reset),
    .valid(line_701_valid)
  );
  GEN_w1_line #(.COVER_INDEX(702)) line_702 (
    .clock(line_702_clock),
    .reset(line_702_reset),
    .valid(line_702_valid)
  );
  assign data_arrays_0_0_rdata_data_en = data_arrays_0_0_rdata_data_en_pipe_0;
  assign data_arrays_0_0_rdata_data_addr = data_arrays_0_0_rdata_data_addr_pipe_0;
  assign data_arrays_0_0_rdata_data_data = data_arrays_0_0[data_arrays_0_0_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_0_rdata_MPORT_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_0_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_0_rdata_MPORT_mask = io_req_bits_eccMask[0];
  assign data_arrays_0_0_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_1_rdata_data_en = data_arrays_0_1_rdata_data_en_pipe_0;
  assign data_arrays_0_1_rdata_data_addr = data_arrays_0_1_rdata_data_addr_pipe_0;
  assign data_arrays_0_1_rdata_data_data = data_arrays_0_1[data_arrays_0_1_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_1_rdata_MPORT_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_1_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_1_rdata_MPORT_mask = io_req_bits_eccMask[1];
  assign data_arrays_0_1_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_2_rdata_data_en = data_arrays_0_2_rdata_data_en_pipe_0;
  assign data_arrays_0_2_rdata_data_addr = data_arrays_0_2_rdata_data_addr_pipe_0;
  assign data_arrays_0_2_rdata_data_data = data_arrays_0_2[data_arrays_0_2_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_2_rdata_MPORT_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_2_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_2_rdata_MPORT_mask = io_req_bits_eccMask[2];
  assign data_arrays_0_2_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_3_rdata_data_en = data_arrays_0_3_rdata_data_en_pipe_0;
  assign data_arrays_0_3_rdata_data_addr = data_arrays_0_3_rdata_data_addr_pipe_0;
  assign data_arrays_0_3_rdata_data_data = data_arrays_0_3[data_arrays_0_3_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_3_rdata_MPORT_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_3_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_3_rdata_MPORT_mask = io_req_bits_eccMask[3];
  assign data_arrays_0_3_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_4_rdata_data_en = data_arrays_0_4_rdata_data_en_pipe_0;
  assign data_arrays_0_4_rdata_data_addr = data_arrays_0_4_rdata_data_addr_pipe_0;
  assign data_arrays_0_4_rdata_data_data = data_arrays_0_4[data_arrays_0_4_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_4_rdata_MPORT_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_4_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_4_rdata_MPORT_mask = io_req_bits_eccMask[4];
  assign data_arrays_0_4_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_5_rdata_data_en = data_arrays_0_5_rdata_data_en_pipe_0;
  assign data_arrays_0_5_rdata_data_addr = data_arrays_0_5_rdata_data_addr_pipe_0;
  assign data_arrays_0_5_rdata_data_data = data_arrays_0_5[data_arrays_0_5_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_5_rdata_MPORT_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_5_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_5_rdata_MPORT_mask = io_req_bits_eccMask[5];
  assign data_arrays_0_5_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_6_rdata_data_en = data_arrays_0_6_rdata_data_en_pipe_0;
  assign data_arrays_0_6_rdata_data_addr = data_arrays_0_6_rdata_data_addr_pipe_0;
  assign data_arrays_0_6_rdata_data_data = data_arrays_0_6[data_arrays_0_6_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_6_rdata_MPORT_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_6_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_6_rdata_MPORT_mask = io_req_bits_eccMask[6];
  assign data_arrays_0_6_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_7_rdata_data_en = data_arrays_0_7_rdata_data_en_pipe_0;
  assign data_arrays_0_7_rdata_data_addr = data_arrays_0_7_rdata_data_addr_pipe_0;
  assign data_arrays_0_7_rdata_data_data = data_arrays_0_7[data_arrays_0_7_rdata_data_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_7_rdata_MPORT_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_7_rdata_MPORT_addr = io_req_bits_addr[5:3];
  assign data_arrays_0_7_rdata_MPORT_mask = io_req_bits_eccMask[7];
  assign data_arrays_0_7_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign line_693_clock = clock;
  assign line_693_reset = reset;
  assign line_693_valid = _rdata_T ^ line_693_valid_reg;
  assign line_694_clock = clock;
  assign line_694_reset = reset;
  assign line_694_valid = eccMask_0 ^ line_694_valid_reg;
  assign line_695_clock = clock;
  assign line_695_reset = reset;
  assign line_695_valid = eccMask_1 ^ line_695_valid_reg;
  assign line_696_clock = clock;
  assign line_696_reset = reset;
  assign line_696_valid = eccMask_2 ^ line_696_valid_reg;
  assign line_697_clock = clock;
  assign line_697_reset = reset;
  assign line_697_valid = eccMask_3 ^ line_697_valid_reg;
  assign line_698_clock = clock;
  assign line_698_reset = reset;
  assign line_698_valid = eccMask_4 ^ line_698_valid_reg;
  assign line_699_clock = clock;
  assign line_699_reset = reset;
  assign line_699_valid = eccMask_5 ^ line_699_valid_reg;
  assign line_700_clock = clock;
  assign line_700_reset = reset;
  assign line_700_valid = eccMask_6 ^ line_700_valid_reg;
  assign line_701_clock = clock;
  assign line_701_reset = reset;
  assign line_701_valid = eccMask_7 ^ line_701_valid_reg;
  assign line_702_clock = clock;
  assign line_702_reset = reset;
  assign line_702_valid = _rdata_data_T_1 ^ line_702_valid_reg;
  assign io_resp_0 = {rdata_hi,rdata_lo}; // @[src/main/scala/util/package.scala 37:27]
  always @(posedge clock) begin
    if (data_arrays_0_0_rdata_MPORT_en & data_arrays_0_0_rdata_MPORT_mask) begin
      data_arrays_0_0[data_arrays_0_0_rdata_MPORT_addr] <= data_arrays_0_0_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_0_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_0_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_1_rdata_MPORT_en & data_arrays_0_1_rdata_MPORT_mask) begin
      data_arrays_0_1[data_arrays_0_1_rdata_MPORT_addr] <= data_arrays_0_1_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_1_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_1_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_2_rdata_MPORT_en & data_arrays_0_2_rdata_MPORT_mask) begin
      data_arrays_0_2[data_arrays_0_2_rdata_MPORT_addr] <= data_arrays_0_2_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_2_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_2_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_3_rdata_MPORT_en & data_arrays_0_3_rdata_MPORT_mask) begin
      data_arrays_0_3[data_arrays_0_3_rdata_MPORT_addr] <= data_arrays_0_3_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_3_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_3_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_4_rdata_MPORT_en & data_arrays_0_4_rdata_MPORT_mask) begin
      data_arrays_0_4[data_arrays_0_4_rdata_MPORT_addr] <= data_arrays_0_4_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_4_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_4_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_5_rdata_MPORT_en & data_arrays_0_5_rdata_MPORT_mask) begin
      data_arrays_0_5[data_arrays_0_5_rdata_MPORT_addr] <= data_arrays_0_5_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_5_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_5_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_6_rdata_MPORT_en & data_arrays_0_6_rdata_MPORT_mask) begin
      data_arrays_0_6[data_arrays_0_6_rdata_MPORT_addr] <= data_arrays_0_6_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_6_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_6_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    if (data_arrays_0_7_rdata_MPORT_en & data_arrays_0_7_rdata_MPORT_mask) begin
      data_arrays_0_7[data_arrays_0_7_rdata_MPORT_addr] <= data_arrays_0_7_rdata_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_7_rdata_data_en_pipe_0 <= io_req_valid & _rdata_data_T;
    if (io_req_valid & _rdata_data_T) begin
      data_arrays_0_7_rdata_data_addr_pipe_0 <= io_req_bits_addr[5:3];
    end
    line_693_valid_reg <= _rdata_T;
    line_694_valid_reg <= eccMask_0;
    line_695_valid_reg <= eccMask_1;
    line_696_valid_reg <= eccMask_2;
    line_697_valid_reg <= eccMask_3;
    line_698_valid_reg <= eccMask_4;
    line_699_valid_reg <= eccMask_5;
    line_700_valid_reg <= eccMask_6;
    line_701_valid_reg <= eccMask_7;
    line_702_valid_reg <= _rdata_data_T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_0[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_3[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_6[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_9[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_4[initvar] = _RAND_12[7:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_5[initvar] = _RAND_15[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_6[initvar] = _RAND_18[7:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_7[initvar] = _RAND_21[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_arrays_0_0_rdata_data_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_arrays_0_0_rdata_data_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  data_arrays_0_1_rdata_data_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data_arrays_0_1_rdata_data_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  data_arrays_0_2_rdata_data_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  data_arrays_0_2_rdata_data_addr_pipe_0 = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  data_arrays_0_3_rdata_data_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  data_arrays_0_3_rdata_data_addr_pipe_0 = _RAND_11[2:0];
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_4_rdata_data_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_4_rdata_data_addr_pipe_0 = _RAND_14[2:0];
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_5_rdata_data_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_5_rdata_data_addr_pipe_0 = _RAND_17[2:0];
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_6_rdata_data_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_6_rdata_data_addr_pipe_0 = _RAND_20[2:0];
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_7_rdata_data_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_7_rdata_data_addr_pipe_0 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  line_693_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_694_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_695_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_696_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_697_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_698_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_699_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_700_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_701_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_702_valid_reg = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCacheModuleImpl_Anon_2(
  input         clock,
  input         reset,
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [5:0]  io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_bits_write, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [7:0]  io_in_0_bits_eccMask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [5:0]  io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_bits_write, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_2_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [5:0]  io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_2_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_3_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_3_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [5:0]  io_in_3_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [63:0] io_in_3_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_3_bits_wordMask, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [5:0]  io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_write, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [7:0]  io_out_bits_eccMask // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  line_703_clock;
  wire  line_703_reset;
  wire  line_703_valid;
  reg  line_703_valid_reg;
  wire [5:0] _GEN_4 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  wire [63:0] _GEN_6 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  wire  line_704_clock;
  wire  line_704_reset;
  wire  line_704_valid;
  reg  line_704_valid_reg;
  wire [5:0] _GEN_11 = io_in_1_valid ? io_in_1_bits_addr : _GEN_4; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire [63:0] _GEN_13 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_6; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  wire  line_705_clock;
  wire  line_705_reset;
  wire  line_705_valid;
  reg  line_705_valid_reg;
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  GEN_w1_line #(.COVER_INDEX(703)) line_703 (
    .clock(line_703_clock),
    .reset(line_703_reset),
    .valid(line_703_valid)
  );
  GEN_w1_line #(.COVER_INDEX(704)) line_704 (
    .clock(line_704_clock),
    .reset(line_704_reset),
    .valid(line_704_valid)
  );
  GEN_w1_line #(.COVER_INDEX(705)) line_705 (
    .clock(line_705_clock),
    .reset(line_705_reset),
    .valid(line_705_valid)
  );
  assign line_703_clock = clock;
  assign line_703_reset = reset;
  assign line_703_valid = io_in_2_valid ^ line_703_valid_reg;
  assign line_704_clock = clock;
  assign line_704_reset = reset;
  assign line_704_valid = io_in_1_valid ^ line_704_valid_reg;
  assign line_705_clock = clock;
  assign line_705_reset = reset;
  assign line_705_valid = io_in_0_valid ^ line_705_valid_reg;
  assign io_in_1_ready = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_2_ready = ~(io_in_0_valid | io_in_1_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_in_3_ready = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_11; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : io_in_1_valid & io_in_1_bits_write; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_13; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : 8'hff; // @[src/main/scala/chisel3/util/Arbiter.scala 139:26 141:19]
  always @(posedge clock) begin
    line_703_valid_reg <= io_in_2_valid;
    line_704_valid_reg <= io_in_1_valid;
    line_705_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_703_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_704_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_705_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DelayReg(
  input   clock,
  input   reset,
  input   i_valid, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input   i_success, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  output  o_valid, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output  o_success // @[difftest/src/main/scala/util/Delayer.scala 24:13]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_success; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  assign o_valid = REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_success = REG_success; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_valid <= i_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_success <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_success <= i_success; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_success = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper(
  input   clock,
  input   reset,
  input   io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input   io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input   io_bits_success // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_success; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestLrScEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_success(dpic_io_success),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_success = io_bits_success; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DelayReg_1(
  input         clock,
  input         reset,
  input         i_valid, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [63:0] i_addr, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [63:0] i_data, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [7:0]  i_mask, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  output        o_valid, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [63:0] o_addr, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [63:0] o_data, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [7:0]  o_mask // @[difftest/src/main/scala/util/Delayer.scala 24:13]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg  REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [7:0] REG_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_1_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_1_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_1_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [7:0] REG_1_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_2_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_2_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_2_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [7:0] REG_2_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  assign o_valid = REG_2_valid; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_addr = REG_2_addr; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_data = REG_2_data; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_mask = REG_2_mask; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_valid <= i_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_addr <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_addr <= i_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_data <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_data <= i_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_mask <= 8'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_mask <= i_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_1_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_1_valid <= REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_1_addr <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_1_addr <= REG_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_1_data <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_1_data <= REG_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_1_mask <= 8'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_1_mask <= REG_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_2_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_2_valid <= REG_1_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_2_addr <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_2_addr <= REG_1_addr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_2_data <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_2_data <= REG_1_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_2_mask <= 8'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_2_mask <= REG_1_mask; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  REG_data = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  REG_mask = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  REG_1_addr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  REG_1_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  REG_1_mask = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  REG_2_valid = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  REG_2_addr = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  REG_2_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  REG_2_mask = _RAND_11[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_1(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_addr, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_mask // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_addr; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_mask; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestStoreEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_addr(dpic_io_addr),
    .io_data(dpic_io_data),
    .io_mask(dpic_io_mask),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_addr = io_bits_addr; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mask = io_bits_mask; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module AMOALU(
  input         clock,
  input         reset,
  input  [7:0]  io_mask, // @[src/main/scala/rocket/AMOALU.scala 57:14]
  input  [4:0]  io_cmd, // @[src/main/scala/rocket/AMOALU.scala 57:14]
  input  [63:0] io_lhs, // @[src/main/scala/rocket/AMOALU.scala 57:14]
  input  [63:0] io_rhs, // @[src/main/scala/rocket/AMOALU.scala 57:14]
  output [63:0] io_out // @[src/main/scala/rocket/AMOALU.scala 57:14]
);
  wire  max = io_cmd == 5'hd | io_cmd == 5'hf; // @[src/main/scala/rocket/AMOALU.scala 66:33]
  wire  min = io_cmd == 5'hc | io_cmd == 5'he; // @[src/main/scala/rocket/AMOALU.scala 67:33]
  wire  add = io_cmd == 5'h8; // @[src/main/scala/rocket/AMOALU.scala 68:20]
  wire  _logic_and_T = io_cmd == 5'ha; // @[src/main/scala/rocket/AMOALU.scala 69:26]
  wire  logic_and = io_cmd == 5'ha | io_cmd == 5'hb; // @[src/main/scala/rocket/AMOALU.scala 69:38]
  wire  logic_xor = io_cmd == 5'h9 | _logic_and_T; // @[src/main/scala/rocket/AMOALU.scala 70:39]
  wire  _adder_out_mask_T_1 = ~io_mask[3]; // @[src/main/scala/rocket/AMOALU.scala 74:61]
  wire [31:0] _adder_out_mask_T_2 = {_adder_out_mask_T_1, 31'h0}; // @[src/main/scala/rocket/AMOALU.scala 74:77]
  wire [63:0] _adder_out_mask_T_3 = {{32'd0}, _adder_out_mask_T_2}; // @[src/main/scala/rocket/AMOALU.scala 74:96]
  wire [63:0] adder_out_mask = ~_adder_out_mask_T_3; // @[src/main/scala/rocket/AMOALU.scala 74:16]
  wire [63:0] _adder_out_T = io_lhs & adder_out_mask; // @[src/main/scala/rocket/AMOALU.scala 75:13]
  wire [63:0] _adder_out_T_1 = io_rhs & adder_out_mask; // @[src/main/scala/rocket/AMOALU.scala 75:31]
  wire [63:0] adder_out = _adder_out_T + _adder_out_T_1; // @[src/main/scala/rocket/AMOALU.scala 75:21]
  wire [4:0] _less_signed_T = io_cmd & 5'h2; // @[src/main/scala/rocket/AMOALU.scala 88:17]
  wire  less_signed = _less_signed_T == 5'h0; // @[src/main/scala/rocket/AMOALU.scala 88:25]
  wire  _less_T_12 = io_lhs[31:0] < io_rhs[31:0]; // @[src/main/scala/rocket/AMOALU.scala 81:35]
  wire  _less_T_14 = io_lhs[63:32] < io_rhs[63:32] | io_lhs[63:32] == io_rhs[63:32] & _less_T_12; // @[src/main/scala/rocket/AMOALU.scala 82:38]
  wire  _less_T_17 = less_signed ? io_lhs[63] : io_rhs[63]; // @[src/main/scala/rocket/AMOALU.scala 90:58]
  wire  _less_T_18 = io_lhs[63] == io_rhs[63] ? _less_T_14 : _less_T_17; // @[src/main/scala/rocket/AMOALU.scala 90:10]
  wire  _less_T_28 = less_signed ? io_lhs[31] : io_rhs[31]; // @[src/main/scala/rocket/AMOALU.scala 90:58]
  wire  _less_T_29 = io_lhs[31] == io_rhs[31] ? _less_T_12 : _less_T_28; // @[src/main/scala/rocket/AMOALU.scala 90:10]
  wire  less = io_mask[4] ? _less_T_18 : _less_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  _minmax_T = less ? min : max; // @[src/main/scala/rocket/AMOALU.scala 96:23]
  wire [63:0] minmax = _minmax_T ? io_lhs : io_rhs; // @[src/main/scala/rocket/AMOALU.scala 96:19]
  wire [63:0] _logic_T = io_lhs & io_rhs; // @[src/main/scala/rocket/AMOALU.scala 98:27]
  wire [63:0] _logic_T_1 = logic_and ? _logic_T : 64'h0; // @[src/main/scala/rocket/AMOALU.scala 98:8]
  wire [63:0] _logic_T_2 = io_lhs ^ io_rhs; // @[src/main/scala/rocket/AMOALU.scala 99:27]
  wire [63:0] _logic_T_3 = logic_xor ? _logic_T_2 : 64'h0; // @[src/main/scala/rocket/AMOALU.scala 99:8]
  wire [63:0] logic_ = _logic_T_1 | _logic_T_3; // @[src/main/scala/rocket/AMOALU.scala 98:42]
  wire [63:0] _out_T_1 = logic_and | logic_xor ? logic_ : minmax; // @[src/main/scala/rocket/AMOALU.scala 102:8]
  wire [63:0] out = add ? adder_out : _out_T_1; // @[src/main/scala/rocket/AMOALU.scala 101:8]
  wire [7:0] _wmask_T_8 = io_mask[0] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_9 = io_mask[1] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_10 = io_mask[2] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_11 = io_mask[3] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_12 = io_mask[4] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_13 = io_mask[5] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_14 = io_mask[6] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [7:0] _wmask_T_15 = io_mask[7] ? 8'hff : 8'h0; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [63:0] wmask = {_wmask_T_15,_wmask_T_14,_wmask_T_13,_wmask_T_12,_wmask_T_11,_wmask_T_10,_wmask_T_9,_wmask_T_8}; // @[src/main/scala/rocket/AMOALU.scala 105:30]
  wire [63:0] _io_out_T = wmask & out; // @[src/main/scala/rocket/AMOALU.scala 106:19]
  wire [63:0] _io_out_T_1 = ~wmask; // @[src/main/scala/rocket/AMOALU.scala 106:27]
  wire [63:0] _io_out_T_2 = _io_out_T_1 & io_lhs; // @[src/main/scala/rocket/AMOALU.scala 106:34]
  assign io_out = _io_out_T | _io_out_T_2; // @[src/main/scala/rocket/AMOALU.scala 106:25]
endmodule
module DCache(
  input         clock,
  input         reset,
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        io_cpu_req_ready, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_cpu_req_valid, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [39:0] io_cpu_req_bits_addr, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [6:0]  io_cpu_req_bits_tag, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [4:0]  io_cpu_req_bits_cmd, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [1:0]  io_cpu_req_bits_size, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_cpu_req_bits_signed, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [1:0]  io_cpu_req_bits_dprv, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_cpu_req_bits_phys, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_cpu_s1_kill, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [63:0] io_cpu_s1_data_data, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [7:0]  io_cpu_s1_data_mask, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_nack, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_resp_valid, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [39:0] io_cpu_resp_bits_addr, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [6:0]  io_cpu_resp_bits_tag, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [4:0]  io_cpu_resp_bits_cmd, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [1:0]  io_cpu_resp_bits_size, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_resp_bits_signed, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [1:0]  io_cpu_resp_bits_dprv, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_resp_bits_dv, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [63:0] io_cpu_resp_bits_data, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [7:0]  io_cpu_resp_bits_mask, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_resp_bits_replay, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_resp_bits_has_data, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [63:0] io_cpu_resp_bits_data_word_bypass, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [63:0] io_cpu_resp_bits_data_raw, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [63:0] io_cpu_resp_bits_store_data, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_replay_next, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_ma_ld, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_ma_st, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_pf_ld, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_pf_st, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_gf_ld, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_gf_st, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_ae_ld, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_s2_xcpt_ae_st, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_ordered, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_perf_release, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_cpu_perf_grant, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_req_ready, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_ptw_req_valid, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output [26:0] io_ptw_req_bits_bits_addr, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  output        io_ptw_req_bits_bits_need_gpa, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_valid, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_ae_ptw, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_ae_final, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pf, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [43:0] io_ptw_resp_bits_pte_ppn, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_d, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_a, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_g, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_u, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_x, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_w, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_r, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_pte_v, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [1:0]  io_ptw_resp_bits_level, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_resp_bits_homogeneous, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input  [3:0]  io_ptw_ptbr_mode, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_status_mxr, // @[src/main/scala/rocket/HellaCache.scala 234:14]
  input         io_ptw_status_sum // @[src/main/scala/rocket/HellaCache.scala 234:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_reset; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_req_ready; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_req_valid; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_req_bits_passthrough; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [1:0] tlb_io_req_bits_size; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [4:0] tlb_io_req_bits_cmd; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [1:0] tlb_io_req_bits_prv; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_miss; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [31:0] tlb_io_resp_paddr; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_pf_ld; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_pf_st; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_ae_ld; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_ae_st; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_ma_ld; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_ma_st; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_resp_cacheable; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_sfence_valid; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_sfence_bits_rs1; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_sfence_bits_rs2; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_req_ready; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_req_valid; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_req_bits_valid; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_valid; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pf; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [43:0] tlb_io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_status_mxr; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  tlb_io_ptw_status_sum; // @[src/main/scala/rocket/DCache.scala 114:19]
  wire  pma_checker_clock; // @[src/main/scala/rocket/DCache.scala 115:27]
  wire  pma_checker_reset; // @[src/main/scala/rocket/DCache.scala 115:27]
  wire [39:0] pma_checker_io_req_bits_vaddr; // @[src/main/scala/rocket/DCache.scala 115:27]
  wire  lfsr_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  lfsr_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  lfsr_prng_io_increment; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  metaArb_clock; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_reset; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_0_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_0_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_0_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_2_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_2_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_2_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_in_2_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_3_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_3_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_3_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_in_3_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_4_ready; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_4_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_4_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_4_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_in_4_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_5_ready; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_5_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_5_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_5_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_6_ready; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_6_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_6_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_6_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_in_6_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_7_ready; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_7_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_in_7_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_in_7_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_in_7_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_out_valid; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [39:0] metaArb_io_out_bits_addr; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire  metaArb_io_out_bits_idx; // @[src/main/scala/rocket/DCache.scala 119:23]
  wire [27:0] metaArb_io_out_bits_data; // @[src/main/scala/rocket/DCache.scala 119:23]
  reg [27:0] tag_array_0 [0:1]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_s1_meta_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_s1_meta_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [27:0] tag_array_0_s1_meta_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [27:0] tag_array_0_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  tag_array_0_s1_meta_en_pipe_0;
  reg  tag_array_0_s1_meta_addr_pipe_0;
  wire  data_clock; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire  data_reset; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire  data_io_req_valid; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire [5:0] data_io_req_bits_addr; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire  data_io_req_bits_write; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire [63:0] data_io_req_bits_wdata; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire [7:0] data_io_req_bits_eccMask; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire [63:0] data_io_resp_0; // @[src/main/scala/rocket/DCache.scala 129:20]
  wire  dataArb_clock; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_reset; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_0_valid; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [5:0] dataArb_io_in_0_bits_addr; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_0_bits_write; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [63:0] dataArb_io_in_0_bits_wdata; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [7:0] dataArb_io_in_0_bits_eccMask; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_1_ready; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_1_valid; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [5:0] dataArb_io_in_1_bits_addr; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_1_bits_write; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [63:0] dataArb_io_in_1_bits_wdata; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_2_ready; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_2_valid; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [5:0] dataArb_io_in_2_bits_addr; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [63:0] dataArb_io_in_2_bits_wdata; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_3_ready; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_3_valid; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [5:0] dataArb_io_in_3_bits_addr; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [63:0] dataArb_io_in_3_bits_wdata; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_in_3_bits_wordMask; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_out_valid; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [5:0] dataArb_io_out_bits_addr; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  dataArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [63:0] dataArb_io_out_bits_wdata; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire [7:0] dataArb_io_out_bits_eccMask; // @[src/main/scala/rocket/DCache.scala 130:23]
  wire  difftest_delayer_clock; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_reset; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_success; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_success; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_success; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_delayer_1_clock; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_reset; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_i_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_i_addr; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_i_data; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_1_i_mask; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_o_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_o_addr; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_o_data; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_1_o_mask; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_module_1_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_addr; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_1_io_bits_mask; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  amoalus_0_clock; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire  amoalus_0_reset; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire [7:0] amoalus_0_io_mask; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire [4:0] amoalus_0_io_cmd; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire [63:0] amoalus_0_io_lhs; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire [63:0] amoalus_0_io_rhs; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire [63:0] amoalus_0_io_out; // @[src/main/scala/rocket/DCache.scala 979:26]
  wire  _s1_valid_T = io_cpu_req_ready & io_cpu_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  s1_valid; // @[src/main/scala/rocket/DCache.scala 160:25]
  reg [2:0] blockProbeAfterGrantCount; // @[src/main/scala/rocket/DCache.scala 652:42]
  wire  _block_probe_for_core_progress_T = blockProbeAfterGrantCount > 3'h0; // @[src/main/scala/rocket/DCache.scala 750:65]
  reg [6:0] lrscCount; // @[src/main/scala/rocket/DCache.scala 450:26]
  wire  lrscValid = lrscCount > 7'h3; // @[src/main/scala/rocket/DCache.scala 451:29]
  wire  block_probe_for_core_progress = blockProbeAfterGrantCount > 3'h0 | lrscValid; // @[src/main/scala/rocket/DCache.scala 750:71]
  reg  s1_probe; // @[src/main/scala/rocket/DCache.scala 161:25]
  reg  s2_probe; // @[src/main/scala/rocket/DCache.scala 311:25]
  reg [3:0] release_state; // @[src/main/scala/rocket/DCache.scala 206:30]
  wire  releaseInFlight = s1_probe | s2_probe | release_state != 4'h0; // @[src/main/scala/rocket/DCache.scala 312:46]
  reg  release_ack_wait; // @[src/main/scala/rocket/DCache.scala 204:33]
  reg [31:0] release_ack_addr; // @[src/main/scala/rocket/DCache.scala 205:29]
  wire [31:0] _block_probe_for_pending_release_ack_T = auto_out_b_bits_address ^ release_ack_addr; // @[src/main/scala/rocket/DCache.scala 751:88]
  wire  block_probe_for_pending_release_ack = release_ack_wait & _block_probe_for_pending_release_ack_T[20:5] == 16'h0; // @[src/main/scala/rocket/DCache.scala 751:62]
  reg  grantInProgress; // @[src/main/scala/rocket/DCache.scala 651:32]
  wire  block_probe_for_ordering = releaseInFlight | block_probe_for_pending_release_ack | grantInProgress; // @[src/main/scala/rocket/DCache.scala 752:89]
  reg  s2_valid; // @[src/main/scala/rocket/DCache.scala 309:25]
  wire  nodeOut_b_ready = metaArb_io_in_6_ready & ~(block_probe_for_core_progress | block_probe_for_ordering | s1_valid
     | s2_valid); // @[src/main/scala/rocket/DCache.scala 754:44]
  wire  _s1_probe_T = nodeOut_b_ready & auto_out_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [1:0] probe_bits_param; // @[src/main/scala/rocket/DCache.scala 162:29]
  reg [2:0] probe_bits_size; // @[src/main/scala/rocket/DCache.scala 162:29]
  reg  probe_bits_source; // @[src/main/scala/rocket/DCache.scala 162:29]
  reg [31:0] probe_bits_address; // @[src/main/scala/rocket/DCache.scala 162:29]
  wire  line_706_clock;
  wire  line_706_reset;
  wire  line_706_valid;
  reg  line_706_valid_reg;
  wire  s1_valid_masked = s1_valid & ~io_cpu_s1_kill; // @[src/main/scala/rocket/DCache.scala 164:34]
  reg [1:0] s2_probe_state_state; // @[src/main/scala/rocket/DCache.scala 362:33]
  wire [3:0] _T_98 = {probe_bits_param,s2_probe_state_state}; // @[src/main/scala/tilelink/Metadata.scala 120:19]
  wire  _T_155 = 4'h3 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_151 = 4'h2 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_147 = 4'h1 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_143 = 4'h0 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_139 = 4'h7 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_135 = 4'h6 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_131 = 4'h5 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_127 = 4'h4 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_123 = 4'hb == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_119 = 4'ha == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_115 = 4'h9 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_111 = 4'h8 == _T_98; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_128 = _T_127 ? 1'h0 : _T_123; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_132 = _T_131 ? 1'h0 : _T_128; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_136 = _T_135 ? 1'h0 : _T_132; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_144 = _T_143 ? 1'h0 : _T_139 | _T_136; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_148 = _T_147 ? 1'h0 : _T_144; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_152 = _T_151 ? 1'h0 : _T_148; // @[src/main/scala/util/Misc.scala 38:9]
  wire  s2_prb_ack_data = _T_155 | _T_152; // @[src/main/scala/util/Misc.scala 38:9]
  wire  _T_284 = s2_probe_state_state > 2'h0; // @[src/main/scala/tilelink/Metadata.scala 50:45]
  reg [1:0] counter_1; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire  _T_289 = release_state == 4'h1; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_290 = release_state == 4'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_291 = release_state == 4'h9; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_293 = _T_289 | _T_290 | _T_291; // @[src/main/scala/util/package.scala 73:59]
  wire [2:0] _GEN_444 = _T_291 ? 3'h6 : 3'h7; // @[src/main/scala/rocket/DCache.scala 848:52 849:23 854:23]
  wire  _T_288 = release_state == 4'h2; // @[src/main/scala/rocket/DCache.scala 843:25]
  wire  _T_287 = release_state == 4'h3; // @[src/main/scala/rocket/DCache.scala 838:25]
  wire [2:0] _GEN_436 = release_state == 4'h2 ? 3'h5 : 3'h4; // @[src/main/scala/rocket/DCache.scala 843:48 844:21]
  wire [2:0] nodeOut_c_bits_opcode = _T_293 ? _GEN_444 : _GEN_436; // @[src/main/scala/rocket/DCache.scala 847:102]
  wire  beats1_opdata_1 = nodeOut_c_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 102:36]
  wire [2:0] nodeOut_c_bits_size = _T_293 ? 3'h5 : probe_bits_size; // @[src/main/scala/rocket/DCache.scala 847:102]
  wire [11:0] _beats1_decode_T_5 = 12'h1f << nodeOut_c_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beats1_decode_T_7 = ~_beats1_decode_T_5[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beats1_decode_1 = _beats1_decode_T_7[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire [1:0] beats1_1 = beats1_opdata_1 ? beats1_decode_1 : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire  c_last = counter_1 == 2'h1 | beats1_1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  _T_286 = release_state == 4'h5; // @[src/main/scala/rocket/DCache.scala 834:25]
  reg  s2_release_data_valid; // @[src/main/scala/rocket/DCache.scala 786:38]
  wire  c_first = counter_1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  _GEN_385 = s2_prb_ack_data ? s2_release_data_valid & ~(c_first & release_ack_wait) : 1'h1; // @[src/main/scala/rocket/DCache.scala 794:18 812:36]
  wire  _GEN_406 = s2_probe ? _GEN_385 : s2_release_data_valid & ~(c_first & release_ack_wait); // @[src/main/scala/rocket/DCache.scala 794:18 808:21]
  wire  _GEN_423 = release_state == 4'h5 | _GEN_406; // @[src/main/scala/rocket/DCache.scala 834:47 835:22]
  wire  nodeOut_c_valid = release_state == 4'h3 | _GEN_423; // @[src/main/scala/rocket/DCache.scala 838:48 839:22]
  wire  _T_278 = auto_out_c_ready & nodeOut_c_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  releaseDone = c_last & _T_278; // @[src/main/scala/tilelink/Edges.scala 233:22]
  wire  _GEN_383 = _T_284 | ~releaseDone; // @[src/main/scala/rocket/DCache.scala 809:34 814:45 820:19]
  wire  probeNack = s2_prb_ack_data | _GEN_383; // @[src/main/scala/rocket/DCache.scala 809:34 812:36]
  reg [4:0] s1_req_cmd; // @[src/main/scala/rocket/DCache.scala 174:25]
  wire  _s1_read_T = s1_req_cmd == 5'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_1 = s1_req_cmd == 5'h10; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_2 = s1_req_cmd == 5'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_3 = s1_req_cmd == 5'h7; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_6 = _s1_read_T | _s1_read_T_1 | _s1_read_T_2 | _s1_read_T_3; // @[src/main/scala/util/package.scala 73:59]
  wire  _s1_read_T_7 = s1_req_cmd == 5'h4; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_8 = s1_req_cmd == 5'h9; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_9 = s1_req_cmd == 5'ha; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_10 = s1_req_cmd == 5'hb; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_13 = _s1_read_T_7 | _s1_read_T_8 | _s1_read_T_9 | _s1_read_T_10; // @[src/main/scala/util/package.scala 73:59]
  wire  _s1_read_T_14 = s1_req_cmd == 5'h8; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_15 = s1_req_cmd == 5'hc; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_16 = s1_req_cmd == 5'hd; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_17 = s1_req_cmd == 5'he; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_18 = s1_req_cmd == 5'hf; // @[src/main/scala/util/package.scala 16:47]
  wire  _s1_read_T_22 = _s1_read_T_14 | _s1_read_T_15 | _s1_read_T_16 | _s1_read_T_17 | _s1_read_T_18; // @[src/main/scala/util/package.scala 73:59]
  wire  _s1_read_T_23 = _s1_read_T_13 | _s1_read_T_22; // @[src/main/scala/rocket/Consts.scala 83:44]
  wire  s1_read = _s1_read_T_6 | _s1_read_T_23; // @[src/main/scala/rocket/Consts.scala 85:68]
  reg [4:0] s2_req_cmd; // @[src/main/scala/rocket/DCache.scala 317:19]
  wire  _s2_write_T_1 = s2_req_cmd == 5'h11; // @[src/main/scala/rocket/Consts.scala 86:49]
  wire  _s2_write_T_3 = s2_req_cmd == 5'h7; // @[src/main/scala/rocket/Consts.scala 86:66]
  wire  _s2_write_T_5 = s2_req_cmd == 5'h4; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_6 = s2_req_cmd == 5'h9; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_7 = s2_req_cmd == 5'ha; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_8 = s2_req_cmd == 5'hb; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_11 = _s2_write_T_5 | _s2_write_T_6 | _s2_write_T_7 | _s2_write_T_8; // @[src/main/scala/util/package.scala 73:59]
  wire  _s2_write_T_12 = s2_req_cmd == 5'h8; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_13 = s2_req_cmd == 5'hc; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_14 = s2_req_cmd == 5'hd; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_15 = s2_req_cmd == 5'he; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_16 = s2_req_cmd == 5'hf; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_write_T_20 = _s2_write_T_12 | _s2_write_T_13 | _s2_write_T_14 | _s2_write_T_15 | _s2_write_T_16; // @[src/main/scala/util/package.scala 73:59]
  wire  _s2_write_T_21 = _s2_write_T_11 | _s2_write_T_20; // @[src/main/scala/rocket/Consts.scala 83:44]
  wire  s2_write = s2_req_cmd == 5'h1 | s2_req_cmd == 5'h11 | s2_req_cmd == 5'h7 | _s2_write_T_21; // @[src/main/scala/rocket/Consts.scala 86:76]
  reg  pstore1_held; // @[src/main/scala/rocket/DCache.scala 488:29]
  wire  pstore1_valid_likely = s2_valid & s2_write | pstore1_held; // @[src/main/scala/rocket/DCache.scala 489:51]
  reg [39:0] pstore1_addr; // @[src/main/scala/rocket/DCache.scala 477:31]
  reg [39:0] s1_req_addr; // @[src/main/scala/rocket/DCache.scala 174:25]
  wire [39:0] s1_vaddr = {s1_req_addr[39:6],s1_req_addr[5:0]}; // @[src/main/scala/rocket/DCache.scala 175:21]
  wire  _s1_write_T_1 = s1_req_cmd == 5'h11; // @[src/main/scala/rocket/Consts.scala 86:49]
  wire  s1_write = s1_req_cmd == 5'h1 | s1_req_cmd == 5'h11 | _s1_read_T_3 | _s1_read_T_23; // @[src/main/scala/rocket/Consts.scala 86:76]
  reg [7:0] pstore1_mask; // @[src/main/scala/rocket/DCache.scala 480:31]
  wire  _s1_hazard_T_18 = |pstore1_mask[7]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_17 = |pstore1_mask[6]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_16 = |pstore1_mask[5]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_15 = |pstore1_mask[4]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_14 = |pstore1_mask[3]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_13 = |pstore1_mask[2]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_12 = |pstore1_mask[1]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_11 = |pstore1_mask[0]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire [7:0] _s1_hazard_T_19 = {_s1_hazard_T_18,_s1_hazard_T_17,_s1_hazard_T_16,_s1_hazard_T_15,_s1_hazard_T_14,
    _s1_hazard_T_13,_s1_hazard_T_12,_s1_hazard_T_11}; // @[src/main/scala/util/package.scala 37:27]
  wire [7:0] _s1_hazard_T_28 = {_s1_hazard_T_19[7],_s1_hazard_T_19[6],_s1_hazard_T_19[5],_s1_hazard_T_19[4],
    _s1_hazard_T_19[3],_s1_hazard_T_19[2],_s1_hazard_T_19[1],_s1_hazard_T_19[0]}; // @[src/main/scala/rocket/DCache.scala 1179:52]
  reg [1:0] s1_req_size; // @[src/main/scala/rocket/DCache.scala 174:25]
  wire  s1_mask_xwr_upper = s1_req_addr[0] | s1_req_size >= 2'h1; // @[src/main/scala/rocket/AMOALU.scala 19:42]
  wire  s1_mask_xwr_lower = s1_req_addr[0] ? 1'h0 : 1'h1; // @[src/main/scala/rocket/AMOALU.scala 20:22]
  wire [1:0] _s1_mask_xwr_T = {s1_mask_xwr_upper,s1_mask_xwr_lower}; // @[src/main/scala/rocket/AMOALU.scala 21:16]
  wire [1:0] _s1_mask_xwr_upper_T_5 = s1_req_addr[1] ? _s1_mask_xwr_T : 2'h0; // @[src/main/scala/rocket/AMOALU.scala 19:22]
  wire [1:0] _s1_mask_xwr_upper_T_7 = s1_req_size >= 2'h2 ? 2'h3 : 2'h0; // @[src/main/scala/rocket/AMOALU.scala 19:47]
  wire [1:0] s1_mask_xwr_upper_1 = _s1_mask_xwr_upper_T_5 | _s1_mask_xwr_upper_T_7; // @[src/main/scala/rocket/AMOALU.scala 19:42]
  wire [1:0] s1_mask_xwr_lower_1 = s1_req_addr[1] ? 2'h0 : _s1_mask_xwr_T; // @[src/main/scala/rocket/AMOALU.scala 20:22]
  wire [3:0] _s1_mask_xwr_T_1 = {s1_mask_xwr_upper_1,s1_mask_xwr_lower_1}; // @[src/main/scala/rocket/AMOALU.scala 21:16]
  wire [3:0] _s1_mask_xwr_upper_T_9 = s1_req_addr[2] ? _s1_mask_xwr_T_1 : 4'h0; // @[src/main/scala/rocket/AMOALU.scala 19:22]
  wire [3:0] _s1_mask_xwr_upper_T_11 = s1_req_size >= 2'h3 ? 4'hf : 4'h0; // @[src/main/scala/rocket/AMOALU.scala 19:47]
  wire [3:0] s1_mask_xwr_upper_2 = _s1_mask_xwr_upper_T_9 | _s1_mask_xwr_upper_T_11; // @[src/main/scala/rocket/AMOALU.scala 19:42]
  wire [3:0] s1_mask_xwr_lower_2 = s1_req_addr[2] ? 4'h0 : _s1_mask_xwr_T_1; // @[src/main/scala/rocket/AMOALU.scala 20:22]
  wire [7:0] s1_mask_xwr = {s1_mask_xwr_upper_2,s1_mask_xwr_lower_2}; // @[src/main/scala/rocket/AMOALU.scala 21:16]
  wire  _s1_hazard_T_44 = |s1_mask_xwr[7]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_43 = |s1_mask_xwr[6]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_42 = |s1_mask_xwr[5]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_41 = |s1_mask_xwr[4]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_40 = |s1_mask_xwr[3]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_39 = |s1_mask_xwr[2]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_38 = |s1_mask_xwr[1]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_37 = |s1_mask_xwr[0]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire [7:0] _s1_hazard_T_45 = {_s1_hazard_T_44,_s1_hazard_T_43,_s1_hazard_T_42,_s1_hazard_T_41,_s1_hazard_T_40,
    _s1_hazard_T_39,_s1_hazard_T_38,_s1_hazard_T_37}; // @[src/main/scala/util/package.scala 37:27]
  wire [7:0] _s1_hazard_T_54 = {_s1_hazard_T_45[7],_s1_hazard_T_45[6],_s1_hazard_T_45[5],_s1_hazard_T_45[4],
    _s1_hazard_T_45[3],_s1_hazard_T_45[2],_s1_hazard_T_45[1],_s1_hazard_T_45[0]}; // @[src/main/scala/rocket/DCache.scala 1179:52]
  wire [7:0] _s1_hazard_T_55 = _s1_hazard_T_28 & _s1_hazard_T_54; // @[src/main/scala/rocket/DCache.scala 546:38]
  wire [7:0] _s1_hazard_T_57 = pstore1_mask & s1_mask_xwr; // @[src/main/scala/rocket/DCache.scala 546:77]
  wire  _s1_hazard_T_59 = s1_write ? |_s1_hazard_T_55 : |_s1_hazard_T_57; // @[src/main/scala/rocket/DCache.scala 546:8]
  wire  _s1_hazard_T_60 = pstore1_addr[5:3] == s1_vaddr[5:3] & _s1_hazard_T_59; // @[src/main/scala/rocket/DCache.scala 545:65]
  reg  pstore2_valid; // @[src/main/scala/rocket/DCache.scala 485:30]
  reg [39:0] pstore2_addr; // @[src/main/scala/rocket/DCache.scala 508:31]
  reg [7:0] pstore2_storegen_mask; // @[src/main/scala/rocket/DCache.scala 515:19]
  wire  _s1_hazard_T_80 = |pstore2_storegen_mask[7]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_79 = |pstore2_storegen_mask[6]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_78 = |pstore2_storegen_mask[5]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_77 = |pstore2_storegen_mask[4]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_76 = |pstore2_storegen_mask[3]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_75 = |pstore2_storegen_mask[2]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_74 = |pstore2_storegen_mask[1]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _s1_hazard_T_73 = |pstore2_storegen_mask[0]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire [7:0] _s1_hazard_T_81 = {_s1_hazard_T_80,_s1_hazard_T_79,_s1_hazard_T_78,_s1_hazard_T_77,_s1_hazard_T_76,
    _s1_hazard_T_75,_s1_hazard_T_74,_s1_hazard_T_73}; // @[src/main/scala/util/package.scala 37:27]
  wire [7:0] _s1_hazard_T_90 = {_s1_hazard_T_81[7],_s1_hazard_T_81[6],_s1_hazard_T_81[5],_s1_hazard_T_81[4],
    _s1_hazard_T_81[3],_s1_hazard_T_81[2],_s1_hazard_T_81[1],_s1_hazard_T_81[0]}; // @[src/main/scala/rocket/DCache.scala 1179:52]
  wire [7:0] _s1_hazard_T_117 = _s1_hazard_T_90 & _s1_hazard_T_54; // @[src/main/scala/rocket/DCache.scala 546:38]
  wire [7:0] _s1_hazard_T_119 = pstore2_storegen_mask & s1_mask_xwr; // @[src/main/scala/rocket/DCache.scala 546:77]
  wire  _s1_hazard_T_121 = s1_write ? |_s1_hazard_T_117 : |_s1_hazard_T_119; // @[src/main/scala/rocket/DCache.scala 546:8]
  wire  _s1_hazard_T_122 = pstore2_addr[5:3] == s1_vaddr[5:3] & _s1_hazard_T_121; // @[src/main/scala/rocket/DCache.scala 545:65]
  wire  _s1_hazard_T_123 = pstore2_valid & _s1_hazard_T_122; // @[src/main/scala/rocket/DCache.scala 549:21]
  wire  s1_hazard = pstore1_valid_likely & _s1_hazard_T_60 | _s1_hazard_T_123; // @[src/main/scala/rocket/DCache.scala 548:69]
  wire  s1_raw_hazard = s1_read & s1_hazard; // @[src/main/scala/rocket/DCache.scala 550:31]
  wire  _T_243 = s1_valid & s1_raw_hazard; // @[src/main/scala/rocket/DCache.scala 555:18]
  wire [7:0] _s2_valid_no_xcpt_T = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,
    io_cpu_s2_xcpt_gf_ld,io_cpu_s2_xcpt_gf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[src/main/scala/rocket/DCache.scala 310:54]
  wire  s2_valid_no_xcpt = s2_valid & ~(|_s2_valid_no_xcpt_T); // @[src/main/scala/rocket/DCache.scala 310:35]
  reg  s2_not_nacked_in_s1; // @[src/main/scala/rocket/DCache.scala 313:36]
  wire  s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1; // @[src/main/scala/rocket/DCache.scala 315:42]
  wire  _c_cat_T_48 = s2_req_cmd == 5'h6; // @[src/main/scala/rocket/Consts.scala 87:71]
  wire  _c_cat_T_49 = s2_write | s2_req_cmd == 5'h3 | s2_req_cmd == 5'h6; // @[src/main/scala/rocket/Consts.scala 87:64]
  reg [1:0] s2_hit_state_state; // @[src/main/scala/rocket/DCache.scala 364:31]
  wire [3:0] _T_31 = {s2_write,_c_cat_T_49,s2_hit_state_state}; // @[src/main/scala/tilelink/Metadata.scala 58:19]
  wire  _T_89 = 4'h3 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_86 = 4'h2 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_83 = 4'h1 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_80 = 4'h7 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_77 = 4'h6 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_74 = 4'hf == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_71 = 4'he == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_68 = 4'h0 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_65 = 4'h5 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_62 = 4'h4 == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_59 = 4'hd == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  _T_56 = 4'hc == _T_31; // @[src/main/scala/util/Misc.scala 49:20]
  wire  s2_hit = _T_89 | (_T_86 | (_T_83 | (_T_80 | (_T_77 | (_T_74 | _T_71))))); // @[src/main/scala/util/Misc.scala 35:9]
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = s2_valid_masked & s2_hit; // @[src/main/scala/rocket/DCache.scala 375:89]
  wire  _s2_read_T = s2_req_cmd == 5'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_read_T_1 = s2_req_cmd == 5'h10; // @[src/main/scala/util/package.scala 16:47]
  wire  _s2_read_T_6 = _s2_read_T | _s2_read_T_1 | _c_cat_T_48 | _s2_write_T_3; // @[src/main/scala/util/package.scala 73:59]
  wire  s2_read = _s2_read_T_6 | _s2_write_T_21; // @[src/main/scala/rocket/Consts.scala 85:68]
  wire  s2_readwrite = s2_read | s2_write; // @[src/main/scala/rocket/DCache.scala 332:30]
  wire  s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite; // @[src/main/scala/rocket/DCache.scala 396:89]
  wire [1:0] _T_58 = _T_56 ? 2'h1 : 2'h0; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_61 = _T_59 ? 2'h2 : _T_58; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_64 = _T_62 ? 2'h1 : _T_61; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_67 = _T_65 ? 2'h2 : _T_64; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_70 = _T_68 ? 2'h0 : _T_67; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_73 = _T_71 ? 2'h3 : _T_70; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_76 = _T_74 ? 2'h3 : _T_73; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_79 = _T_77 ? 2'h2 : _T_76; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_82 = _T_80 ? 2'h3 : _T_79; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_85 = _T_83 ? 2'h1 : _T_82; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] _T_88 = _T_86 ? 2'h2 : _T_85; // @[src/main/scala/util/Misc.scala 35:36]
  wire [1:0] s2_grow_param = _T_89 ? 2'h3 : _T_88; // @[src/main/scala/util/Misc.scala 35:36]
  wire  _s2_update_meta_T = s2_hit_state_state == s2_grow_param; // @[src/main/scala/tilelink/Metadata.scala 46:46]
  wire  s2_update_meta = ~_s2_update_meta_T; // @[src/main/scala/tilelink/Metadata.scala 47:40]
  wire  _T_223 = io_cpu_s2_nack | s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[src/main/scala/rocket/DCache.scala 424:24]
  wire  s1_readwrite = s1_read | s1_write; // @[src/main/scala/rocket/DCache.scala 190:30]
  wire  s1_flush_line = s1_req_cmd == 5'h5 & s1_req_size[0]; // @[src/main/scala/rocket/DCache.scala 192:50]
  wire  s1_cmd_uses_tlb = s1_readwrite | s1_flush_line | s1_req_cmd == 5'h17; // @[src/main/scala/rocket/DCache.scala 248:55]
  wire  _T_14 = s1_valid & s1_cmd_uses_tlb & tlb_io_resp_miss; // @[src/main/scala/rocket/DCache.scala 254:58]
  wire  _GEN_235 = io_cpu_s2_nack | s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta | _T_14; // @[src/main/scala/rocket/DCache.scala 424:{82,92}]
  wire  _GEN_259 = s1_valid & s1_raw_hazard | _GEN_235; // @[src/main/scala/rocket/DCache.scala 555:{36,46}]
  wire  _GEN_404 = probeNack | _GEN_259; // @[src/main/scala/rocket/DCache.scala 823:{24,34}]
  wire  s1_nack = s2_probe ? _GEN_404 : _GEN_259; // @[src/main/scala/rocket/DCache.scala 808:21]
  wire  _s1_valid_not_nacked_T = ~s1_nack; // @[src/main/scala/rocket/DCache.scala 165:41]
  wire  s1_valid_not_nacked = s1_valid & ~s1_nack; // @[src/main/scala/rocket/DCache.scala 165:38]
  wire  _s0_clk_en_T = ~metaArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 168:43]
  wire  s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 168:40]
  wire [39:0] s0_req_addr = {metaArb_io_out_bits_addr[39:5],io_cpu_req_bits_addr[4:0]}; // @[src/main/scala/rocket/DCache.scala 171:21]
  wire  _T = ~metaArb_io_in_7_ready; // @[src/main/scala/rocket/DCache.scala 173:9]
  wire  line_707_clock;
  wire  line_707_reset;
  wire  line_707_valid;
  reg  line_707_valid_reg;
  wire  s0_req_phys = ~metaArb_io_in_7_ready | io_cpu_req_bits_phys; // @[src/main/scala/rocket/DCache.scala 170:24 173:{34,48}]
  reg [6:0] s1_req_tag; // @[src/main/scala/rocket/DCache.scala 174:25]
  reg  s1_req_signed; // @[src/main/scala/rocket/DCache.scala 174:25]
  reg [1:0] s1_req_dprv; // @[src/main/scala/rocket/DCache.scala 174:25]
  wire  line_708_clock;
  wire  line_708_reset;
  wire  line_708_valid;
  reg  line_708_valid_reg;
  reg [39:0] s1_tlb_req_vaddr; // @[src/main/scala/rocket/DCache.scala 186:29]
  reg  s1_tlb_req_passthrough; // @[src/main/scala/rocket/DCache.scala 186:29]
  reg [1:0] s1_tlb_req_size; // @[src/main/scala/rocket/DCache.scala 186:29]
  reg [4:0] s1_tlb_req_cmd; // @[src/main/scala/rocket/DCache.scala 186:29]
  reg [1:0] s1_tlb_req_prv; // @[src/main/scala/rocket/DCache.scala 186:29]
  wire  line_709_clock;
  wire  line_709_reset;
  wire  line_709_valid;
  reg  line_709_valid_reg;
  wire  s1_sfence = s1_req_cmd == 5'h14 | s1_req_cmd == 5'h15 | s1_req_cmd == 5'h16; // @[src/main/scala/rocket/DCache.scala 191:71]
  reg  s1_flush_valid; // @[src/main/scala/rocket/DCache.scala 193:27]
  reg  cached_grant_wait; // @[src/main/scala/rocket/DCache.scala 201:34]
  reg  resetting; // @[src/main/scala/rocket/DCache.scala 202:26]
  reg  flushCounter; // @[src/main/scala/rocket/DCache.scala 203:29]
  wire  inWriteback = _T_289 | _T_288; // @[src/main/scala/util/package.scala 73:59]
  wire  _io_cpu_req_ready_T = release_state == 4'h0; // @[src/main/scala/rocket/DCache.scala 211:38]
  wire  _io_cpu_req_ready_T_1 = ~cached_grant_wait; // @[src/main/scala/rocket/DCache.scala 211:54]
  reg  uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 214:33]
  reg [39:0] uncachedReqs_0_addr; // @[src/main/scala/rocket/DCache.scala 215:25]
  reg [6:0] uncachedReqs_0_tag; // @[src/main/scala/rocket/DCache.scala 215:25]
  reg [1:0] uncachedReqs_0_size; // @[src/main/scala/rocket/DCache.scala 215:25]
  reg  uncachedReqs_0_signed; // @[src/main/scala/rocket/DCache.scala 215:25]
  wire  _s0_read_T = io_cpu_req_bits_cmd == 5'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_1 = io_cpu_req_bits_cmd == 5'h10; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_2 = io_cpu_req_bits_cmd == 5'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_3 = io_cpu_req_bits_cmd == 5'h7; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_6 = _s0_read_T | _s0_read_T_1 | _s0_read_T_2 | _s0_read_T_3; // @[src/main/scala/util/package.scala 73:59]
  wire  _s0_read_T_7 = io_cpu_req_bits_cmd == 5'h4; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_8 = io_cpu_req_bits_cmd == 5'h9; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_9 = io_cpu_req_bits_cmd == 5'ha; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_10 = io_cpu_req_bits_cmd == 5'hb; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_13 = _s0_read_T_7 | _s0_read_T_8 | _s0_read_T_9 | _s0_read_T_10; // @[src/main/scala/util/package.scala 73:59]
  wire  _s0_read_T_14 = io_cpu_req_bits_cmd == 5'h8; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_15 = io_cpu_req_bits_cmd == 5'hc; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_16 = io_cpu_req_bits_cmd == 5'hd; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_17 = io_cpu_req_bits_cmd == 5'he; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_18 = io_cpu_req_bits_cmd == 5'hf; // @[src/main/scala/util/package.scala 16:47]
  wire  _s0_read_T_22 = _s0_read_T_14 | _s0_read_T_15 | _s0_read_T_16 | _s0_read_T_17 | _s0_read_T_18; // @[src/main/scala/util/package.scala 73:59]
  wire  _s0_read_T_23 = _s0_read_T_13 | _s0_read_T_22; // @[src/main/scala/rocket/Consts.scala 83:44]
  wire  s0_read = _s0_read_T_6 | _s0_read_T_23; // @[src/main/scala/rocket/Consts.scala 85:68]
  wire  _dataArb_io_in_3_valid_res_T = io_cpu_req_bits_cmd == 5'h1; // @[src/main/scala/util/package.scala 16:47]
  wire  _dataArb_io_in_3_valid_res_T_1 = io_cpu_req_bits_cmd == 5'h3; // @[src/main/scala/util/package.scala 16:47]
  wire  _dataArb_io_in_3_valid_res_T_2 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_res_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  dataArb_io_in_3_valid_res = ~_dataArb_io_in_3_valid_res_T_2; // @[src/main/scala/rocket/DCache.scala 1182:15]
  wire  _dataArb_io_in_3_valid_T_26 = io_cpu_req_bits_cmd == 5'h11; // @[src/main/scala/rocket/Consts.scala 86:49]
  wire  _dataArb_io_in_3_valid_T_47 = _dataArb_io_in_3_valid_res_T | io_cpu_req_bits_cmd == 5'h11 | _s0_read_T_3 |
    _s0_read_T_23; // @[src/main/scala/rocket/Consts.scala 86:76]
  wire  _dataArb_io_in_3_valid_T_51 = _dataArb_io_in_3_valid_T_47 & _dataArb_io_in_3_valid_T_26; // @[src/main/scala/rocket/DCache.scala 1188:23]
  wire  _dataArb_io_in_3_valid_T_52 = s0_read | _dataArb_io_in_3_valid_T_51; // @[src/main/scala/rocket/DCache.scala 1187:21]
  wire  _dataArb_io_in_3_valid_T_56 = ~reset; // @[src/main/scala/rocket/DCache.scala 1183:11]
  wire  line_710_clock;
  wire  line_710_reset;
  wire  line_710_valid;
  reg  line_710_valid_reg;
  wire  _dataArb_io_in_3_valid_T_57 = ~(~_dataArb_io_in_3_valid_T_52 | dataArb_io_in_3_valid_res); // @[src/main/scala/rocket/DCache.scala 1183:11]
  wire  line_711_clock;
  wire  line_711_reset;
  wire  line_711_valid;
  reg  line_711_valid_reg;
  wire  _dataArb_io_in_3_valid_T_58 = io_cpu_req_valid & dataArb_io_in_3_valid_res; // @[src/main/scala/rocket/DCache.scala 220:46]
  wire [39:0] _dataArb_io_in_3_bits_addr_T_2 = {io_cpu_req_bits_addr[39:6],io_cpu_req_bits_addr[5:0]}; // @[src/main/scala/rocket/DCache.scala 223:36]
  wire  _T_4 = ~dataArb_io_in_3_ready & s0_read; // @[src/main/scala/rocket/DCache.scala 236:33]
  wire  line_712_clock;
  wire  line_712_reset;
  wire  line_712_valid;
  reg  line_712_valid_reg;
  wire  _GEN_156 = ~dataArb_io_in_3_ready & s0_read ? 1'h0 : release_state == 4'h0 & ~cached_grant_wait &
    _s1_valid_not_nacked_T; // @[src/main/scala/rocket/DCache.scala 211:20 236:{45,64}]
  reg  s1_did_read; // @[src/main/scala/rocket/DCache.scala 237:30]
  wire  line_713_clock;
  wire  line_713_reset;
  wire  line_713_valid;
  reg  line_713_valid_reg;
  reg  s1_read_mask; // @[src/main/scala/rocket/DCache.scala 238:31]
  wire  line_714_clock;
  wire  line_714_reset;
  wire  line_714_valid;
  reg  line_714_valid_reg;
  wire  line_715_clock;
  wire  line_715_reset;
  wire  line_715_valid;
  reg  line_715_valid_reg;
  wire  _GEN_159 = _T ? 1'h0 : _GEN_156; // @[src/main/scala/rocket/DCache.scala 245:{34,53}]
  wire  _T_10 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid & ~io_cpu_req_bits_phys; // @[src/main/scala/rocket/DCache.scala 253:53]
  wire  line_716_clock;
  wire  line_716_reset;
  wire  line_716_valid;
  reg  line_716_valid_reg;
  wire  _GEN_160 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid & ~io_cpu_req_bits_phys ? 1'h0 : _GEN_159; // @[src/main/scala/rocket/DCache.scala 253:{79,98}]
  wire  line_717_clock;
  wire  line_717_reset;
  wire  line_717_valid;
  reg  line_717_valid_reg;
  wire [31:0] s1_paddr = {tlb_io_resp_paddr[31:12],s1_req_addr[11:0]}; // @[src/main/scala/rocket/DCache.scala 276:21]
  wire  _T_19 = metaArb_io_out_valid & metaArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 288:27]
  wire  line_718_clock;
  wire  line_718_reset;
  wire  line_718_valid;
  reg  line_718_valid_reg;
  wire  line_719_clock;
  wire  line_719_reset;
  wire  line_719_valid;
  reg  line_719_valid_reg;
  wire [27:0] _s1_meta_uncorrected_WIRE = tag_array_0_s1_meta_data; // @[src/main/scala/rocket/DCache.scala 293:{80,80}]
  wire [25:0] s1_meta_uncorrected_0_tag = _s1_meta_uncorrected_WIRE[25:0]; // @[src/main/scala/rocket/DCache.scala 293:80]
  wire [1:0] s1_meta_uncorrected_0_coh_state = _s1_meta_uncorrected_WIRE[27:26]; // @[src/main/scala/rocket/DCache.scala 293:80]
  wire [25:0] s1_tag = s1_paddr[31:6]; // @[src/main/scala/rocket/DCache.scala 294:29]
  wire  _s1_meta_hit_way_T_1 = s1_meta_uncorrected_0_tag == s1_tag; // @[src/main/scala/rocket/DCache.scala 295:83]
  wire  _s1_meta_hit_state_T_1 = ~s1_flush_valid; // @[src/main/scala/rocket/DCache.scala 297:62]
  wire [31:0] tl_d_data_encoded_lo = {auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8]
    ,auto_out_d_bits_data[7:0]}; // @[src/main/scala/util/package.scala 37:27]
  wire [31:0] tl_d_data_encoded_hi = {auto_out_d_bits_data[63:56],auto_out_d_bits_data[55:48],auto_out_d_bits_data[47:40
    ],auto_out_d_bits_data[39:32]}; // @[src/main/scala/util/package.scala 37:27]
  wire [63:0] _tl_d_data_encoded_T_8 = {auto_out_d_bits_data[63:56],auto_out_d_bits_data[55:48],auto_out_d_bits_data[47:
    40],auto_out_d_bits_data[39:32],auto_out_d_bits_data[31:24],auto_out_d_bits_data[23:16],auto_out_d_bits_data[15:8],
    auto_out_d_bits_data[7:0]}; // @[src/main/scala/util/package.scala 37:27]
  wire [7:0] _T_23 = ~io_cpu_s1_data_mask; // @[src/main/scala/rocket/DCache.scala 307:71]
  wire [7:0] _T_24 = s1_mask_xwr | _T_23; // @[src/main/scala/rocket/DCache.scala 307:69]
  wire  line_720_clock;
  wire  line_720_reset;
  wire  line_720_valid;
  reg  line_720_valid_reg;
  wire  _T_29 = ~(~(s1_valid_masked & _s1_write_T_1) | &_T_24); // @[src/main/scala/rocket/DCache.scala 307:9]
  wire  line_721_clock;
  wire  line_721_reset;
  wire  line_721_valid;
  reg  line_721_valid_reg;
  reg [39:0] s2_req_addr; // @[src/main/scala/rocket/DCache.scala 317:19]
  reg [6:0] s2_req_tag; // @[src/main/scala/rocket/DCache.scala 317:19]
  reg [1:0] s2_req_size; // @[src/main/scala/rocket/DCache.scala 317:19]
  reg  s2_req_signed; // @[src/main/scala/rocket/DCache.scala 317:19]
  reg [1:0] s2_req_dprv; // @[src/main/scala/rocket/DCache.scala 317:19]
  wire  _s2_cmd_flush_all_T = s2_req_cmd == 5'h5; // @[src/main/scala/rocket/DCache.scala 318:37]
  wire  s2_cmd_flush_line = _s2_cmd_flush_all_T & s2_req_size[0]; // @[src/main/scala/rocket/DCache.scala 319:54]
  reg  s2_tlb_xcpt_pf_ld; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_tlb_xcpt_pf_st; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_tlb_xcpt_ae_ld; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_tlb_xcpt_ae_st; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_tlb_xcpt_ma_ld; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_tlb_xcpt_ma_st; // @[src/main/scala/rocket/DCache.scala 320:24]
  reg  s2_pma_cacheable; // @[src/main/scala/rocket/DCache.scala 321:19]
  reg [39:0] s2_uncached_resp_addr; // @[src/main/scala/rocket/DCache.scala 322:34]
  wire  _T_30 = s1_valid_not_nacked | s1_flush_valid; // @[src/main/scala/rocket/DCache.scala 323:29]
  wire  line_722_clock;
  wire  line_722_reset;
  wire  line_722_valid;
  reg  line_722_valid_reg;
  wire [39:0] _GEN_174 = s1_valid_not_nacked | s1_flush_valid ? {{8'd0}, s1_paddr} : s2_req_addr; // @[src/main/scala/rocket/DCache.scala 323:48 325:17 317:19]
  wire [6:0] _GEN_175 = s1_valid_not_nacked | s1_flush_valid ? s1_req_tag : s2_req_tag; // @[src/main/scala/rocket/DCache.scala 323:48 324:12 317:19]
  wire [4:0] _GEN_176 = s1_valid_not_nacked | s1_flush_valid ? s1_req_cmd : s2_req_cmd; // @[src/main/scala/rocket/DCache.scala 323:48 324:12 317:19]
  wire [1:0] _GEN_177 = s1_valid_not_nacked | s1_flush_valid ? s1_req_size : s2_req_size; // @[src/main/scala/rocket/DCache.scala 323:48 324:12 317:19]
  wire  _GEN_178 = s1_valid_not_nacked | s1_flush_valid ? s1_req_signed : s2_req_signed; // @[src/main/scala/rocket/DCache.scala 323:48 324:12 317:19]
  reg [39:0] s2_vaddr_r; // @[src/main/scala/rocket/DCache.scala 329:31]
  wire  line_723_clock;
  wire  line_723_reset;
  wire  line_723_valid;
  reg  line_723_valid_reg;
  wire [39:0] s2_vaddr = {s2_vaddr_r[39:6],s2_req_addr[5:0]}; // @[src/main/scala/rocket/DCache.scala 329:21]
  reg  s2_flush_valid_pre_tag_ecc; // @[src/main/scala/rocket/DCache.scala 333:43]
  wire  s1_meta_clk_en = _T_30 | s1_probe; // @[src/main/scala/rocket/DCache.scala 335:62]
  wire  line_724_clock;
  wire  line_724_reset;
  wire  line_724_valid;
  reg  line_724_valid_reg;
  wire  line_725_clock;
  wire  line_725_reset;
  wire  line_725_valid;
  reg  line_725_valid_reg;
  reg [27:0] s2_meta_corrected_r; // @[src/main/scala/rocket/DCache.scala 339:61]
  wire  line_726_clock;
  wire  line_726_reset;
  wire  line_726_valid;
  reg  line_726_valid_reg;
  wire [25:0] s2_meta_corrected_0_tag = s2_meta_corrected_r[25:0]; // @[src/main/scala/rocket/DCache.scala 339:99]
  wire [1:0] s2_meta_corrected_0_coh_state = s2_meta_corrected_r[27:26]; // @[src/main/scala/rocket/DCache.scala 339:99]
  wire  s2_data_en = s1_valid | inWriteback | io_cpu_replay_next; // @[src/main/scala/rocket/DCache.scala 344:38]
  wire  s2_data_word_en = inWriteback | s1_did_read & s1_read_mask; // @[src/main/scala/rocket/DCache.scala 345:22]
  wire [63:0] s1_all_data_ways_0 = data_io_resp_0; // @[src/main/scala/rocket/DCache.scala 303:{33,33}]
  wire  s2_data_s1_word_en = ~io_cpu_replay_next ? s2_data_word_en : 1'h1; // @[src/main/scala/rocket/DCache.scala 355:27]
  wire  grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[src/main/scala/util/package.scala 16:47]
  reg  blockUncachedGrant; // @[src/main/scala/rocket/DCache.scala 734:33]
  wire  _T_275 = grantIsUncachedData & (blockUncachedGrant | s1_valid); // @[src/main/scala/rocket/DCache.scala 736:31]
  wire  grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[src/main/scala/rocket/DCache.scala 650:29]
  wire  _T_272 = ~dataArb_io_in_1_ready; // @[src/main/scala/rocket/DCache.scala 706:26]
  wire  _T_273 = grantIsRefill & ~dataArb_io_in_1_ready; // @[src/main/scala/rocket/DCache.scala 706:23]
  wire  _grantIsCached_T = auto_out_d_bits_opcode == 3'h4; // @[src/main/scala/util/package.scala 16:47]
  wire  grantIsCached = _grantIsCached_T | grantIsRefill; // @[src/main/scala/util/package.scala 73:59]
  reg [1:0] counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire  d_first = counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  canAcceptCachedGrant = ~_T_293; // @[src/main/scala/rocket/DCache.scala 654:30]
  wire  _nodeOut_d_ready_T_3 = grantIsCached ? (~d_first | auto_out_e_ready) & canAcceptCachedGrant : 1'h1; // @[src/main/scala/rocket/DCache.scala 655:24]
  wire  _GEN_354 = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : _nodeOut_d_ready_T_3; // @[src/main/scala/rocket/DCache.scala 655:18 706:51 708:20]
  wire  nodeOut_d_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_354; // @[src/main/scala/rocket/DCache.scala 736:68 737:22]
  wire  _T_252 = nodeOut_d_ready & auto_out_d_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_248 = auto_out_d_bits_opcode == 3'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_249 = auto_out_d_bits_opcode == 3'h2; // @[src/main/scala/util/package.scala 16:47]
  wire  grantIsUncached = grantIsUncachedData | _T_248 | _T_249; // @[src/main/scala/util/package.scala 73:59]
  wire [1:0] _GEN_310 = grantIsUncachedData ? 2'h2 : 2'h1; // @[src/main/scala/rocket/DCache.scala 675:34 678:25 301:32]
  wire [1:0] _GEN_319 = grantIsUncached ? _GEN_310 : 2'h1; // @[src/main/scala/rocket/DCache.scala 301:32 668:35]
  wire [1:0] _GEN_332 = grantIsCached ? 2'h1 : _GEN_319; // @[src/main/scala/rocket/DCache.scala 659:26 301:32]
  wire [1:0] s1_data_way = _T_252 ? _GEN_332 : 2'h1; // @[src/main/scala/rocket/DCache.scala 658:24 301:32]
  wire [1:0] _s2_data_T_1 = s2_data_s1_word_en ? s1_data_way : 2'h0; // @[src/main/scala/rocket/DCache.scala 357:28]
  wire [63:0] _s2_data_T_4 = _s2_data_T_1[0] ? s1_all_data_ways_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _s2_data_T_5 = _s2_data_T_1[1] ? _tl_d_data_encoded_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _s2_data_T_6 = _s2_data_T_4 | _s2_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg [63:0] s2_data; // @[src/main/scala/rocket/DCache.scala 357:18]
  wire  line_727_clock;
  wire  line_727_reset;
  wire  line_727_valid;
  reg  line_727_valid_reg;
  wire  line_728_clock;
  wire  line_728_reset;
  wire  line_728_valid;
  reg  line_728_valid_reg;
  wire  line_729_clock;
  wire  line_729_reset;
  wire  line_729_valid;
  reg  line_729_valid_reg;
  wire  line_730_clock;
  wire  line_730_reset;
  wire  line_730_valid;
  reg  line_730_valid_reg;
  wire  line_731_clock;
  wire  line_731_reset;
  wire  line_731_valid;
  reg  line_731_valid_reg;
  wire  line_732_clock;
  wire  line_732_reset;
  wire  line_732_valid;
  reg  line_732_valid_reg;
  wire  s2_hit_valid = s2_hit_state_state > 2'h0; // @[src/main/scala/tilelink/Metadata.scala 50:45]
  wire [31:0] s2_data_corrected_lo = {s2_data[31:24],s2_data[23:16],s2_data[15:8],s2_data[7:0]}; // @[src/main/scala/util/package.scala 37:27]
  wire [31:0] s2_data_corrected_hi = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32]}; // @[src/main/scala/util/package.scala 37:27]
  wire [63:0] s2_data_corrected = {s2_data[63:56],s2_data[55:48],s2_data[47:40],s2_data[39:32],s2_data[31:24],s2_data[23
    :16],s2_data[15:8],s2_data[7:0]}; // @[src/main/scala/util/package.scala 37:27]
  wire  s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line; // @[src/main/scala/rocket/DCache.scala 397:75]
  wire  s2_valid_miss = s2_valid_masked & s2_readwrite & ~s2_hit; // @[src/main/scala/rocket/DCache.scala 401:73]
  wire  s2_uncached = ~s2_pma_cacheable; // @[src/main/scala/rocket/DCache.scala 402:21]
  wire  _s2_valid_cached_miss_T = ~s2_uncached; // @[src/main/scala/rocket/DCache.scala 403:47]
  wire  _s2_valid_cached_miss_T_2 = |uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 403:88]
  wire  s2_valid_cached_miss = s2_valid_miss & ~s2_uncached & ~(|uncachedInFlight_0); // @[src/main/scala/rocket/DCache.scala 403:60]
  wire  s2_want_victimize = s2_valid_cached_miss | s2_valid_flush_line | s2_flush_valid_pre_tag_ecc; // @[src/main/scala/rocket/DCache.scala 405:123]
  wire  _s2_cannot_victimize_T = ~s2_flush_valid_pre_tag_ecc; // @[src/main/scala/rocket/DCache.scala 406:29]
  wire  s2_valid_uncached_pending = s2_valid_miss & s2_uncached & ~(&uncachedInFlight_0); // @[src/main/scala/rocket/DCache.scala 408:64]
  wire  line_733_clock;
  wire  line_733_reset;
  wire  line_733_valid;
  reg  line_733_valid_reg;
  wire [25:0] s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:6] : s2_meta_corrected_0_tag; // @[src/main/scala/rocket/DCache.scala 411:26]
  wire [1:0] s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : s2_meta_corrected_0_coh_state; // @[src/main/scala/rocket/DCache.scala 412:28]
  wire [2:0] _T_113 = _T_111 ? 3'h5 : 3'h0; // @[src/main/scala/util/Misc.scala 38:36]
  wire [2:0] _T_117 = _T_115 ? 3'h2 : _T_113; // @[src/main/scala/util/Misc.scala 38:36]
  wire [2:0] _T_121 = _T_119 ? 3'h1 : _T_117; // @[src/main/scala/util/Misc.scala 38:36]
  wire [2:0] _T_125 = _T_123 ? 3'h1 : _T_121; // @[src/main/scala/util/Misc.scala 38:36]
  wire [2:0] _T_129 = _T_127 ? 3'h5 : _T_125; // @[src/main/scala/util/Misc.scala 38:36]
  wire [2:0] _T_133 = _T_131 ? 3'h4 : _T_129; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_134 = _T_131 ? 2'h1 : 2'h0; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] _T_137 = _T_135 ? 3'h0 : _T_133; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_138 = _T_135 ? 2'h1 : _T_134; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] _T_141 = _T_139 ? 3'h0 : _T_137; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_142 = _T_139 ? 2'h1 : _T_138; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] _T_145 = _T_143 ? 3'h5 : _T_141; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_146 = _T_143 ? 2'h0 : _T_142; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] _T_149 = _T_147 ? 3'h4 : _T_145; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_150 = _T_147 ? 2'h1 : _T_146; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] _T_153 = _T_151 ? 3'h3 : _T_149; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_154 = _T_151 ? 2'h2 : _T_150; // @[src/main/scala/util/Misc.scala 38:63]
  wire [2:0] s2_report_param = _T_155 ? 3'h3 : _T_153; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] probeNewCoh_state = _T_155 ? 2'h2 : _T_154; // @[src/main/scala/util/Misc.scala 38:63]
  wire [3:0] _T_163 = {2'h2,s2_victim_state_state}; // @[src/main/scala/tilelink/Metadata.scala 120:19]
  wire  _T_176 = 4'h8 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire [2:0] _T_178 = _T_176 ? 3'h5 : 3'h0; // @[src/main/scala/util/Misc.scala 38:36]
  wire  _T_180 = 4'h9 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire [2:0] _T_182 = _T_180 ? 3'h2 : _T_178; // @[src/main/scala/util/Misc.scala 38:36]
  wire  _T_184 = 4'ha == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire [2:0] _T_186 = _T_184 ? 3'h1 : _T_182; // @[src/main/scala/util/Misc.scala 38:36]
  wire  _T_188 = 4'hb == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire [2:0] _T_190 = _T_188 ? 3'h1 : _T_186; // @[src/main/scala/util/Misc.scala 38:36]
  wire  _T_192 = 4'h4 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_193 = _T_192 ? 1'h0 : _T_188; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_194 = _T_192 ? 3'h5 : _T_190; // @[src/main/scala/util/Misc.scala 38:36]
  wire  _T_196 = 4'h5 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_197 = _T_196 ? 1'h0 : _T_193; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_198 = _T_196 ? 3'h4 : _T_194; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_199 = _T_196 ? 2'h1 : 2'h0; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_200 = 4'h6 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_201 = _T_200 ? 1'h0 : _T_197; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_202 = _T_200 ? 3'h0 : _T_198; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_203 = _T_200 ? 2'h1 : _T_199; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_204 = 4'h7 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire [2:0] _T_206 = _T_204 ? 3'h0 : _T_202; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_207 = _T_204 ? 2'h1 : _T_203; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_208 = 4'h0 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_209 = _T_208 ? 1'h0 : _T_204 | _T_201; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_210 = _T_208 ? 3'h5 : _T_206; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_211 = _T_208 ? 2'h0 : _T_207; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_212 = 4'h1 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_213 = _T_212 ? 1'h0 : _T_209; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_214 = _T_212 ? 3'h4 : _T_210; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_215 = _T_212 ? 2'h1 : _T_211; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_216 = 4'h2 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  _T_217 = _T_216 ? 1'h0 : _T_213; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] _T_218 = _T_216 ? 3'h3 : _T_214; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] _T_219 = _T_216 ? 2'h2 : _T_215; // @[src/main/scala/util/Misc.scala 38:63]
  wire  _T_220 = 4'h3 == _T_163; // @[src/main/scala/util/Misc.scala 56:20]
  wire  s2_victim_dirty = _T_220 | _T_217; // @[src/main/scala/util/Misc.scala 38:9]
  wire [2:0] s2_shrink_param = _T_220 ? 3'h3 : _T_218; // @[src/main/scala/util/Misc.scala 38:36]
  wire [1:0] voluntaryNewCoh_state = _T_220 ? 2'h2 : _T_219; // @[src/main/scala/util/Misc.scala 38:63]
  wire  s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready; // @[src/main/scala/rocket/DCache.scala 418:57]
  wire  _s2_dont_nack_misc_T_10 = s2_req_cmd == 5'h17; // @[src/main/scala/rocket/DCache.scala 422:17]
  wire  s2_dont_nack_misc = s2_valid_masked & _s2_dont_nack_misc_T_10; // @[src/main/scala/rocket/DCache.scala 419:61]
  wire  _io_cpu_s2_nack_T_4 = ~s2_valid_hit_pre_data_ecc_and_waw; // @[src/main/scala/rocket/DCache.scala 423:89]
  wire  line_734_clock;
  wire  line_734_reset;
  wire  line_734_valid;
  reg  line_734_valid_reg;
  wire [25:0] metaArb_io_in_2_bits_data_meta_tag = s2_req_addr[31:6]; // @[src/main/scala/rocket/HellaCache.scala 299:20 300:14]
  wire  _lrscBackingOff_T = lrscCount > 7'h0; // @[src/main/scala/rocket/DCache.scala 452:34]
  wire  lrscBackingOff = lrscCount > 7'h0 & ~lrscValid; // @[src/main/scala/rocket/DCache.scala 452:40]
  reg [34:0] lrscAddr; // @[src/main/scala/rocket/DCache.scala 453:21]
  wire  lrscAddrMatch = lrscAddr == s2_req_addr[39:5]; // @[src/main/scala/rocket/DCache.scala 454:32]
  wire  s2_sc_fail = _s2_write_T_3 & ~(lrscValid & lrscAddrMatch); // @[src/main/scala/rocket/DCache.scala 455:26]
  wire  _T_227 = s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_48 & _io_cpu_req_ready_T_1 | s2_valid_cached_miss; // @[src/main/scala/rocket/DCache.scala 456:54]
  wire  line_735_clock;
  wire  line_735_reset;
  wire  line_735_valid;
  reg  line_735_valid_reg;
  wire [6:0] _lrscCount_T = s2_hit ? 7'h4f : 7'h0; // @[src/main/scala/rocket/DCache.scala 457:21]
  wire [6:0] _GEN_237 = s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_48 & _io_cpu_req_ready_T_1 | s2_valid_cached_miss
     ? _lrscCount_T : lrscCount; // @[src/main/scala/rocket/DCache.scala 456:99 457:15 450:26]
  wire  line_736_clock;
  wire  line_736_reset;
  wire  line_736_valid;
  reg  line_736_valid_reg;
  wire [6:0] _lrscCount_T_2 = lrscCount - 7'h1; // @[src/main/scala/rocket/DCache.scala 460:51]
  wire  _T_231 = s2_valid_masked & lrscValid; // @[src/main/scala/rocket/DCache.scala 461:29]
  wire  line_737_clock;
  wire  line_737_reset;
  wire  line_737_valid;
  reg  line_737_valid_reg;
  wire  line_738_clock;
  wire  line_738_reset;
  wire  line_738_valid;
  reg  line_738_valid_reg;
  wire  _pstore1_cmd_T = s1_valid_not_nacked & s1_write; // @[src/main/scala/rocket/DCache.scala 476:63]
  reg [4:0] pstore1_cmd; // @[src/main/scala/rocket/DCache.scala 476:30]
  wire  line_739_clock;
  wire  line_739_reset;
  wire  line_739_valid;
  reg  line_739_valid_reg;
  wire  line_740_clock;
  wire  line_740_reset;
  wire  line_740_valid;
  reg  line_740_valid_reg;
  reg [63:0] pstore1_data; // @[src/main/scala/rocket/DCache.scala 478:31]
  wire  line_741_clock;
  wire  line_741_reset;
  wire  line_741_valid;
  reg  line_741_valid_reg;
  wire  line_742_clock;
  wire  line_742_reset;
  wire  line_742_valid;
  reg  line_742_valid_reg;
  wire  line_743_clock;
  wire  line_743_reset;
  wire  line_743_valid;
  reg  line_743_valid_reg;
  wire  _pstore1_rmw_T_51 = s1_write & _s1_write_T_1; // @[src/main/scala/rocket/DCache.scala 1188:23]
  wire  _pstore1_rmw_T_52 = s1_read | _pstore1_rmw_T_51; // @[src/main/scala/rocket/DCache.scala 1187:21]
  reg  pstore1_rmw_r; // @[src/main/scala/rocket/DCache.scala 482:44]
  wire  line_744_clock;
  wire  line_744_reset;
  wire  line_744_valid;
  reg  line_744_valid_reg;
  wire  _pstore1_merge_T = s2_valid_hit_pre_data_ecc_and_waw & s2_write; // @[src/main/scala/rocket/DCache.scala 474:46]
  wire  _pstore1_merge_T_2 = s2_valid_hit_pre_data_ecc_and_waw & s2_write & ~s2_sc_fail; // @[src/main/scala/rocket/DCache.scala 474:58]
  wire  line_745_clock;
  wire  line_745_reset;
  wire  line_745_valid;
  reg  line_745_valid_reg;
  wire  line_746_clock;
  wire  line_746_reset;
  wire  line_746_valid;
  reg  line_746_valid_reg;
  wire  pstore_drain_opportunistic = ~_dataArb_io_in_3_valid_T_58; // @[src/main/scala/rocket/DCache.scala 486:36]
  reg  pstore_drain_on_miss_REG; // @[src/main/scala/rocket/DCache.scala 487:56]
  wire  pstore_drain_on_miss = releaseInFlight | pstore_drain_on_miss_REG; // @[src/main/scala/rocket/DCache.scala 487:46]
  wire  pstore1_valid = _pstore1_merge_T_2 | pstore1_held; // @[src/main/scala/rocket/DCache.scala 491:38]
  wire  pstore_drain_structural = pstore1_valid_likely & pstore2_valid & (s1_valid & s1_write | pstore1_rmw_r); // @[src/main/scala/rocket/DCache.scala 493:71]
  wire  _T_235 = _pstore1_merge_T | pstore1_held; // @[src/main/scala/rocket/DCache.scala 490:96]
  wire  line_747_clock;
  wire  line_747_reset;
  wire  line_747_valid;
  reg  line_747_valid_reg;
  wire  _T_240 = ~(pstore1_rmw_r | _T_235 == pstore1_valid); // @[src/main/scala/rocket/DCache.scala 494:9]
  wire  line_748_clock;
  wire  line_748_reset;
  wire  line_748_valid;
  reg  line_748_valid_reg;
  wire  _pstore_drain_T_10 = (_T_235 & ~pstore1_rmw_r | pstore2_valid) & (pstore_drain_opportunistic |
    pstore_drain_on_miss); // @[src/main/scala/rocket/DCache.scala 502:76]
  wire  pstore_drain = pstore_drain_structural | _pstore_drain_T_10; // @[src/main/scala/rocket/DCache.scala 501:44]
  wire  _pstore1_held_T_9 = ~pstore_drain; // @[src/main/scala/rocket/DCache.scala 505:91]
  wire  advance_pstore1 = pstore1_valid & pstore2_valid == pstore_drain; // @[src/main/scala/rocket/DCache.scala 506:61]
  wire  line_749_clock;
  wire  line_749_reset;
  wire  line_749_valid;
  reg  line_749_valid_reg;
  wire  line_750_clock;
  wire  line_750_reset;
  wire  line_750_valid;
  reg  line_750_valid_reg;
  wire [63:0] pstore1_storegen_data = amoalus_0_io_out; // @[src/main/scala/rocket/DCache.scala 481:42 986:27]
  reg [7:0] pstore2_storegen_data_r; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_751_clock;
  wire  line_751_reset;
  wire  line_751_valid;
  reg  line_751_valid_reg;
  reg [7:0] pstore2_storegen_data_r_1; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_752_clock;
  wire  line_752_reset;
  wire  line_752_valid;
  reg  line_752_valid_reg;
  reg [7:0] pstore2_storegen_data_r_2; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_753_clock;
  wire  line_753_reset;
  wire  line_753_valid;
  reg  line_753_valid_reg;
  reg [7:0] pstore2_storegen_data_r_3; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_754_clock;
  wire  line_754_reset;
  wire  line_754_valid;
  reg  line_754_valid_reg;
  reg [7:0] pstore2_storegen_data_r_4; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_755_clock;
  wire  line_755_reset;
  wire  line_755_valid;
  reg  line_755_valid_reg;
  reg [7:0] pstore2_storegen_data_r_5; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_756_clock;
  wire  line_756_reset;
  wire  line_756_valid;
  reg  line_756_valid_reg;
  reg [7:0] pstore2_storegen_data_r_6; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_757_clock;
  wire  line_757_reset;
  wire  line_757_valid;
  reg  line_757_valid_reg;
  reg [7:0] pstore2_storegen_data_r_7; // @[src/main/scala/rocket/DCache.scala 512:22]
  wire  line_758_clock;
  wire  line_758_reset;
  wire  line_758_valid;
  reg  line_758_valid_reg;
  wire [63:0] pstore2_storegen_data = {pstore2_storegen_data_r_7,pstore2_storegen_data_r_6,pstore2_storegen_data_r_5,
    pstore2_storegen_data_r_4,pstore2_storegen_data_r_3,pstore2_storegen_data_r_2,pstore2_storegen_data_r_1,
    pstore2_storegen_data_r}; // @[src/main/scala/util/package.scala 37:27]
  wire  line_759_clock;
  wire  line_759_reset;
  wire  line_759_valid;
  reg  line_759_valid_reg;
  wire [7:0] _pstore2_storegen_mask_mask_T = ~pstore1_mask; // @[src/main/scala/rocket/DCache.scala 518:37]
  wire [7:0] _pstore2_storegen_mask_mask_T_2 = ~_pstore2_storegen_mask_mask_T; // @[src/main/scala/rocket/DCache.scala 518:15]
  wire [39:0] _dataArb_io_in_0_bits_addr_T = pstore2_valid ? pstore2_addr : pstore1_addr; // @[src/main/scala/rocket/DCache.scala 533:36]
  wire [63:0] _dataArb_io_in_0_bits_wdata_T = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[src/main/scala/rocket/DCache.scala 535:63]
  wire [31:0] dataArb_io_in_0_bits_wdata_lo = {_dataArb_io_in_0_bits_wdata_T[31:24],_dataArb_io_in_0_bits_wdata_T[23:16]
    ,_dataArb_io_in_0_bits_wdata_T[15:8],_dataArb_io_in_0_bits_wdata_T[7:0]}; // @[src/main/scala/util/package.scala 37:27]
  wire [31:0] dataArb_io_in_0_bits_wdata_hi = {_dataArb_io_in_0_bits_wdata_T[63:56],_dataArb_io_in_0_bits_wdata_T[55:48]
    ,_dataArb_io_in_0_bits_wdata_T[47:40],_dataArb_io_in_0_bits_wdata_T[39:32]}; // @[src/main/scala/util/package.scala 37:27]
  wire [7:0] _dataArb_io_in_0_bits_eccMask_T = pstore2_valid ? pstore2_storegen_mask : pstore1_mask; // @[src/main/scala/rocket/DCache.scala 541:47]
  wire  _dataArb_io_in_0_bits_eccMask_T_9 = |_dataArb_io_in_0_bits_eccMask_T[0]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_10 = |_dataArb_io_in_0_bits_eccMask_T[1]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_11 = |_dataArb_io_in_0_bits_eccMask_T[2]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_12 = |_dataArb_io_in_0_bits_eccMask_T[3]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_13 = |_dataArb_io_in_0_bits_eccMask_T[4]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_14 = |_dataArb_io_in_0_bits_eccMask_T[5]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_15 = |_dataArb_io_in_0_bits_eccMask_T[6]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire  _dataArb_io_in_0_bits_eccMask_T_16 = |_dataArb_io_in_0_bits_eccMask_T[7]; // @[src/main/scala/rocket/DCache.scala 1178:66]
  wire [3:0] dataArb_io_in_0_bits_eccMask_lo = {_dataArb_io_in_0_bits_eccMask_T_12,_dataArb_io_in_0_bits_eccMask_T_11,
    _dataArb_io_in_0_bits_eccMask_T_10,_dataArb_io_in_0_bits_eccMask_T_9}; // @[src/main/scala/util/package.scala 37:27]
  wire [3:0] dataArb_io_in_0_bits_eccMask_hi = {_dataArb_io_in_0_bits_eccMask_T_16,_dataArb_io_in_0_bits_eccMask_T_15,
    _dataArb_io_in_0_bits_eccMask_T_14,_dataArb_io_in_0_bits_eccMask_T_13}; // @[src/main/scala/util/package.scala 37:27]
  wire  line_760_clock;
  wire  line_760_reset;
  wire  line_760_valid;
  reg  line_760_valid_reg;
  wire  _a_source_T = ~uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 561:34]
  wire [1:0] _a_source_T_1 = {_a_source_T, 1'h0}; // @[src/main/scala/rocket/DCache.scala 561:59]
  wire  a_source = _a_source_T_1[0] ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [39:0] acquire_address = {s2_req_addr[39:5], 5'h0}; // @[src/main/scala/rocket/DCache.scala 562:49]
  wire [22:0] a_mask = {{15'd0}, pstore1_mask}; // @[src/main/scala/rocket/DCache.scala 566:29]
  wire [2:0] _get_a_mask_sizeOH_T = {{1'd0}, s2_req_size}; // @[src/main/scala/util/Misc.scala 202:34]
  wire [1:0] get_a_mask_sizeOH_shiftAmount = _get_a_mask_sizeOH_T[1:0]; // @[src/main/scala/chisel3/util/OneHot.scala 64:49]
  wire [3:0] _get_a_mask_sizeOH_T_1 = 4'h1 << get_a_mask_sizeOH_shiftAmount; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire [2:0] get_a_mask_sizeOH = _get_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[src/main/scala/util/Misc.scala 202:81]
  wire  _get_a_mask_T = s2_req_size >= 2'h3; // @[src/main/scala/util/Misc.scala 206:21]
  wire  get_a_mask_size = get_a_mask_sizeOH[2]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  get_a_mask_bit = s2_req_addr[2]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  get_a_mask_nbit = ~get_a_mask_bit; // @[src/main/scala/util/Misc.scala 211:20]
  wire  get_a_mask_acc = _get_a_mask_T | get_a_mask_size & get_a_mask_nbit; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_acc_1 = _get_a_mask_T | get_a_mask_size & get_a_mask_bit; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_size_1 = get_a_mask_sizeOH[1]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  get_a_mask_bit_1 = s2_req_addr[1]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  get_a_mask_nbit_1 = ~get_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 211:20]
  wire  get_a_mask_eq_2 = get_a_mask_nbit & get_a_mask_nbit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_2 = get_a_mask_acc | get_a_mask_size_1 & get_a_mask_eq_2; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_3 = get_a_mask_nbit & get_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_3 = get_a_mask_acc | get_a_mask_size_1 & get_a_mask_eq_3; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_4 = get_a_mask_bit & get_a_mask_nbit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_4 = get_a_mask_acc_1 | get_a_mask_size_1 & get_a_mask_eq_4; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_5 = get_a_mask_bit & get_a_mask_bit_1; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_5 = get_a_mask_acc_1 | get_a_mask_size_1 & get_a_mask_eq_5; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_size_2 = get_a_mask_sizeOH[0]; // @[src/main/scala/util/Misc.scala 209:26]
  wire  get_a_mask_bit_2 = s2_req_addr[0]; // @[src/main/scala/util/Misc.scala 210:26]
  wire  get_a_mask_nbit_2 = ~get_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 211:20]
  wire  get_a_mask_eq_6 = get_a_mask_eq_2 & get_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_6 = get_a_mask_acc_2 | get_a_mask_size_2 & get_a_mask_eq_6; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_7 = get_a_mask_eq_2 & get_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_7 = get_a_mask_acc_2 | get_a_mask_size_2 & get_a_mask_eq_7; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_8 = get_a_mask_eq_3 & get_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_8 = get_a_mask_acc_3 | get_a_mask_size_2 & get_a_mask_eq_8; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_9 = get_a_mask_eq_3 & get_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_9 = get_a_mask_acc_3 | get_a_mask_size_2 & get_a_mask_eq_9; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_10 = get_a_mask_eq_4 & get_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_10 = get_a_mask_acc_4 | get_a_mask_size_2 & get_a_mask_eq_10; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_11 = get_a_mask_eq_4 & get_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_11 = get_a_mask_acc_4 | get_a_mask_size_2 & get_a_mask_eq_11; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_12 = get_a_mask_eq_5 & get_a_mask_nbit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_12 = get_a_mask_acc_5 | get_a_mask_size_2 & get_a_mask_eq_12; // @[src/main/scala/util/Misc.scala 215:29]
  wire  get_a_mask_eq_13 = get_a_mask_eq_5 & get_a_mask_bit_2; // @[src/main/scala/util/Misc.scala 214:27]
  wire  get_a_mask_acc_13 = get_a_mask_acc_5 | get_a_mask_size_2 & get_a_mask_eq_13; // @[src/main/scala/util/Misc.scala 215:29]
  wire [7:0] get_mask = {get_a_mask_acc_13,get_a_mask_acc_12,get_a_mask_acc_11,get_a_mask_acc_10,get_a_mask_acc_9,
    get_a_mask_acc_8,get_a_mask_acc_7,get_a_mask_acc_6}; // @[src/main/scala/util/Misc.scala 222:10]
  wire [39:0] _GEN_478 = {{8'd0}, release_ack_addr}; // @[src/main/scala/rocket/DCache.scala 590:43]
  wire [39:0] _tl_out_a_valid_T_1 = s2_req_addr ^ _GEN_478; // @[src/main/scala/rocket/DCache.scala 590:43]
  wire  _tl_out_a_valid_T_5 = ~(release_ack_wait & _tl_out_a_valid_T_1[20:5] == 16'h0); // @[src/main/scala/rocket/DCache.scala 590:8]
  wire  _tl_out_a_valid_T_6 = s2_valid_cached_miss & _tl_out_a_valid_T_5; // @[src/main/scala/rocket/DCache.scala 589:29]
  wire  _tl_out_a_valid_T_7 = ~release_ack_wait; // @[src/main/scala/rocket/DCache.scala 591:47]
  wire  _tl_out_a_valid_T_10 = ~s2_victim_dirty; // @[src/main/scala/rocket/DCache.scala 591:91]
  wire  _tl_out_a_valid_T_12 = _tl_out_a_valid_T_6 & _tl_out_a_valid_T_10; // @[src/main/scala/rocket/DCache.scala 590:127]
  wire  tl_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12; // @[src/main/scala/rocket/DCache.scala 588:32]
  wire  line_761_clock;
  wire  line_761_reset;
  wire  line_761_valid;
  reg  line_761_valid_reg;
  wire  _atomics_T_6 = ~(~(tl_out_a_valid & s2_read & s2_write & s2_uncached)); // @[src/main/scala/rocket/DCache.scala 583:12]
  wire  line_762_clock;
  wire  line_762_reset;
  wire  line_762_valid;
  reg  line_762_valid_reg;
  wire [2:0] _tl_out_a_bits_T_6_size = ~s2_read ? _get_a_mask_sizeOH_T : 3'h0; // @[src/main/scala/rocket/DCache.scala 595:8]
  wire  _tl_out_a_bits_T_6_source = ~s2_read & a_source; // @[src/main/scala/rocket/DCache.scala 595:8]
  wire [31:0] put_address = s2_req_addr[31:0]; // @[src/main/scala/tilelink/Edges.scala 480:17 485:15]
  wire [31:0] _tl_out_a_bits_T_6_address = ~s2_read ? put_address : 32'h0; // @[src/main/scala/rocket/DCache.scala 595:8]
  wire [7:0] _tl_out_a_bits_T_6_mask = ~s2_read ? get_mask : 8'h0; // @[src/main/scala/rocket/DCache.scala 595:8]
  wire [63:0] _tl_out_a_bits_T_6_data = ~s2_read ? pstore1_data : 64'h0; // @[src/main/scala/rocket/DCache.scala 595:8]
  wire [2:0] _tl_out_a_bits_T_7_opcode = _s2_write_T_1 ? 3'h1 : 3'h0; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire [2:0] _tl_out_a_bits_T_7_size = _s2_write_T_1 ? _get_a_mask_sizeOH_T : _tl_out_a_bits_T_6_size; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire  _tl_out_a_bits_T_7_source = _s2_write_T_1 ? a_source : _tl_out_a_bits_T_6_source; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire [31:0] _tl_out_a_bits_T_7_address = _s2_write_T_1 ? put_address : _tl_out_a_bits_T_6_address; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire [7:0] putpartial_mask = a_mask[7:0]; // @[src/main/scala/tilelink/Edges.scala 500:17 508:15]
  wire [7:0] _tl_out_a_bits_T_7_mask = _s2_write_T_1 ? putpartial_mask : _tl_out_a_bits_T_6_mask; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire [63:0] _tl_out_a_bits_T_7_data = _s2_write_T_1 ? pstore1_data : _tl_out_a_bits_T_6_data; // @[src/main/scala/rocket/DCache.scala 594:8]
  wire [2:0] _tl_out_a_bits_T_8_opcode = ~s2_write ? 3'h4 : _tl_out_a_bits_T_7_opcode; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire [2:0] _tl_out_a_bits_T_8_size = ~s2_write ? _get_a_mask_sizeOH_T : _tl_out_a_bits_T_7_size; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire  _tl_out_a_bits_T_8_source = ~s2_write ? a_source : _tl_out_a_bits_T_7_source; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire [31:0] _tl_out_a_bits_T_8_address = ~s2_write ? put_address : _tl_out_a_bits_T_7_address; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire [7:0] _tl_out_a_bits_T_8_mask = ~s2_write ? get_mask : _tl_out_a_bits_T_7_mask; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire [63:0] _tl_out_a_bits_T_8_data = ~s2_write ? 64'h0 : _tl_out_a_bits_T_7_data; // @[src/main/scala/rocket/DCache.scala 593:8]
  wire [2:0] tl_out_a_bits_a_param = {{1'd0}, s2_grow_param}; // @[src/main/scala/tilelink/Edges.scala 346:17 348:15]
  wire [31:0] tl_out_a_bits_a_address = acquire_address[31:0]; // @[src/main/scala/tilelink/Edges.scala 346:17 351:15]
  wire [1:0] _a_sel_T = 2'h1 << a_source; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  a_sel = _a_sel_T[1]; // @[src/main/scala/rocket/DCache.scala 614:66]
  wire  _T_244 = auto_out_a_ready & tl_out_a_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_763_clock;
  wire  line_763_reset;
  wire  line_763_valid;
  reg  line_763_valid_reg;
  wire  line_764_clock;
  wire  line_764_reset;
  wire  line_764_valid;
  reg  line_764_valid_reg;
  wire  line_765_clock;
  wire  line_765_reset;
  wire  line_765_valid;
  reg  line_765_valid_reg;
  wire  _GEN_260 = a_sel | uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 618:18 619:13 214:33]
  wire  line_766_clock;
  wire  line_766_reset;
  wire  line_766_valid;
  reg  line_766_valid_reg;
  wire  _GEN_273 = s2_uncached ? _GEN_260 : uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 616:24 214:33]
  wire  _GEN_286 = s2_uncached ? cached_grant_wait : 1'h1; // @[src/main/scala/rocket/DCache.scala 616:24 201:34 625:25]
  wire  _GEN_288 = _T_244 ? _GEN_273 : uncachedInFlight_0; // @[src/main/scala/rocket/DCache.scala 615:24 214:33]
  wire  _GEN_301 = _T_244 ? _GEN_286 : cached_grant_wait; // @[src/main/scala/rocket/DCache.scala 615:24 201:34]
  wire [11:0] _beats1_decode_T_1 = 12'h1f << auto_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beats1_decode = _beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire  beats1_opdata = auto_out_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  wire [1:0] beats1 = beats1_opdata ? beats1_decode : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  wire [1:0] counter1 = counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  d_last = counter == 2'h1 | beats1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  d_done = d_last & _T_252; // @[src/main/scala/tilelink/Edges.scala 233:22]
  wire [1:0] _count_T = ~counter1; // @[src/main/scala/tilelink/Edges.scala 234:27]
  wire [1:0] count = beats1 & _count_T; // @[src/main/scala/tilelink/Edges.scala 234:25]
  wire  line_767_clock;
  wire  line_767_reset;
  wire  line_767_valid;
  reg  line_767_valid_reg;
  wire [4:0] d_address_inc = {count, 3'h0}; // @[src/main/scala/tilelink/Edges.scala 269:29]
  wire  _tl_d_data_encoded_T_11 = ~grantIsUncached; // @[src/main/scala/rocket/DCache.scala 647:129]
  wire  grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[src/main/scala/rocket/DCache.scala 649:32]
  wire  line_768_clock;
  wire  line_768_reset;
  wire  line_768_valid;
  reg  line_768_valid_reg;
  wire [2:0] _blockProbeAfterGrantCount_T_1 = blockProbeAfterGrantCount - 3'h1; // @[src/main/scala/rocket/DCache.scala 653:99]
  wire [2:0] _GEN_304 = _block_probe_for_core_progress_T ? _blockProbeAfterGrantCount_T_1 : blockProbeAfterGrantCount; // @[src/main/scala/rocket/DCache.scala 652:42 653:{42,70}]
  wire [1:0] _uncachedRespIdxOH_T = 2'h1 << auto_out_d_bits_source; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  uncachedRespIdxOH = _uncachedRespIdxOH_T[1]; // @[src/main/scala/rocket/DCache.scala 656:90]
  wire  line_769_clock;
  wire  line_769_reset;
  wire  line_769_valid;
  reg  line_769_valid_reg;
  wire  line_770_clock;
  wire  line_770_reset;
  wire  line_770_valid;
  reg  line_770_valid_reg;
  wire  line_771_clock;
  wire  line_771_reset;
  wire  line_771_valid;
  reg  line_771_valid_reg;
  wire  line_772_clock;
  wire  line_772_reset;
  wire  line_772_valid;
  reg  line_772_valid_reg;
  wire  line_773_clock;
  wire  line_773_reset;
  wire  line_773_valid;
  reg  line_773_valid_reg;
  wire  line_774_clock;
  wire  line_774_reset;
  wire  line_774_valid;
  reg  line_774_valid_reg;
  wire  line_775_clock;
  wire  line_775_reset;
  wire  line_775_valid;
  reg  line_775_valid_reg;
  wire  _T_257 = uncachedRespIdxOH & d_last; // @[src/main/scala/rocket/DCache.scala 670:17]
  wire  line_776_clock;
  wire  line_776_reset;
  wire  line_776_valid;
  reg  line_776_valid_reg;
  wire  line_777_clock;
  wire  line_777_reset;
  wire  line_777_valid;
  reg  line_777_valid_reg;
  wire  line_778_clock;
  wire  line_778_reset;
  wire  line_778_valid;
  reg  line_778_valid_reg;
  wire  _GEN_309 = uncachedRespIdxOH & d_last ? 1'h0 : _GEN_288; // @[src/main/scala/rocket/DCache.scala 670:28 672:13]
  wire  line_779_clock;
  wire  line_779_reset;
  wire  line_779_valid;
  reg  line_779_valid_reg;
  wire [31:0] s2_req_addr_dontCareBits = {s1_paddr[31:3], 3'h0}; // @[src/main/scala/rocket/DCache.scala 685:55]
  wire [31:0] _GEN_479 = {{29'd0}, uncachedReqs_0_addr[2:0]}; // @[src/main/scala/rocket/DCache.scala 686:26]
  wire [31:0] _s2_req_addr_T_1 = s2_req_addr_dontCareBits | _GEN_479; // @[src/main/scala/rocket/DCache.scala 686:26]
  wire  line_780_clock;
  wire  line_780_reset;
  wire  line_780_valid;
  reg  line_780_valid_reg;
  wire  line_781_clock;
  wire  line_781_reset;
  wire  line_781_valid;
  reg  line_781_valid_reg;
  wire  line_782_clock;
  wire  line_782_reset;
  wire  line_782_valid;
  reg  line_782_valid_reg;
  wire  line_783_clock;
  wire  line_783_reset;
  wire  line_783_valid;
  reg  line_783_valid_reg;
  wire  _GEN_317 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[src/main/scala/rocket/DCache.scala 691:36 693:24 204:33]
  wire  _GEN_326 = grantIsUncached ? release_ack_wait : _GEN_317; // @[src/main/scala/rocket/DCache.scala 204:33 668:35]
  wire  _GEN_330 = grantIsCached & d_last; // @[src/main/scala/rocket/DCache.scala 659:26 src/main/scala/util/Replacement.scala 38:11]
  wire  _GEN_339 = grantIsCached ? release_ack_wait : _GEN_326; // @[src/main/scala/rocket/DCache.scala 659:26 204:33]
  wire  _GEN_352 = _T_252 ? _GEN_339 : release_ack_wait; // @[src/main/scala/rocket/DCache.scala 658:24 204:33]
  wire  nodeOut_e_valid = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : auto_out_d_valid & d_first & grantIsCached &
    canAcceptCachedGrant; // @[src/main/scala/rocket/DCache.scala 698:18 706:51 707:20]
  wire  _T_264 = auto_out_e_ready & nodeOut_e_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_784_clock;
  wire  line_784_reset;
  wire  line_784_valid;
  reg  line_784_valid_reg;
  wire  _T_271 = ~(_T_264 == (_T_252 & d_first & grantIsCached)); // @[src/main/scala/rocket/DCache.scala 700:9]
  wire  line_785_clock;
  wire  line_785_reset;
  wire  line_785_valid;
  reg  line_785_valid_reg;
  wire  line_786_clock;
  wire  line_786_reset;
  wire  line_786_valid;
  reg  line_786_valid_reg;
  wire [39:0] _dataArb_io_in_1_bits_addr_T_1 = {s2_vaddr[39:5], 5'h0}; // @[src/main/scala/rocket/DCache.scala 712:57]
  wire [39:0] _GEN_480 = {{35'd0}, d_address_inc}; // @[src/main/scala/rocket/DCache.scala 712:67]
  wire [39:0] _dataArb_io_in_1_bits_addr_T_2 = _dataArb_io_in_1_bits_addr_T_1 | _GEN_480; // @[src/main/scala/rocket/DCache.scala 712:67]
  wire [3:0] _metaArb_io_in_3_bits_data_T_1 = {s2_write,_c_cat_T_49,auto_out_d_bits_param}; // @[src/main/scala/tilelink/Metadata.scala 84:18]
  wire [1:0] _metaArb_io_in_3_bits_data_T_11 = 4'h1 == _metaArb_io_in_3_bits_data_T_1 ? 2'h1 : 2'h0; // @[src/main/scala/tilelink/Metadata.scala 84:38]
  wire [1:0] _metaArb_io_in_3_bits_data_T_13 = 4'h0 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_11; // @[src/main/scala/tilelink/Metadata.scala 84:38]
  wire [1:0] _metaArb_io_in_3_bits_data_T_15 = 4'h4 == _metaArb_io_in_3_bits_data_T_1 ? 2'h2 :
    _metaArb_io_in_3_bits_data_T_13; // @[src/main/scala/tilelink/Metadata.scala 84:38]
  wire [1:0] metaArb_io_in_3_bits_data_meta_state = 4'hc == _metaArb_io_in_3_bits_data_T_1 ? 2'h3 :
    _metaArb_io_in_3_bits_data_T_15; // @[src/main/scala/tilelink/Metadata.scala 84:38]
  wire  line_787_clock;
  wire  line_787_reset;
  wire  line_787_valid;
  reg  line_787_valid_reg;
  wire  line_788_clock;
  wire  line_788_reset;
  wire  line_788_valid;
  reg  line_788_valid_reg;
  wire  _GEN_355 = auto_out_d_valid ? 1'h0 : _GEN_160; // @[src/main/scala/rocket/DCache.scala 739:29 740:26]
  wire  _GEN_356 = auto_out_d_valid | auto_out_d_valid & grantIsRefill & canAcceptCachedGrant; // @[src/main/scala/rocket/DCache.scala 705:26 739:29 741:32]
  wire  _GEN_357 = auto_out_d_valid ? 1'h0 : 1'h1; // @[src/main/scala/rocket/DCache.scala 739:29 711:33 742:37]
  wire [39:0] _metaArb_io_in_6_bits_addr_T_1 = {io_cpu_req_bits_addr[39:32],auto_out_b_bits_address}; // @[src/main/scala/rocket/DCache.scala 757:36]
  wire [1:0] counter1_1 = counter_1 - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire [1:0] _count_T_1 = ~counter1_1; // @[src/main/scala/tilelink/Edges.scala 234:27]
  wire [1:0] c_count = beats1_1 & _count_T_1; // @[src/main/scala/tilelink/Edges.scala 234:25]
  wire  line_789_clock;
  wire  line_789_reset;
  wire  line_789_valid;
  reg  line_789_valid_reg;
  reg  s1_release_data_valid; // @[src/main/scala/rocket/DCache.scala 785:38]
  wire  releaseRejected = s2_release_data_valid & ~_T_278; // @[src/main/scala/rocket/DCache.scala 787:44]
  wire [2:0] _releaseDataBeat_T = {1'h0,c_count}; // @[src/main/scala/rocket/DCache.scala 788:28]
  wire [1:0] _releaseDataBeat_T_1 = {1'h0,s2_release_data_valid}; // @[src/main/scala/rocket/DCache.scala 788:98]
  wire [1:0] _GEN_481 = {{1'd0}, s1_release_data_valid}; // @[src/main/scala/rocket/DCache.scala 788:93]
  wire [1:0] _releaseDataBeat_T_3 = _GEN_481 + _releaseDataBeat_T_1; // @[src/main/scala/rocket/DCache.scala 788:93]
  wire [1:0] _releaseDataBeat_T_4 = releaseRejected ? 2'h0 : _releaseDataBeat_T_3; // @[src/main/scala/rocket/DCache.scala 788:48]
  wire [2:0] _GEN_482 = {{1'd0}, _releaseDataBeat_T_4}; // @[src/main/scala/rocket/DCache.scala 788:43]
  wire [2:0] releaseDataBeat = _releaseDataBeat_T + _GEN_482; // @[src/main/scala/rocket/DCache.scala 788:43]
  wire  line_790_clock;
  wire  line_790_reset;
  wire  line_790_valid;
  reg  line_790_valid_reg;
  wire  line_791_clock;
  wire  line_791_reset;
  wire  line_791_valid;
  reg  line_791_valid_reg;
  wire  _T_283 = ~(s2_valid_flush_line | s2_flush_valid_pre_tag_ecc | io_cpu_s2_nack); // @[src/main/scala/rocket/DCache.scala 801:13]
  wire  line_792_clock;
  wire  line_792_reset;
  wire  line_792_valid;
  reg  line_792_valid_reg;
  wire  discard_line = s2_valid_flush_line & s2_req_size[1]; // @[src/main/scala/rocket/DCache.scala 802:46]
  wire [3:0] _release_state_T_14 = s2_victim_dirty & ~discard_line ? 4'h1 : 4'h6; // @[src/main/scala/rocket/DCache.scala 803:27]
  wire [26:0] _probe_bits_T_2 = {s2_victim_tag,s2_req_addr[5]}; // @[src/main/scala/rocket/DCache.scala 806:49]
  wire [31:0] probe_bits_res_address = {_probe_bits_T_2, 5'h0}; // @[src/main/scala/rocket/DCache.scala 806:96]
  wire [3:0] _GEN_365 = s2_want_victimize ? _release_state_T_14 : release_state; // @[src/main/scala/rocket/DCache.scala 800:25 803:21 206:30]
  wire  line_793_clock;
  wire  line_793_reset;
  wire  line_793_valid;
  reg  line_793_valid_reg;
  wire  line_794_clock;
  wire  line_794_reset;
  wire  line_794_valid;
  reg  line_794_valid_reg;
  wire  line_795_clock;
  wire  line_795_reset;
  wire  line_795_valid;
  reg  line_795_valid_reg;
  wire  line_796_clock;
  wire  line_796_reset;
  wire  line_796_valid;
  reg  line_796_valid_reg;
  wire [3:0] _release_state_T_15 = releaseDone ? 4'h7 : 4'h3; // @[src/main/scala/rocket/DCache.scala 817:29]
  wire  line_797_clock;
  wire  line_797_reset;
  wire  line_797_valid;
  reg  line_797_valid_reg;
  wire [3:0] _release_state_T_16 = releaseDone ? 4'h0 : 4'h5; // @[src/main/scala/rocket/DCache.scala 821:29]
  wire [2:0] _GEN_376 = _T_284 ? s2_report_param : 3'h5; // @[src/main/scala/rocket/DCache.scala 795:17 814:45 816:23]
  wire [3:0] _GEN_382 = _T_284 ? _release_state_T_15 : _release_state_T_16; // @[src/main/scala/rocket/DCache.scala 814:45 817:23 821:23]
  wire [3:0] _GEN_384 = s2_prb_ack_data ? 4'h2 : _GEN_382; // @[src/main/scala/rocket/DCache.scala 812:36 813:23]
  wire [2:0] _GEN_387 = s2_prb_ack_data ? 3'h5 : _GEN_376; // @[src/main/scala/rocket/DCache.scala 795:17 812:36]
  wire  line_798_clock;
  wire  line_798_reset;
  wire  line_798_valid;
  reg  line_798_valid_reg;
  wire [3:0] _GEN_405 = s2_probe ? _GEN_384 : _GEN_365; // @[src/main/scala/rocket/DCache.scala 808:21]
  wire [2:0] _GEN_408 = s2_probe ? _GEN_387 : 3'h5; // @[src/main/scala/rocket/DCache.scala 795:17 808:21]
  wire  _T_285 = release_state == 4'h4; // @[src/main/scala/rocket/DCache.scala 825:25]
  wire  line_799_clock;
  wire  line_799_reset;
  wire  line_799_valid;
  reg  line_799_valid_reg;
  wire [39:0] _metaArb_io_in_6_bits_addr_T_3 = {io_cpu_req_bits_addr[39:32],probe_bits_address}; // @[src/main/scala/rocket/DCache.scala 828:40]
  wire  line_800_clock;
  wire  line_800_reset;
  wire  line_800_valid;
  reg  line_800_valid_reg;
  wire [3:0] _GEN_415 = metaArb_io_in_6_ready ? 4'h0 : _GEN_405; // @[src/main/scala/rocket/DCache.scala 829:37 830:23]
  wire  _GEN_416 = metaArb_io_in_6_ready | _s1_probe_T; // @[src/main/scala/rocket/DCache.scala 829:37 831:18 161:25]
  wire [3:0] _GEN_420 = release_state == 4'h4 ? _GEN_415 : _GEN_405; // @[src/main/scala/rocket/DCache.scala 825:44]
  wire  line_801_clock;
  wire  line_801_reset;
  wire  line_801_valid;
  reg  line_801_valid_reg;
  wire  line_802_clock;
  wire  line_802_reset;
  wire  line_802_valid;
  reg  line_802_valid_reg;
  wire [3:0] _GEN_422 = releaseDone ? 4'h0 : _GEN_420; // @[src/main/scala/rocket/DCache.scala 836:{26,42}]
  wire [3:0] _GEN_424 = release_state == 4'h5 ? _GEN_422 : _GEN_420; // @[src/main/scala/rocket/DCache.scala 834:47]
  wire  line_803_clock;
  wire  line_803_reset;
  wire  line_803_valid;
  reg  line_803_valid_reg;
  wire  line_804_clock;
  wire  line_804_reset;
  wire  line_804_valid;
  reg  line_804_valid_reg;
  wire [3:0] _GEN_425 = releaseDone ? 4'h7 : _GEN_424; // @[src/main/scala/rocket/DCache.scala 841:{26,42}]
  wire [2:0] _GEN_428 = release_state == 4'h3 ? s2_report_param : _GEN_408; // @[src/main/scala/rocket/DCache.scala 838:48 840:21]
  wire [3:0] _GEN_434 = release_state == 4'h3 ? _GEN_425 : _GEN_424; // @[src/main/scala/rocket/DCache.scala 838:48]
  wire  line_805_clock;
  wire  line_805_reset;
  wire  line_805_valid;
  reg  line_805_valid_reg;
  wire  line_806_clock;
  wire  line_806_reset;
  wire  line_806_valid;
  reg  line_806_valid_reg;
  wire [3:0] _GEN_435 = releaseDone ? 4'h7 : _GEN_434; // @[src/main/scala/rocket/DCache.scala 845:{26,42}]
  wire [2:0] _GEN_437 = release_state == 4'h2 ? s2_report_param : _GEN_428; // @[src/main/scala/rocket/DCache.scala 843:48 844:21]
  wire [3:0] _GEN_443 = release_state == 4'h2 ? _GEN_435 : _GEN_434; // @[src/main/scala/rocket/DCache.scala 843:48]
  wire  line_807_clock;
  wire  line_807_reset;
  wire  line_807_valid;
  reg  line_807_valid_reg;
  wire  line_808_clock;
  wire  line_808_reset;
  wire  line_808_valid;
  reg  line_808_valid_reg;
  wire  line_809_clock;
  wire  line_809_reset;
  wire  line_809_valid;
  reg  line_809_valid_reg;
  wire  line_810_clock;
  wire  line_810_reset;
  wire  line_810_valid;
  reg  line_810_valid_reg;
  wire  _T_296 = _T_278 & c_first; // @[src/main/scala/rocket/DCache.scala 863:27]
  wire  line_811_clock;
  wire  line_811_reset;
  wire  line_811_valid;
  reg  line_811_valid_reg;
  wire  _GEN_452 = _T_278 & c_first | _GEN_352; // @[src/main/scala/rocket/DCache.scala 863:39 864:26]
  wire [1:0] newCoh_state = _T_293 ? voluntaryNewCoh_state : probeNewCoh_state; // @[src/main/scala/rocket/DCache.scala 847:102 860:14 796:27]
  wire [5:0] _dataArb_io_in_2_bits_addr_T_1 = {probe_bits_address[5], 5'h0}; // @[src/main/scala/rocket/DCache.scala 887:55]
  wire [4:0] _dataArb_io_in_2_bits_addr_T_3 = {releaseDataBeat[1:0], 3'h0}; // @[src/main/scala/rocket/DCache.scala 887:117]
  wire [5:0] _GEN_485 = {{1'd0}, _dataArb_io_in_2_bits_addr_T_3}; // @[src/main/scala/rocket/DCache.scala 887:72]
  wire  _metaArb_io_in_4_valid_T_1 = release_state == 4'h7; // @[src/main/scala/util/package.scala 16:47]
  wire [25:0] metaArb_io_in_4_bits_data_meta_tag = probe_bits_address[31:6]; // @[src/main/scala/rocket/DCache.scala 897:78]
  wire  _T_297 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_812_clock;
  wire  line_812_reset;
  wire  line_812_valid;
  reg  line_812_valid_reg;
  reg  io_cpu_s2_xcpt_REG; // @[src/main/scala/rocket/DCache.scala 916:32]
  wire  line_813_clock;
  wire  line_813_reset;
  wire  line_813_valid;
  reg  line_813_valid_reg;
  reg  doUncachedResp; // @[src/main/scala/rocket/DCache.scala 931:31]
  wire  line_814_clock;
  wire  line_814_reset;
  wire  line_814_valid;
  reg  line_814_valid_reg;
  wire  line_815_clock;
  wire  line_815_reset;
  wire  line_815_valid;
  reg  line_815_valid_reg;
  wire  _T_303 = ~_io_cpu_s2_nack_T_4; // @[src/main/scala/rocket/DCache.scala 935:11]
  wire  line_816_clock;
  wire  line_816_reset;
  wire  line_816_valid;
  reg  line_816_valid_reg;
  wire [31:0] io_cpu_resp_bits_data_shifted = get_a_mask_bit ? s2_data_corrected[63:32] : s2_data_corrected[31:0]; // @[src/main/scala/rocket/AMOALU.scala 41:24]
  wire [31:0] _io_cpu_resp_bits_data_T_4 = s2_req_signed & io_cpu_resp_bits_data_shifted[31] ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/AMOALU.scala 44:49]
  wire [31:0] _io_cpu_resp_bits_data_T_6 = s2_req_size == 2'h2 ? _io_cpu_resp_bits_data_T_4 : s2_data_corrected[63:32]; // @[src/main/scala/rocket/AMOALU.scala 44:20]
  wire [63:0] _io_cpu_resp_bits_data_T_7 = {_io_cpu_resp_bits_data_T_6,io_cpu_resp_bits_data_shifted}; // @[src/main/scala/rocket/AMOALU.scala 44:16]
  wire [15:0] io_cpu_resp_bits_data_shifted_1 = get_a_mask_bit_1 ? _io_cpu_resp_bits_data_T_7[31:16] :
    _io_cpu_resp_bits_data_T_7[15:0]; // @[src/main/scala/rocket/AMOALU.scala 41:24]
  wire [47:0] _io_cpu_resp_bits_data_T_12 = s2_req_signed & io_cpu_resp_bits_data_shifted_1[15] ? 48'hffffffffffff : 48'h0
    ; // @[src/main/scala/rocket/AMOALU.scala 44:49]
  wire [47:0] _io_cpu_resp_bits_data_T_14 = s2_req_size == 2'h1 ? _io_cpu_resp_bits_data_T_12 :
    _io_cpu_resp_bits_data_T_7[63:16]; // @[src/main/scala/rocket/AMOALU.scala 44:20]
  wire [63:0] _io_cpu_resp_bits_data_T_15 = {_io_cpu_resp_bits_data_T_14,io_cpu_resp_bits_data_shifted_1}; // @[src/main/scala/rocket/AMOALU.scala 44:16]
  wire [7:0] io_cpu_resp_bits_data_shifted_2 = get_a_mask_bit_2 ? _io_cpu_resp_bits_data_T_15[15:8] :
    _io_cpu_resp_bits_data_T_15[7:0]; // @[src/main/scala/rocket/AMOALU.scala 41:24]
  wire [7:0] io_cpu_resp_bits_data_zeroed_2 = _s2_write_T_3 ? 8'h0 : io_cpu_resp_bits_data_shifted_2; // @[src/main/scala/rocket/AMOALU.scala 43:23]
  wire [55:0] _io_cpu_resp_bits_data_T_20 = s2_req_signed & io_cpu_resp_bits_data_zeroed_2[7] ? 56'hffffffffffffff : 56'h0
    ; // @[src/main/scala/rocket/AMOALU.scala 44:49]
  wire [55:0] _io_cpu_resp_bits_data_T_22 = s2_req_size == 2'h0 | _s2_write_T_3 ? _io_cpu_resp_bits_data_T_20 :
    _io_cpu_resp_bits_data_T_15[63:8]; // @[src/main/scala/rocket/AMOALU.scala 44:20]
  wire [63:0] _io_cpu_resp_bits_data_T_23 = {_io_cpu_resp_bits_data_T_22,io_cpu_resp_bits_data_zeroed_2}; // @[src/main/scala/rocket/AMOALU.scala 44:16]
  wire [63:0] _GEN_486 = {{63'd0}, s2_sc_fail}; // @[src/main/scala/rocket/DCache.scala 957:41]
  wire [6:0] _mask_T = 7'h1 << io_cpu_resp_bits_size; // @[src/main/scala/rocket/DCache.scala 970:36]
  wire [135:0] _mask_T_1 = 136'h1 << _mask_T; // @[src/main/scala/rocket/DCache.scala 970:23]
  wire [135:0] _mask_T_3 = _mask_T_1 - 136'h1; // @[src/main/scala/rocket/DCache.scala 970:56]
  wire [7:0] mask = _mask_T_3[7:0]; // @[src/main/scala/rocket/DCache.scala 969:20 970:10]
  wire [7:0] _masked_data_T_8 = mask[0] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_9 = mask[1] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_10 = mask[2] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_11 = mask[3] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_12 = mask[4] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_13 = mask[5] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_14 = mask[6] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [7:0] _masked_data_T_15 = mask[7] ? 8'hff : 8'h0; // @[src/main/scala/rocket/DCache.scala 971:38]
  wire [63:0] _masked_data_T_16 = {_masked_data_T_15,_masked_data_T_14,_masked_data_T_13,_masked_data_T_12,
    _masked_data_T_11,_masked_data_T_10,_masked_data_T_9,_masked_data_T_8}; // @[src/main/scala/rocket/DCache.scala 971:38]
  reg  REG; // @[src/main/scala/rocket/DCache.scala 1005:18]
  wire  line_817_clock;
  wire  line_817_reset;
  wire  line_817_valid;
  reg  line_817_valid_reg;
  wire  _GEN_470 = REG | resetting; // @[src/main/scala/rocket/DCache.scala 1005:{34,46} 202:26]
  wire [1:0] flushCounterNext = flushCounter + 1'h1; // @[src/main/scala/rocket/DCache.scala 1006:39]
  wire  flushDone = flushCounterNext[1]; // @[src/main/scala/rocket/DCache.scala 1007:37]
  wire  _s1_flush_valid_T = metaArb_io_in_5_ready & metaArb_io_in_5_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [5:0] _metaArb_io_in_5_bits_addr_T_1 = {metaArb_io_in_5_bits_idx, 5'h0}; // @[src/main/scala/rocket/DCache.scala 1015:98]
  wire  line_818_clock;
  wire  line_818_reset;
  wire  line_818_valid;
  reg  line_818_valid_reg;
  wire  line_819_clock;
  wire  line_819_reset;
  wire  line_819_valid;
  reg  line_819_valid_reg;
  wire [1:0] _GEN_472 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[src/main/scala/rocket/DCache.scala 1048:20 1049:18 203:29]
  wire  line_820_clock;
  wire  line_820_reset;
  wire  line_820_valid;
  reg  line_820_valid_reg;
  reg [1:0] io_cpu_perf_release_counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] io_cpu_perf_release_counter1 = io_cpu_perf_release_counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  io_cpu_perf_release_first = io_cpu_perf_release_counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  io_cpu_perf_release_last = io_cpu_perf_release_counter == 2'h1 | beats1_1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  line_821_clock;
  wire  line_821_reset;
  wire  line_821_valid;
  reg  line_821_valid_reg;
  wire  _io_cpu_perf_blocked_near_end_of_refill_T_1 = _T_252 & grantIsRefill; // @[src/main/scala/rocket/DCache.scala 1100:27]
  wire  line_822_clock;
  wire  line_822_reset;
  wire  line_822_valid;
  reg  line_822_valid_reg;
  wire  _T_313 = ~grantIsCached; // @[src/main/scala/rocket/DCache.scala 1130:35]
  wire [1:0] _GEN_489 = reset ? 2'h0 : _GEN_472; // @[src/main/scala/rocket/DCache.scala 203:{29,29}]
  wire  _GEN_494 = _T_252 & _T_313; // @[src/main/scala/rocket/DCache.scala 671:17]
  TLB tlb ( // @[src/main/scala/rocket/DCache.scala 114:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_req_bits_prv(tlb_io_req_bits_prv),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_req_bits_bits_need_gpa(tlb_io_ptw_req_bits_bits_need_gpa),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_ptw(tlb_io_ptw_resp_bits_ae_ptw),
    .io_ptw_resp_bits_ae_final(tlb_io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pf(tlb_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum)
  );
  DCacheModuleImpl_Anon pma_checker ( // @[src/main/scala/rocket/DCache.scala 115:27]
    .clock(pma_checker_clock),
    .reset(pma_checker_reset),
    .io_req_bits_vaddr(pma_checker_io_req_bits_vaddr)
  );
  MaxPeriodFibonacciLFSR lfsr_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(lfsr_prng_clock),
    .reset(lfsr_prng_reset),
    .io_increment(lfsr_prng_io_increment)
  );
  DCacheModuleImpl_Anon_1 metaArb ( // @[src/main/scala/rocket/DCache.scala 119:23]
    .clock(metaArb_clock),
    .reset(metaArb_reset),
    .io_in_0_valid(metaArb_io_in_0_valid),
    .io_in_0_bits_addr(metaArb_io_in_0_bits_addr),
    .io_in_0_bits_idx(metaArb_io_in_0_bits_idx),
    .io_in_2_valid(metaArb_io_in_2_valid),
    .io_in_2_bits_addr(metaArb_io_in_2_bits_addr),
    .io_in_2_bits_idx(metaArb_io_in_2_bits_idx),
    .io_in_2_bits_data(metaArb_io_in_2_bits_data),
    .io_in_3_valid(metaArb_io_in_3_valid),
    .io_in_3_bits_addr(metaArb_io_in_3_bits_addr),
    .io_in_3_bits_idx(metaArb_io_in_3_bits_idx),
    .io_in_3_bits_data(metaArb_io_in_3_bits_data),
    .io_in_4_ready(metaArb_io_in_4_ready),
    .io_in_4_valid(metaArb_io_in_4_valid),
    .io_in_4_bits_addr(metaArb_io_in_4_bits_addr),
    .io_in_4_bits_idx(metaArb_io_in_4_bits_idx),
    .io_in_4_bits_data(metaArb_io_in_4_bits_data),
    .io_in_5_ready(metaArb_io_in_5_ready),
    .io_in_5_valid(metaArb_io_in_5_valid),
    .io_in_5_bits_addr(metaArb_io_in_5_bits_addr),
    .io_in_5_bits_idx(metaArb_io_in_5_bits_idx),
    .io_in_6_ready(metaArb_io_in_6_ready),
    .io_in_6_valid(metaArb_io_in_6_valid),
    .io_in_6_bits_addr(metaArb_io_in_6_bits_addr),
    .io_in_6_bits_idx(metaArb_io_in_6_bits_idx),
    .io_in_6_bits_data(metaArb_io_in_6_bits_data),
    .io_in_7_ready(metaArb_io_in_7_ready),
    .io_in_7_valid(metaArb_io_in_7_valid),
    .io_in_7_bits_addr(metaArb_io_in_7_bits_addr),
    .io_in_7_bits_idx(metaArb_io_in_7_bits_idx),
    .io_in_7_bits_data(metaArb_io_in_7_bits_data),
    .io_out_valid(metaArb_io_out_valid),
    .io_out_bits_write(metaArb_io_out_bits_write),
    .io_out_bits_addr(metaArb_io_out_bits_addr),
    .io_out_bits_idx(metaArb_io_out_bits_idx),
    .io_out_bits_data(metaArb_io_out_bits_data)
  );
  DCacheDataArray data ( // @[src/main/scala/rocket/DCache.scala 129:20]
    .clock(data_clock),
    .reset(data_reset),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_resp_0(data_io_resp_0)
  );
  DCacheModuleImpl_Anon_2 dataArb ( // @[src/main/scala/rocket/DCache.scala 130:23]
    .clock(dataArb_clock),
    .reset(dataArb_reset),
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_wordMask(dataArb_io_in_3_bits_wordMask),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_eccMask(dataArb_io_out_bits_eccMask)
  );
  DelayReg difftest_delayer ( // @[difftest/src/main/scala/util/Delayer.scala 54:15]
    .clock(difftest_delayer_clock),
    .reset(difftest_delayer_reset),
    .i_valid(difftest_delayer_i_valid),
    .i_success(difftest_delayer_i_success),
    .o_valid(difftest_delayer_o_valid),
    .o_success(difftest_delayer_o_success)
  );
  DummyDPICWrapper difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_success(difftest_module_io_bits_success)
  );
  DelayReg_1 difftest_delayer_1 ( // @[difftest/src/main/scala/util/Delayer.scala 54:15]
    .clock(difftest_delayer_1_clock),
    .reset(difftest_delayer_1_reset),
    .i_valid(difftest_delayer_1_i_valid),
    .i_addr(difftest_delayer_1_i_addr),
    .i_data(difftest_delayer_1_i_data),
    .i_mask(difftest_delayer_1_i_mask),
    .o_valid(difftest_delayer_1_o_valid),
    .o_addr(difftest_delayer_1_o_addr),
    .o_data(difftest_delayer_1_o_data),
    .o_mask(difftest_delayer_1_o_mask)
  );
  DummyDPICWrapper_1 difftest_module_1 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_1_clock),
    .reset(difftest_module_1_reset),
    .io_valid(difftest_module_1_io_valid),
    .io_bits_valid(difftest_module_1_io_bits_valid),
    .io_bits_addr(difftest_module_1_io_bits_addr),
    .io_bits_data(difftest_module_1_io_bits_data),
    .io_bits_mask(difftest_module_1_io_bits_mask)
  );
  AMOALU amoalus_0 ( // @[src/main/scala/rocket/DCache.scala 979:26]
    .clock(amoalus_0_clock),
    .reset(amoalus_0_reset),
    .io_mask(amoalus_0_io_mask),
    .io_cmd(amoalus_0_io_cmd),
    .io_lhs(amoalus_0_io_lhs),
    .io_rhs(amoalus_0_io_rhs),
    .io_out(amoalus_0_io_out)
  );
  GEN_w1_line #(.COVER_INDEX(706)) line_706 (
    .clock(line_706_clock),
    .reset(line_706_reset),
    .valid(line_706_valid)
  );
  GEN_w1_line #(.COVER_INDEX(707)) line_707 (
    .clock(line_707_clock),
    .reset(line_707_reset),
    .valid(line_707_valid)
  );
  GEN_w1_line #(.COVER_INDEX(708)) line_708 (
    .clock(line_708_clock),
    .reset(line_708_reset),
    .valid(line_708_valid)
  );
  GEN_w1_line #(.COVER_INDEX(709)) line_709 (
    .clock(line_709_clock),
    .reset(line_709_reset),
    .valid(line_709_valid)
  );
  GEN_w1_line #(.COVER_INDEX(710)) line_710 (
    .clock(line_710_clock),
    .reset(line_710_reset),
    .valid(line_710_valid)
  );
  GEN_w1_line #(.COVER_INDEX(711)) line_711 (
    .clock(line_711_clock),
    .reset(line_711_reset),
    .valid(line_711_valid)
  );
  GEN_w1_line #(.COVER_INDEX(712)) line_712 (
    .clock(line_712_clock),
    .reset(line_712_reset),
    .valid(line_712_valid)
  );
  GEN_w1_line #(.COVER_INDEX(713)) line_713 (
    .clock(line_713_clock),
    .reset(line_713_reset),
    .valid(line_713_valid)
  );
  GEN_w1_line #(.COVER_INDEX(714)) line_714 (
    .clock(line_714_clock),
    .reset(line_714_reset),
    .valid(line_714_valid)
  );
  GEN_w1_line #(.COVER_INDEX(715)) line_715 (
    .clock(line_715_clock),
    .reset(line_715_reset),
    .valid(line_715_valid)
  );
  GEN_w1_line #(.COVER_INDEX(716)) line_716 (
    .clock(line_716_clock),
    .reset(line_716_reset),
    .valid(line_716_valid)
  );
  GEN_w1_line #(.COVER_INDEX(717)) line_717 (
    .clock(line_717_clock),
    .reset(line_717_reset),
    .valid(line_717_valid)
  );
  GEN_w1_line #(.COVER_INDEX(718)) line_718 (
    .clock(line_718_clock),
    .reset(line_718_reset),
    .valid(line_718_valid)
  );
  GEN_w1_line #(.COVER_INDEX(719)) line_719 (
    .clock(line_719_clock),
    .reset(line_719_reset),
    .valid(line_719_valid)
  );
  GEN_w1_line #(.COVER_INDEX(720)) line_720 (
    .clock(line_720_clock),
    .reset(line_720_reset),
    .valid(line_720_valid)
  );
  GEN_w1_line #(.COVER_INDEX(721)) line_721 (
    .clock(line_721_clock),
    .reset(line_721_reset),
    .valid(line_721_valid)
  );
  GEN_w1_line #(.COVER_INDEX(722)) line_722 (
    .clock(line_722_clock),
    .reset(line_722_reset),
    .valid(line_722_valid)
  );
  GEN_w1_line #(.COVER_INDEX(723)) line_723 (
    .clock(line_723_clock),
    .reset(line_723_reset),
    .valid(line_723_valid)
  );
  GEN_w1_line #(.COVER_INDEX(724)) line_724 (
    .clock(line_724_clock),
    .reset(line_724_reset),
    .valid(line_724_valid)
  );
  GEN_w1_line #(.COVER_INDEX(725)) line_725 (
    .clock(line_725_clock),
    .reset(line_725_reset),
    .valid(line_725_valid)
  );
  GEN_w1_line #(.COVER_INDEX(726)) line_726 (
    .clock(line_726_clock),
    .reset(line_726_reset),
    .valid(line_726_valid)
  );
  GEN_w1_line #(.COVER_INDEX(727)) line_727 (
    .clock(line_727_clock),
    .reset(line_727_reset),
    .valid(line_727_valid)
  );
  GEN_w1_line #(.COVER_INDEX(728)) line_728 (
    .clock(line_728_clock),
    .reset(line_728_reset),
    .valid(line_728_valid)
  );
  GEN_w1_line #(.COVER_INDEX(729)) line_729 (
    .clock(line_729_clock),
    .reset(line_729_reset),
    .valid(line_729_valid)
  );
  GEN_w1_line #(.COVER_INDEX(730)) line_730 (
    .clock(line_730_clock),
    .reset(line_730_reset),
    .valid(line_730_valid)
  );
  GEN_w1_line #(.COVER_INDEX(731)) line_731 (
    .clock(line_731_clock),
    .reset(line_731_reset),
    .valid(line_731_valid)
  );
  GEN_w1_line #(.COVER_INDEX(732)) line_732 (
    .clock(line_732_clock),
    .reset(line_732_reset),
    .valid(line_732_valid)
  );
  GEN_w1_line #(.COVER_INDEX(733)) line_733 (
    .clock(line_733_clock),
    .reset(line_733_reset),
    .valid(line_733_valid)
  );
  GEN_w1_line #(.COVER_INDEX(734)) line_734 (
    .clock(line_734_clock),
    .reset(line_734_reset),
    .valid(line_734_valid)
  );
  GEN_w1_line #(.COVER_INDEX(735)) line_735 (
    .clock(line_735_clock),
    .reset(line_735_reset),
    .valid(line_735_valid)
  );
  GEN_w1_line #(.COVER_INDEX(736)) line_736 (
    .clock(line_736_clock),
    .reset(line_736_reset),
    .valid(line_736_valid)
  );
  GEN_w1_line #(.COVER_INDEX(737)) line_737 (
    .clock(line_737_clock),
    .reset(line_737_reset),
    .valid(line_737_valid)
  );
  GEN_w1_line #(.COVER_INDEX(738)) line_738 (
    .clock(line_738_clock),
    .reset(line_738_reset),
    .valid(line_738_valid)
  );
  GEN_w1_line #(.COVER_INDEX(739)) line_739 (
    .clock(line_739_clock),
    .reset(line_739_reset),
    .valid(line_739_valid)
  );
  GEN_w1_line #(.COVER_INDEX(740)) line_740 (
    .clock(line_740_clock),
    .reset(line_740_reset),
    .valid(line_740_valid)
  );
  GEN_w1_line #(.COVER_INDEX(741)) line_741 (
    .clock(line_741_clock),
    .reset(line_741_reset),
    .valid(line_741_valid)
  );
  GEN_w1_line #(.COVER_INDEX(742)) line_742 (
    .clock(line_742_clock),
    .reset(line_742_reset),
    .valid(line_742_valid)
  );
  GEN_w1_line #(.COVER_INDEX(743)) line_743 (
    .clock(line_743_clock),
    .reset(line_743_reset),
    .valid(line_743_valid)
  );
  GEN_w1_line #(.COVER_INDEX(744)) line_744 (
    .clock(line_744_clock),
    .reset(line_744_reset),
    .valid(line_744_valid)
  );
  GEN_w1_line #(.COVER_INDEX(745)) line_745 (
    .clock(line_745_clock),
    .reset(line_745_reset),
    .valid(line_745_valid)
  );
  GEN_w1_line #(.COVER_INDEX(746)) line_746 (
    .clock(line_746_clock),
    .reset(line_746_reset),
    .valid(line_746_valid)
  );
  GEN_w1_line #(.COVER_INDEX(747)) line_747 (
    .clock(line_747_clock),
    .reset(line_747_reset),
    .valid(line_747_valid)
  );
  GEN_w1_line #(.COVER_INDEX(748)) line_748 (
    .clock(line_748_clock),
    .reset(line_748_reset),
    .valid(line_748_valid)
  );
  GEN_w1_line #(.COVER_INDEX(749)) line_749 (
    .clock(line_749_clock),
    .reset(line_749_reset),
    .valid(line_749_valid)
  );
  GEN_w1_line #(.COVER_INDEX(750)) line_750 (
    .clock(line_750_clock),
    .reset(line_750_reset),
    .valid(line_750_valid)
  );
  GEN_w1_line #(.COVER_INDEX(751)) line_751 (
    .clock(line_751_clock),
    .reset(line_751_reset),
    .valid(line_751_valid)
  );
  GEN_w1_line #(.COVER_INDEX(752)) line_752 (
    .clock(line_752_clock),
    .reset(line_752_reset),
    .valid(line_752_valid)
  );
  GEN_w1_line #(.COVER_INDEX(753)) line_753 (
    .clock(line_753_clock),
    .reset(line_753_reset),
    .valid(line_753_valid)
  );
  GEN_w1_line #(.COVER_INDEX(754)) line_754 (
    .clock(line_754_clock),
    .reset(line_754_reset),
    .valid(line_754_valid)
  );
  GEN_w1_line #(.COVER_INDEX(755)) line_755 (
    .clock(line_755_clock),
    .reset(line_755_reset),
    .valid(line_755_valid)
  );
  GEN_w1_line #(.COVER_INDEX(756)) line_756 (
    .clock(line_756_clock),
    .reset(line_756_reset),
    .valid(line_756_valid)
  );
  GEN_w1_line #(.COVER_INDEX(757)) line_757 (
    .clock(line_757_clock),
    .reset(line_757_reset),
    .valid(line_757_valid)
  );
  GEN_w1_line #(.COVER_INDEX(758)) line_758 (
    .clock(line_758_clock),
    .reset(line_758_reset),
    .valid(line_758_valid)
  );
  GEN_w1_line #(.COVER_INDEX(759)) line_759 (
    .clock(line_759_clock),
    .reset(line_759_reset),
    .valid(line_759_valid)
  );
  GEN_w1_line #(.COVER_INDEX(760)) line_760 (
    .clock(line_760_clock),
    .reset(line_760_reset),
    .valid(line_760_valid)
  );
  GEN_w1_line #(.COVER_INDEX(761)) line_761 (
    .clock(line_761_clock),
    .reset(line_761_reset),
    .valid(line_761_valid)
  );
  GEN_w1_line #(.COVER_INDEX(762)) line_762 (
    .clock(line_762_clock),
    .reset(line_762_reset),
    .valid(line_762_valid)
  );
  GEN_w1_line #(.COVER_INDEX(763)) line_763 (
    .clock(line_763_clock),
    .reset(line_763_reset),
    .valid(line_763_valid)
  );
  GEN_w1_line #(.COVER_INDEX(764)) line_764 (
    .clock(line_764_clock),
    .reset(line_764_reset),
    .valid(line_764_valid)
  );
  GEN_w1_line #(.COVER_INDEX(765)) line_765 (
    .clock(line_765_clock),
    .reset(line_765_reset),
    .valid(line_765_valid)
  );
  GEN_w1_line #(.COVER_INDEX(766)) line_766 (
    .clock(line_766_clock),
    .reset(line_766_reset),
    .valid(line_766_valid)
  );
  GEN_w1_line #(.COVER_INDEX(767)) line_767 (
    .clock(line_767_clock),
    .reset(line_767_reset),
    .valid(line_767_valid)
  );
  GEN_w1_line #(.COVER_INDEX(768)) line_768 (
    .clock(line_768_clock),
    .reset(line_768_reset),
    .valid(line_768_valid)
  );
  GEN_w1_line #(.COVER_INDEX(769)) line_769 (
    .clock(line_769_clock),
    .reset(line_769_reset),
    .valid(line_769_valid)
  );
  GEN_w1_line #(.COVER_INDEX(770)) line_770 (
    .clock(line_770_clock),
    .reset(line_770_reset),
    .valid(line_770_valid)
  );
  GEN_w1_line #(.COVER_INDEX(771)) line_771 (
    .clock(line_771_clock),
    .reset(line_771_reset),
    .valid(line_771_valid)
  );
  GEN_w1_line #(.COVER_INDEX(772)) line_772 (
    .clock(line_772_clock),
    .reset(line_772_reset),
    .valid(line_772_valid)
  );
  GEN_w1_line #(.COVER_INDEX(773)) line_773 (
    .clock(line_773_clock),
    .reset(line_773_reset),
    .valid(line_773_valid)
  );
  GEN_w1_line #(.COVER_INDEX(774)) line_774 (
    .clock(line_774_clock),
    .reset(line_774_reset),
    .valid(line_774_valid)
  );
  GEN_w1_line #(.COVER_INDEX(775)) line_775 (
    .clock(line_775_clock),
    .reset(line_775_reset),
    .valid(line_775_valid)
  );
  GEN_w1_line #(.COVER_INDEX(776)) line_776 (
    .clock(line_776_clock),
    .reset(line_776_reset),
    .valid(line_776_valid)
  );
  GEN_w1_line #(.COVER_INDEX(777)) line_777 (
    .clock(line_777_clock),
    .reset(line_777_reset),
    .valid(line_777_valid)
  );
  GEN_w1_line #(.COVER_INDEX(778)) line_778 (
    .clock(line_778_clock),
    .reset(line_778_reset),
    .valid(line_778_valid)
  );
  GEN_w1_line #(.COVER_INDEX(779)) line_779 (
    .clock(line_779_clock),
    .reset(line_779_reset),
    .valid(line_779_valid)
  );
  GEN_w1_line #(.COVER_INDEX(780)) line_780 (
    .clock(line_780_clock),
    .reset(line_780_reset),
    .valid(line_780_valid)
  );
  GEN_w1_line #(.COVER_INDEX(781)) line_781 (
    .clock(line_781_clock),
    .reset(line_781_reset),
    .valid(line_781_valid)
  );
  GEN_w1_line #(.COVER_INDEX(782)) line_782 (
    .clock(line_782_clock),
    .reset(line_782_reset),
    .valid(line_782_valid)
  );
  GEN_w1_line #(.COVER_INDEX(783)) line_783 (
    .clock(line_783_clock),
    .reset(line_783_reset),
    .valid(line_783_valid)
  );
  GEN_w1_line #(.COVER_INDEX(784)) line_784 (
    .clock(line_784_clock),
    .reset(line_784_reset),
    .valid(line_784_valid)
  );
  GEN_w1_line #(.COVER_INDEX(785)) line_785 (
    .clock(line_785_clock),
    .reset(line_785_reset),
    .valid(line_785_valid)
  );
  GEN_w1_line #(.COVER_INDEX(786)) line_786 (
    .clock(line_786_clock),
    .reset(line_786_reset),
    .valid(line_786_valid)
  );
  GEN_w1_line #(.COVER_INDEX(787)) line_787 (
    .clock(line_787_clock),
    .reset(line_787_reset),
    .valid(line_787_valid)
  );
  GEN_w1_line #(.COVER_INDEX(788)) line_788 (
    .clock(line_788_clock),
    .reset(line_788_reset),
    .valid(line_788_valid)
  );
  GEN_w1_line #(.COVER_INDEX(789)) line_789 (
    .clock(line_789_clock),
    .reset(line_789_reset),
    .valid(line_789_valid)
  );
  GEN_w1_line #(.COVER_INDEX(790)) line_790 (
    .clock(line_790_clock),
    .reset(line_790_reset),
    .valid(line_790_valid)
  );
  GEN_w1_line #(.COVER_INDEX(791)) line_791 (
    .clock(line_791_clock),
    .reset(line_791_reset),
    .valid(line_791_valid)
  );
  GEN_w1_line #(.COVER_INDEX(792)) line_792 (
    .clock(line_792_clock),
    .reset(line_792_reset),
    .valid(line_792_valid)
  );
  GEN_w1_line #(.COVER_INDEX(793)) line_793 (
    .clock(line_793_clock),
    .reset(line_793_reset),
    .valid(line_793_valid)
  );
  GEN_w1_line #(.COVER_INDEX(794)) line_794 (
    .clock(line_794_clock),
    .reset(line_794_reset),
    .valid(line_794_valid)
  );
  GEN_w1_line #(.COVER_INDEX(795)) line_795 (
    .clock(line_795_clock),
    .reset(line_795_reset),
    .valid(line_795_valid)
  );
  GEN_w1_line #(.COVER_INDEX(796)) line_796 (
    .clock(line_796_clock),
    .reset(line_796_reset),
    .valid(line_796_valid)
  );
  GEN_w1_line #(.COVER_INDEX(797)) line_797 (
    .clock(line_797_clock),
    .reset(line_797_reset),
    .valid(line_797_valid)
  );
  GEN_w1_line #(.COVER_INDEX(798)) line_798 (
    .clock(line_798_clock),
    .reset(line_798_reset),
    .valid(line_798_valid)
  );
  GEN_w1_line #(.COVER_INDEX(799)) line_799 (
    .clock(line_799_clock),
    .reset(line_799_reset),
    .valid(line_799_valid)
  );
  GEN_w1_line #(.COVER_INDEX(800)) line_800 (
    .clock(line_800_clock),
    .reset(line_800_reset),
    .valid(line_800_valid)
  );
  GEN_w1_line #(.COVER_INDEX(801)) line_801 (
    .clock(line_801_clock),
    .reset(line_801_reset),
    .valid(line_801_valid)
  );
  GEN_w1_line #(.COVER_INDEX(802)) line_802 (
    .clock(line_802_clock),
    .reset(line_802_reset),
    .valid(line_802_valid)
  );
  GEN_w1_line #(.COVER_INDEX(803)) line_803 (
    .clock(line_803_clock),
    .reset(line_803_reset),
    .valid(line_803_valid)
  );
  GEN_w1_line #(.COVER_INDEX(804)) line_804 (
    .clock(line_804_clock),
    .reset(line_804_reset),
    .valid(line_804_valid)
  );
  GEN_w1_line #(.COVER_INDEX(805)) line_805 (
    .clock(line_805_clock),
    .reset(line_805_reset),
    .valid(line_805_valid)
  );
  GEN_w1_line #(.COVER_INDEX(806)) line_806 (
    .clock(line_806_clock),
    .reset(line_806_reset),
    .valid(line_806_valid)
  );
  GEN_w1_line #(.COVER_INDEX(807)) line_807 (
    .clock(line_807_clock),
    .reset(line_807_reset),
    .valid(line_807_valid)
  );
  GEN_w1_line #(.COVER_INDEX(808)) line_808 (
    .clock(line_808_clock),
    .reset(line_808_reset),
    .valid(line_808_valid)
  );
  GEN_w1_line #(.COVER_INDEX(809)) line_809 (
    .clock(line_809_clock),
    .reset(line_809_reset),
    .valid(line_809_valid)
  );
  GEN_w1_line #(.COVER_INDEX(810)) line_810 (
    .clock(line_810_clock),
    .reset(line_810_reset),
    .valid(line_810_valid)
  );
  GEN_w1_line #(.COVER_INDEX(811)) line_811 (
    .clock(line_811_clock),
    .reset(line_811_reset),
    .valid(line_811_valid)
  );
  GEN_w1_line #(.COVER_INDEX(812)) line_812 (
    .clock(line_812_clock),
    .reset(line_812_reset),
    .valid(line_812_valid)
  );
  GEN_w1_line #(.COVER_INDEX(813)) line_813 (
    .clock(line_813_clock),
    .reset(line_813_reset),
    .valid(line_813_valid)
  );
  GEN_w1_line #(.COVER_INDEX(814)) line_814 (
    .clock(line_814_clock),
    .reset(line_814_reset),
    .valid(line_814_valid)
  );
  GEN_w1_line #(.COVER_INDEX(815)) line_815 (
    .clock(line_815_clock),
    .reset(line_815_reset),
    .valid(line_815_valid)
  );
  GEN_w1_line #(.COVER_INDEX(816)) line_816 (
    .clock(line_816_clock),
    .reset(line_816_reset),
    .valid(line_816_valid)
  );
  GEN_w1_line #(.COVER_INDEX(817)) line_817 (
    .clock(line_817_clock),
    .reset(line_817_reset),
    .valid(line_817_valid)
  );
  GEN_w1_line #(.COVER_INDEX(818)) line_818 (
    .clock(line_818_clock),
    .reset(line_818_reset),
    .valid(line_818_valid)
  );
  GEN_w1_line #(.COVER_INDEX(819)) line_819 (
    .clock(line_819_clock),
    .reset(line_819_reset),
    .valid(line_819_valid)
  );
  GEN_w1_line #(.COVER_INDEX(820)) line_820 (
    .clock(line_820_clock),
    .reset(line_820_reset),
    .valid(line_820_valid)
  );
  GEN_w1_line #(.COVER_INDEX(821)) line_821 (
    .clock(line_821_clock),
    .reset(line_821_reset),
    .valid(line_821_valid)
  );
  GEN_w1_line #(.COVER_INDEX(822)) line_822 (
    .clock(line_822_clock),
    .reset(line_822_reset),
    .valid(line_822_valid)
  );
  assign tag_array_0_s1_meta_en = tag_array_0_s1_meta_en_pipe_0;
  assign tag_array_0_s1_meta_addr = tag_array_0_s1_meta_addr_pipe_0;
  assign tag_array_0_s1_meta_data = tag_array_0[tag_array_0_s1_meta_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign tag_array_0_MPORT_data = metaArb_io_out_bits_data;
  assign tag_array_0_MPORT_addr = metaArb_io_out_bits_idx;
  assign tag_array_0_MPORT_mask = 1'h1;
  assign tag_array_0_MPORT_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign line_706_clock = clock;
  assign line_706_reset = reset;
  assign line_706_valid = _s1_probe_T ^ line_706_valid_reg;
  assign line_707_clock = clock;
  assign line_707_reset = reset;
  assign line_707_valid = _T ^ line_707_valid_reg;
  assign line_708_clock = clock;
  assign line_708_reset = reset;
  assign line_708_valid = s0_clk_en ^ line_708_valid_reg;
  assign line_709_clock = clock;
  assign line_709_reset = reset;
  assign line_709_valid = s0_clk_en ^ line_709_valid_reg;
  assign line_710_clock = clock;
  assign line_710_reset = reset;
  assign line_710_valid = _dataArb_io_in_3_valid_T_56 ^ line_710_valid_reg;
  assign line_711_clock = clock;
  assign line_711_reset = reset;
  assign line_711_valid = _dataArb_io_in_3_valid_T_57 ^ line_711_valid_reg;
  assign line_712_clock = clock;
  assign line_712_reset = reset;
  assign line_712_valid = _T_4 ^ line_712_valid_reg;
  assign line_713_clock = clock;
  assign line_713_reset = reset;
  assign line_713_valid = s0_clk_en ^ line_713_valid_reg;
  assign line_714_clock = clock;
  assign line_714_reset = reset;
  assign line_714_valid = s0_clk_en ^ line_714_valid_reg;
  assign line_715_clock = clock;
  assign line_715_reset = reset;
  assign line_715_valid = _T ^ line_715_valid_reg;
  assign line_716_clock = clock;
  assign line_716_reset = reset;
  assign line_716_valid = _T_10 ^ line_716_valid_reg;
  assign line_717_clock = clock;
  assign line_717_reset = reset;
  assign line_717_valid = _T_14 ^ line_717_valid_reg;
  assign line_718_clock = clock;
  assign line_718_reset = reset;
  assign line_718_valid = _T_19 ^ line_718_valid_reg;
  assign line_719_clock = clock;
  assign line_719_reset = reset;
  assign line_719_valid = s0_clk_en ^ line_719_valid_reg;
  assign line_720_clock = clock;
  assign line_720_reset = reset;
  assign line_720_valid = _dataArb_io_in_3_valid_T_56 ^ line_720_valid_reg;
  assign line_721_clock = clock;
  assign line_721_reset = reset;
  assign line_721_valid = _T_29 ^ line_721_valid_reg;
  assign line_722_clock = clock;
  assign line_722_reset = reset;
  assign line_722_valid = _T_30 ^ line_722_valid_reg;
  assign line_723_clock = clock;
  assign line_723_reset = reset;
  assign line_723_valid = _T_30 ^ line_723_valid_reg;
  assign line_724_clock = clock;
  assign line_724_reset = reset;
  assign line_724_valid = s1_meta_clk_en ^ line_724_valid_reg;
  assign line_725_clock = clock;
  assign line_725_reset = reset;
  assign line_725_valid = s1_meta_clk_en ^ line_725_valid_reg;
  assign line_726_clock = clock;
  assign line_726_reset = reset;
  assign line_726_valid = s1_meta_clk_en ^ line_726_valid_reg;
  assign line_727_clock = clock;
  assign line_727_reset = reset;
  assign line_727_valid = s2_data_en ^ line_727_valid_reg;
  assign line_728_clock = clock;
  assign line_728_reset = reset;
  assign line_728_valid = s1_probe ^ line_728_valid_reg;
  assign line_729_clock = clock;
  assign line_729_reset = reset;
  assign line_729_valid = s1_probe ^ line_729_valid_reg;
  assign line_730_clock = clock;
  assign line_730_reset = reset;
  assign line_730_valid = s1_valid_not_nacked ^ line_730_valid_reg;
  assign line_731_clock = clock;
  assign line_731_reset = reset;
  assign line_731_valid = _T_30 ^ line_731_valid_reg;
  assign line_732_clock = clock;
  assign line_732_reset = reset;
  assign line_732_valid = s1_valid_not_nacked ^ line_732_valid_reg;
  assign line_733_clock = clock;
  assign line_733_reset = reset;
  assign line_733_valid = _T_30 ^ line_733_valid_reg;
  assign line_734_clock = clock;
  assign line_734_reset = reset;
  assign line_734_valid = _T_223 ^ line_734_valid_reg;
  assign line_735_clock = clock;
  assign line_735_reset = reset;
  assign line_735_valid = _T_227 ^ line_735_valid_reg;
  assign line_736_clock = clock;
  assign line_736_reset = reset;
  assign line_736_valid = _lrscBackingOff_T ^ line_736_valid_reg;
  assign line_737_clock = clock;
  assign line_737_reset = reset;
  assign line_737_valid = _T_231 ^ line_737_valid_reg;
  assign line_738_clock = clock;
  assign line_738_reset = reset;
  assign line_738_valid = s1_probe ^ line_738_valid_reg;
  assign line_739_clock = clock;
  assign line_739_reset = reset;
  assign line_739_valid = _pstore1_cmd_T ^ line_739_valid_reg;
  assign line_740_clock = clock;
  assign line_740_reset = reset;
  assign line_740_valid = _pstore1_cmd_T ^ line_740_valid_reg;
  assign line_741_clock = clock;
  assign line_741_reset = reset;
  assign line_741_valid = _pstore1_cmd_T ^ line_741_valid_reg;
  assign line_742_clock = clock;
  assign line_742_reset = reset;
  assign line_742_valid = _pstore1_cmd_T ^ line_742_valid_reg;
  assign line_743_clock = clock;
  assign line_743_reset = reset;
  assign line_743_valid = _pstore1_cmd_T ^ line_743_valid_reg;
  assign line_744_clock = clock;
  assign line_744_reset = reset;
  assign line_744_valid = _pstore1_cmd_T ^ line_744_valid_reg;
  assign line_745_clock = clock;
  assign line_745_reset = reset;
  assign line_745_valid = _dataArb_io_in_3_valid_T_56 ^ line_745_valid_reg;
  assign line_746_clock = clock;
  assign line_746_reset = reset;
  assign line_746_valid = _dataArb_io_in_3_valid_T_57 ^ line_746_valid_reg;
  assign line_747_clock = clock;
  assign line_747_reset = reset;
  assign line_747_valid = _dataArb_io_in_3_valid_T_56 ^ line_747_valid_reg;
  assign line_748_clock = clock;
  assign line_748_reset = reset;
  assign line_748_valid = _T_240 ^ line_748_valid_reg;
  assign line_749_clock = clock;
  assign line_749_reset = reset;
  assign line_749_valid = advance_pstore1 ^ line_749_valid_reg;
  assign line_750_clock = clock;
  assign line_750_reset = reset;
  assign line_750_valid = advance_pstore1 ^ line_750_valid_reg;
  assign line_751_clock = clock;
  assign line_751_reset = reset;
  assign line_751_valid = advance_pstore1 ^ line_751_valid_reg;
  assign line_752_clock = clock;
  assign line_752_reset = reset;
  assign line_752_valid = advance_pstore1 ^ line_752_valid_reg;
  assign line_753_clock = clock;
  assign line_753_reset = reset;
  assign line_753_valid = advance_pstore1 ^ line_753_valid_reg;
  assign line_754_clock = clock;
  assign line_754_reset = reset;
  assign line_754_valid = advance_pstore1 ^ line_754_valid_reg;
  assign line_755_clock = clock;
  assign line_755_reset = reset;
  assign line_755_valid = advance_pstore1 ^ line_755_valid_reg;
  assign line_756_clock = clock;
  assign line_756_reset = reset;
  assign line_756_valid = advance_pstore1 ^ line_756_valid_reg;
  assign line_757_clock = clock;
  assign line_757_reset = reset;
  assign line_757_valid = advance_pstore1 ^ line_757_valid_reg;
  assign line_758_clock = clock;
  assign line_758_reset = reset;
  assign line_758_valid = advance_pstore1 ^ line_758_valid_reg;
  assign line_759_clock = clock;
  assign line_759_reset = reset;
  assign line_759_valid = advance_pstore1 ^ line_759_valid_reg;
  assign line_760_clock = clock;
  assign line_760_reset = reset;
  assign line_760_valid = _T_243 ^ line_760_valid_reg;
  assign line_761_clock = clock;
  assign line_761_reset = reset;
  assign line_761_valid = _dataArb_io_in_3_valid_T_56 ^ line_761_valid_reg;
  assign line_762_clock = clock;
  assign line_762_reset = reset;
  assign line_762_valid = _atomics_T_6 ^ line_762_valid_reg;
  assign line_763_clock = clock;
  assign line_763_reset = reset;
  assign line_763_valid = _T_244 ^ line_763_valid_reg;
  assign line_764_clock = clock;
  assign line_764_reset = reset;
  assign line_764_valid = s2_uncached ^ line_764_valid_reg;
  assign line_765_clock = clock;
  assign line_765_reset = reset;
  assign line_765_valid = a_sel ^ line_765_valid_reg;
  assign line_766_clock = clock;
  assign line_766_reset = reset;
  assign line_766_valid = s2_uncached ^ line_766_valid_reg;
  assign line_767_clock = clock;
  assign line_767_reset = reset;
  assign line_767_valid = _T_252 ^ line_767_valid_reg;
  assign line_768_clock = clock;
  assign line_768_reset = reset;
  assign line_768_valid = _block_probe_for_core_progress_T ^ line_768_valid_reg;
  assign line_769_clock = clock;
  assign line_769_reset = reset;
  assign line_769_valid = _T_252 ^ line_769_valid_reg;
  assign line_770_clock = clock;
  assign line_770_reset = reset;
  assign line_770_valid = grantIsCached ^ line_770_valid_reg;
  assign line_771_clock = clock;
  assign line_771_reset = reset;
  assign line_771_valid = _dataArb_io_in_3_valid_T_56 ^ line_771_valid_reg;
  assign line_772_clock = clock;
  assign line_772_reset = reset;
  assign line_772_valid = _io_cpu_req_ready_T_1 ^ line_772_valid_reg;
  assign line_773_clock = clock;
  assign line_773_reset = reset;
  assign line_773_valid = d_last ^ line_773_valid_reg;
  assign line_774_clock = clock;
  assign line_774_reset = reset;
  assign line_774_valid = grantIsCached ^ line_774_valid_reg;
  assign line_775_clock = clock;
  assign line_775_reset = reset;
  assign line_775_valid = grantIsUncached ^ line_775_valid_reg;
  assign line_776_clock = clock;
  assign line_776_reset = reset;
  assign line_776_valid = _T_257 ^ line_776_valid_reg;
  assign line_777_clock = clock;
  assign line_777_reset = reset;
  assign line_777_valid = _dataArb_io_in_3_valid_T_56 ^ line_777_valid_reg;
  assign line_778_clock = clock;
  assign line_778_reset = reset;
  assign line_778_valid = _a_source_T ^ line_778_valid_reg;
  assign line_779_clock = clock;
  assign line_779_reset = reset;
  assign line_779_valid = grantIsUncachedData ^ line_779_valid_reg;
  assign line_780_clock = clock;
  assign line_780_reset = reset;
  assign line_780_valid = grantIsUncached ^ line_780_valid_reg;
  assign line_781_clock = clock;
  assign line_781_reset = reset;
  assign line_781_valid = grantIsVoluntary ^ line_781_valid_reg;
  assign line_782_clock = clock;
  assign line_782_reset = reset;
  assign line_782_valid = _dataArb_io_in_3_valid_T_56 ^ line_782_valid_reg;
  assign line_783_clock = clock;
  assign line_783_reset = reset;
  assign line_783_valid = _tl_out_a_valid_T_7 ^ line_783_valid_reg;
  assign line_784_clock = clock;
  assign line_784_reset = reset;
  assign line_784_valid = _dataArb_io_in_3_valid_T_56 ^ line_784_valid_reg;
  assign line_785_clock = clock;
  assign line_785_reset = reset;
  assign line_785_valid = _T_271 ^ line_785_valid_reg;
  assign line_786_clock = clock;
  assign line_786_reset = reset;
  assign line_786_valid = _T_273 ^ line_786_valid_reg;
  assign line_787_clock = clock;
  assign line_787_reset = reset;
  assign line_787_valid = _T_275 ^ line_787_valid_reg;
  assign line_788_clock = clock;
  assign line_788_reset = reset;
  assign line_788_valid = auto_out_d_valid ^ line_788_valid_reg;
  assign line_789_clock = clock;
  assign line_789_reset = reset;
  assign line_789_valid = _T_278 ^ line_789_valid_reg;
  assign line_790_clock = clock;
  assign line_790_reset = reset;
  assign line_790_valid = s2_want_victimize ^ line_790_valid_reg;
  assign line_791_clock = clock;
  assign line_791_reset = reset;
  assign line_791_valid = _dataArb_io_in_3_valid_T_56 ^ line_791_valid_reg;
  assign line_792_clock = clock;
  assign line_792_reset = reset;
  assign line_792_valid = _T_283 ^ line_792_valid_reg;
  assign line_793_clock = clock;
  assign line_793_reset = reset;
  assign line_793_valid = s2_probe ^ line_793_valid_reg;
  assign line_794_clock = clock;
  assign line_794_reset = reset;
  assign line_794_valid = s2_prb_ack_data ^ line_794_valid_reg;
  assign line_795_clock = clock;
  assign line_795_reset = reset;
  assign line_795_valid = s2_prb_ack_data ^ line_795_valid_reg;
  assign line_796_clock = clock;
  assign line_796_reset = reset;
  assign line_796_valid = _T_284 ^ line_796_valid_reg;
  assign line_797_clock = clock;
  assign line_797_reset = reset;
  assign line_797_valid = _T_284 ^ line_797_valid_reg;
  assign line_798_clock = clock;
  assign line_798_reset = reset;
  assign line_798_valid = probeNack ^ line_798_valid_reg;
  assign line_799_clock = clock;
  assign line_799_reset = reset;
  assign line_799_valid = _T_285 ^ line_799_valid_reg;
  assign line_800_clock = clock;
  assign line_800_reset = reset;
  assign line_800_valid = metaArb_io_in_6_ready ^ line_800_valid_reg;
  assign line_801_clock = clock;
  assign line_801_reset = reset;
  assign line_801_valid = _T_286 ^ line_801_valid_reg;
  assign line_802_clock = clock;
  assign line_802_reset = reset;
  assign line_802_valid = releaseDone ^ line_802_valid_reg;
  assign line_803_clock = clock;
  assign line_803_reset = reset;
  assign line_803_valid = _T_287 ^ line_803_valid_reg;
  assign line_804_clock = clock;
  assign line_804_reset = reset;
  assign line_804_valid = releaseDone ^ line_804_valid_reg;
  assign line_805_clock = clock;
  assign line_805_reset = reset;
  assign line_805_valid = _T_288 ^ line_805_valid_reg;
  assign line_806_clock = clock;
  assign line_806_reset = reset;
  assign line_806_valid = releaseDone ^ line_806_valid_reg;
  assign line_807_clock = clock;
  assign line_807_reset = reset;
  assign line_807_valid = _T_293 ^ line_807_valid_reg;
  assign line_808_clock = clock;
  assign line_808_reset = reset;
  assign line_808_valid = _T_291 ^ line_808_valid_reg;
  assign line_809_clock = clock;
  assign line_809_reset = reset;
  assign line_809_valid = _T_291 ^ line_809_valid_reg;
  assign line_810_clock = clock;
  assign line_810_reset = reset;
  assign line_810_valid = releaseDone ^ line_810_valid_reg;
  assign line_811_clock = clock;
  assign line_811_reset = reset;
  assign line_811_valid = _T_296 ^ line_811_valid_reg;
  assign line_812_clock = clock;
  assign line_812_reset = reset;
  assign line_812_valid = _T_297 ^ line_812_valid_reg;
  assign line_813_clock = clock;
  assign line_813_reset = reset;
  assign line_813_valid = io_cpu_replay_next ^ line_813_valid_reg;
  assign line_814_clock = clock;
  assign line_814_reset = reset;
  assign line_814_valid = doUncachedResp ^ line_814_valid_reg;
  assign line_815_clock = clock;
  assign line_815_reset = reset;
  assign line_815_valid = _dataArb_io_in_3_valid_T_56 ^ line_815_valid_reg;
  assign line_816_clock = clock;
  assign line_816_reset = reset;
  assign line_816_valid = _T_303 ^ line_816_valid_reg;
  assign line_817_clock = clock;
  assign line_817_reset = reset;
  assign line_817_valid = REG ^ line_817_valid_reg;
  assign line_818_clock = clock;
  assign line_818_reset = reset;
  assign line_818_valid = resetting ^ line_818_valid_reg;
  assign line_819_clock = clock;
  assign line_819_reset = reset;
  assign line_819_valid = flushDone ^ line_819_valid_reg;
  assign line_820_clock = clock;
  assign line_820_reset = reset;
  assign line_820_valid = _T_244 ^ line_820_valid_reg;
  assign line_821_clock = clock;
  assign line_821_reset = reset;
  assign line_821_valid = _T_278 ^ line_821_valid_reg;
  assign line_822_clock = clock;
  assign line_822_reset = reset;
  assign line_822_valid = _io_cpu_perf_blocked_near_end_of_refill_T_1 ^ line_822_valid_reg;
  assign auto_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12; // @[src/main/scala/rocket/DCache.scala 588:32]
  assign auto_out_a_bits_opcode = _s2_valid_cached_miss_T ? 3'h6 : _tl_out_a_bits_T_8_opcode; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_param = _s2_valid_cached_miss_T ? tl_out_a_bits_a_param : 3'h0; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_size = _s2_valid_cached_miss_T ? 3'h5 : _tl_out_a_bits_T_8_size; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_source = _s2_valid_cached_miss_T ? 1'h0 : _tl_out_a_bits_T_8_source; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_address = _s2_valid_cached_miss_T ? tl_out_a_bits_a_address : _tl_out_a_bits_T_8_address; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_mask = _s2_valid_cached_miss_T ? 8'hff : _tl_out_a_bits_T_8_mask; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_a_bits_data = _s2_valid_cached_miss_T ? 64'h0 : _tl_out_a_bits_T_8_data; // @[src/main/scala/rocket/DCache.scala 592:23]
  assign auto_out_b_ready = metaArb_io_in_6_ready & ~(block_probe_for_core_progress | block_probe_for_ordering |
    s1_valid | s2_valid); // @[src/main/scala/rocket/DCache.scala 754:44]
  assign auto_out_c_valid = release_state == 4'h3 | _GEN_423; // @[src/main/scala/rocket/DCache.scala 838:48 839:22]
  assign auto_out_c_bits_opcode = _T_293 ? _GEN_444 : _GEN_436; // @[src/main/scala/rocket/DCache.scala 847:102]
  assign auto_out_c_bits_param = _T_293 ? s2_shrink_param : _GEN_437; // @[src/main/scala/rocket/DCache.scala 847:102]
  assign auto_out_c_bits_size = _T_293 ? 3'h5 : probe_bits_size; // @[src/main/scala/rocket/DCache.scala 847:102]
  assign auto_out_c_bits_source = probe_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/rocket/DCache.scala 868:26]
  assign auto_out_c_bits_address = probe_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/rocket/DCache.scala 869:27]
  assign auto_out_c_bits_data = {s2_data_corrected_hi,s2_data_corrected_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign auto_out_d_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? 1'h0 : _GEN_354; // @[src/main/scala/rocket/DCache.scala 736:68 737:22]
  assign auto_out_e_valid = grantIsRefill & ~dataArb_io_in_1_ready ? 1'h0 : auto_out_d_valid & d_first & grantIsCached
     & canAcceptCachedGrant; // @[src/main/scala/rocket/DCache.scala 698:18 706:51 707:20]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign io_cpu_req_ready = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_355 : _GEN_160; // @[src/main/scala/rocket/DCache.scala 736:68]
  assign io_cpu_s2_nack = s2_valid_no_xcpt & ~s2_dont_nack_uncached & ~s2_dont_nack_misc & ~
    s2_valid_hit_pre_data_ecc_and_waw; // @[src/main/scala/rocket/DCache.scala 423:86]
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp; // @[src/main/scala/rocket/DCache.scala 932:51]
  assign io_cpu_resp_bits_addr = doUncachedResp ? s2_uncached_resp_addr : s2_req_addr; // @[src/main/scala/rocket/DCache.scala 934:25 937:27 901:37]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_cmd = s2_req_cmd; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_size = s2_req_size; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_signed = s2_req_signed; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_dprv = s2_req_dprv; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_dv = 1'h0; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_data = _io_cpu_resp_bits_data_T_23 | _GEN_486; // @[src/main/scala/rocket/DCache.scala 957:41]
  assign io_cpu_resp_bits_mask = 8'h0; // @[src/main/scala/rocket/DCache.scala 901:37]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[src/main/scala/rocket/DCache.scala 934:25 903:27 936:29]
  assign io_cpu_resp_bits_has_data = _s2_read_T_6 | _s2_write_T_21; // @[src/main/scala/rocket/Consts.scala 85:68]
  assign io_cpu_resp_bits_data_word_bypass = {_io_cpu_resp_bits_data_T_6,io_cpu_resp_bits_data_shifted}; // @[src/main/scala/rocket/AMOALU.scala 44:16]
  assign io_cpu_resp_bits_data_raw = {s2_data_corrected_hi,s2_data_corrected_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign io_cpu_resp_bits_store_data = pstore1_data; // @[src/main/scala/rocket/DCache.scala 960:31]
  assign io_cpu_replay_next = _T_252 & grantIsUncachedData; // @[src/main/scala/rocket/DCache.scala 933:39]
  assign io_cpu_s2_xcpt_ma_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_ld; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_ma_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_st; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_pf_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_ld; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_pf_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_st; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_gf_ld = 1'h0; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_gf_st = 1'h0; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_ae_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_ld; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_s2_xcpt_ae_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_st; // @[src/main/scala/rocket/DCache.scala 916:24]
  assign io_cpu_ordered = ~(s1_valid | s2_valid | cached_grant_wait | _s2_valid_cached_miss_T_2); // @[src/main/scala/rocket/DCache.scala 913:21]
  assign io_cpu_perf_release = io_cpu_perf_release_last & _T_278; // @[src/main/scala/tilelink/Edges.scala 233:22]
  assign io_cpu_perf_grant = auto_out_d_valid & d_last; // @[src/main/scala/rocket/DCache.scala 1075:39]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign io_ptw_req_bits_bits_need_gpa = tlb_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb; // @[src/main/scala/rocket/DCache.scala 251:71]
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr; // @[src/main/scala/rocket/DCache.scala 252:19]
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough; // @[src/main/scala/rocket/DCache.scala 252:19]
  assign tlb_io_req_bits_size = s1_tlb_req_size; // @[src/main/scala/rocket/DCache.scala 252:19]
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd; // @[src/main/scala/rocket/DCache.scala 252:19]
  assign tlb_io_req_bits_prv = s1_tlb_req_prv; // @[src/main/scala/rocket/DCache.scala 252:19]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[src/main/scala/rocket/DCache.scala 256:54]
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0]; // @[src/main/scala/rocket/DCache.scala 257:40]
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1]; // @[src/main/scala/rocket/DCache.scala 258:40]
  assign tlb_io_sfence_bits_addr = s1_req_addr[38:0]; // @[src/main/scala/rocket/DCache.scala 260:27]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_ae_ptw = io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_ae_final = io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pf = io_ptw_resp_bits_pf; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[src/main/scala/rocket/DCache.scala 249:10]
  assign pma_checker_clock = clock;
  assign pma_checker_reset = reset;
  assign pma_checker_io_req_bits_vaddr = s1_req_addr; // @[src/main/scala/rocket/DCache.scala 270:33]
  assign lfsr_prng_clock = clock;
  assign lfsr_prng_reset = reset;
  assign lfsr_prng_io_increment = _T_252 & _GEN_330; // @[src/main/scala/rocket/DCache.scala 658:24 src/main/scala/util/Replacement.scala 38:11]
  assign metaArb_clock = clock;
  assign metaArb_reset = reset;
  assign metaArb_io_in_0_valid = resetting; // @[src/main/scala/rocket/DCache.scala 1043:26]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[src/main/scala/rocket/DCache.scala 1044:25]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[src/main/scala/rocket/DCache.scala 1044:25]
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[src/main/scala/rocket/DCache.scala 440:63]
  assign metaArb_io_in_2_bits_addr = {io_cpu_req_bits_addr[39:6],s2_vaddr[5:0]}; // @[src/main/scala/rocket/DCache.scala 444:36]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[5]; // @[src/main/scala/rocket/DCache.scala 443:40]
  assign metaArb_io_in_2_bits_data = {s2_grow_param,metaArb_io_in_2_bits_data_meta_tag}; // @[src/main/scala/rocket/DCache.scala 445:97]
  assign metaArb_io_in_3_valid = grantIsCached & d_done & ~auto_out_d_bits_denied; // @[src/main/scala/rocket/DCache.scala 725:53]
  assign metaArb_io_in_3_bits_addr = {io_cpu_req_bits_addr[39:6],s2_vaddr[5:0]}; // @[src/main/scala/rocket/DCache.scala 729:36]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[5]; // @[src/main/scala/rocket/DCache.scala 728:40]
  assign metaArb_io_in_3_bits_data = {metaArb_io_in_3_bits_data_meta_state,metaArb_io_in_2_bits_data_meta_tag}; // @[src/main/scala/rocket/DCache.scala 730:134]
  assign metaArb_io_in_4_valid = _T_290 | _metaArb_io_in_4_valid_T_1; // @[src/main/scala/util/package.scala 73:59]
  assign metaArb_io_in_4_bits_addr = {io_cpu_req_bits_addr[39:6],probe_bits_address[5:0]}; // @[src/main/scala/rocket/DCache.scala 896:36]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[5]; // @[src/main/scala/rocket/DCache.scala 1197:47]
  assign metaArb_io_in_4_bits_data = {newCoh_state,metaArb_io_in_4_bits_data_meta_tag}; // @[src/main/scala/rocket/DCache.scala 897:97]
  assign metaArb_io_in_5_valid = 1'h0; // @[src/main/scala/rocket/DCache.scala 1012:38]
  assign metaArb_io_in_5_bits_addr = {io_cpu_req_bits_addr[39:6],_metaArb_io_in_5_bits_addr_T_1}; // @[src/main/scala/rocket/DCache.scala 1015:36]
  assign metaArb_io_in_5_bits_idx = flushCounter; // @[src/main/scala/rocket/DCache.scala 1014:44]
  assign metaArb_io_in_6_valid = release_state == 4'h4 | auto_out_b_valid & (~block_probe_for_core_progress |
    lrscBackingOff); // @[src/main/scala/rocket/DCache.scala 753:26 825:44 826:30]
  assign metaArb_io_in_6_bits_addr = release_state == 4'h4 ? _metaArb_io_in_6_bits_addr_T_3 :
    _metaArb_io_in_6_bits_addr_T_1; // @[src/main/scala/rocket/DCache.scala 757:30 825:44 828:34]
  assign metaArb_io_in_6_bits_idx = release_state == 4'h4 ? probe_bits_address[5] : auto_out_b_bits_address[5]; // @[src/main/scala/rocket/DCache.scala 756:29 825:44 827:33]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[src/main/scala/rocket/DCache.scala 759:30]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[src/main/scala/rocket/DCache.scala 239:26]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[src/main/scala/rocket/DCache.scala 242:30]
  assign metaArb_io_in_7_bits_idx = dataArb_io_in_3_bits_addr[5]; // @[src/main/scala/rocket/DCache.scala 241:58]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[src/main/scala/rocket/DCache.scala 244:30]
  assign data_clock = clock;
  assign data_reset = reset;
  assign data_io_req_valid = dataArb_io_out_valid; // @[src/main/scala/rocket/DCache.scala 133:21]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[src/main/scala/rocket/DCache.scala 132:20]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[src/main/scala/rocket/DCache.scala 132:20]
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata; // @[src/main/scala/rocket/DCache.scala 132:20]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[src/main/scala/rocket/DCache.scala 132:20]
  assign dataArb_clock = clock;
  assign dataArb_reset = reset;
  assign dataArb_io_in_0_valid = pstore_drain_structural | _pstore_drain_T_10; // @[src/main/scala/rocket/DCache.scala 501:44]
  assign dataArb_io_in_0_bits_addr = _dataArb_io_in_0_bits_addr_T[5:0]; // @[src/main/scala/rocket/DCache.scala 533:30]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _pstore_drain_T_10; // @[src/main/scala/rocket/DCache.scala 501:44]
  assign dataArb_io_in_0_bits_wdata = {dataArb_io_in_0_bits_wdata_hi,dataArb_io_in_0_bits_wdata_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign dataArb_io_in_0_bits_eccMask = {dataArb_io_in_0_bits_eccMask_hi,dataArb_io_in_0_bits_eccMask_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign dataArb_io_in_1_valid = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_356 : auto_out_d_valid &
    grantIsRefill & canAcceptCachedGrant; // @[src/main/scala/rocket/DCache.scala 705:26 736:68]
  assign dataArb_io_in_1_bits_addr = _dataArb_io_in_1_bits_addr_T_2[5:0]; // @[src/main/scala/rocket/DCache.scala 712:32]
  assign dataArb_io_in_1_bits_write = grantIsUncachedData & (blockUncachedGrant | s1_valid) ? _GEN_357 : 1'h1; // @[src/main/scala/rocket/DCache.scala 711:33 736:68]
  assign dataArb_io_in_1_bits_wdata = {tl_d_data_encoded_hi,tl_d_data_encoded_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign dataArb_io_in_2_valid = inWriteback & releaseDataBeat < 3'h4; // @[src/main/scala/rocket/DCache.scala 884:41]
  assign dataArb_io_in_2_bits_addr = _dataArb_io_in_2_bits_addr_T_1 | _GEN_485; // @[src/main/scala/rocket/DCache.scala 887:72]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[src/main/scala/rocket/DCache.scala 885:25]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & dataArb_io_in_3_valid_res; // @[src/main/scala/rocket/DCache.scala 220:46]
  assign dataArb_io_in_3_bits_addr = _dataArb_io_in_3_bits_addr_T_2[5:0]; // @[src/main/scala/rocket/DCache.scala 223:30]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[src/main/scala/rocket/DCache.scala 221:25]
  assign dataArb_io_in_3_bits_wordMask = 1'h1; // @[src/main/scala/rocket/DCache.scala 224:34]
  assign difftest_delayer_clock = clock;
  assign difftest_delayer_reset = reset;
  assign difftest_delayer_i_valid = io_cpu_resp_valid & _s2_write_T_3; // @[src/main/scala/rocket/DCache.scala 466:43]
  assign difftest_delayer_i_success = lrscValid & lrscAddrMatch; // @[src/main/scala/rocket/DCache.scala 467:35]
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 158:15]
  assign difftest_module_io_bits_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_io_bits_success = difftest_delayer_o_success; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_delayer_1_clock = clock;
  assign difftest_delayer_1_reset = reset;
  assign difftest_delayer_1_i_valid = io_cpu_resp_valid & ~io_cpu_resp_bits_has_data; // @[src/main/scala/rocket/DCache.scala 966:35]
  assign difftest_delayer_1_i_addr = {{24'd0}, io_cpu_resp_bits_addr}; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/DCache.scala 968:21]
  assign difftest_delayer_1_i_data = _masked_data_T_16 & io_cpu_resp_bits_store_data; // @[src/main/scala/rocket/DCache.scala 971:48]
  assign difftest_delayer_1_i_mask = _mask_T_3[7:0]; // @[src/main/scala/rocket/DCache.scala 969:20 970:10]
  assign difftest_module_1_clock = clock;
  assign difftest_module_1_reset = reset;
  assign difftest_module_1_io_valid = difftest_delayer_1_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 158:15]
  assign difftest_module_1_io_bits_valid = difftest_delayer_1_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_1_io_bits_addr = difftest_delayer_1_o_addr; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_1_io_bits_data = difftest_delayer_1_o_data; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_1_io_bits_mask = difftest_delayer_1_o_mask; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign amoalus_0_clock = clock;
  assign amoalus_0_reset = reset;
  assign amoalus_0_io_mask = pstore1_mask; // @[src/main/scala/rocket/DCache.scala 980:38]
  assign amoalus_0_io_cmd = pstore1_cmd; // @[src/main/scala/rocket/DCache.scala 981:21]
  assign amoalus_0_io_lhs = {s2_data_corrected_hi,s2_data_corrected_lo}; // @[src/main/scala/util/package.scala 37:27]
  assign amoalus_0_io_rhs = pstore1_data; // @[src/main/scala/rocket/DCache.scala 983:37]
  always @(posedge clock) begin
    if (tag_array_0_MPORT_en & tag_array_0_MPORT_mask) begin
      tag_array_0[tag_array_0_MPORT_addr] <= tag_array_0_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    tag_array_0_s1_meta_en_pipe_0 <= metaArb_io_out_valid & _s0_clk_en_T;
    if (metaArb_io_out_valid & _s0_clk_en_T) begin
      tag_array_0_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 160:25]
      s1_valid <= 1'h0; // @[src/main/scala/rocket/DCache.scala 160:25]
    end else begin
      s1_valid <= _s1_valid_T; // @[src/main/scala/rocket/DCache.scala 160:25]
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 652:42]
      blockProbeAfterGrantCount <= 3'h0; // @[src/main/scala/rocket/DCache.scala 652:42]
    end else if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        if (d_last) begin // @[src/main/scala/rocket/DCache.scala 662:20]
          blockProbeAfterGrantCount <= 3'h7; // @[src/main/scala/rocket/DCache.scala 665:35]
        end else begin
          blockProbeAfterGrantCount <= _GEN_304;
        end
      end else begin
        blockProbeAfterGrantCount <= _GEN_304;
      end
    end else begin
      blockProbeAfterGrantCount <= _GEN_304;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 450:26]
      lrscCount <= 7'h0; // @[src/main/scala/rocket/DCache.scala 450:26]
    end else if (s1_probe) begin // @[src/main/scala/rocket/DCache.scala 462:19]
      lrscCount <= 7'h0; // @[src/main/scala/rocket/DCache.scala 462:31]
    end else if (s2_valid_masked & lrscValid) begin // @[src/main/scala/rocket/DCache.scala 461:43]
      lrscCount <= 7'h3; // @[src/main/scala/rocket/DCache.scala 461:55]
    end else if (_lrscBackingOff_T) begin // @[src/main/scala/rocket/DCache.scala 460:26]
      lrscCount <= _lrscCount_T_2; // @[src/main/scala/rocket/DCache.scala 460:38]
    end else begin
      lrscCount <= _GEN_237;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 161:25]
      s1_probe <= 1'h0; // @[src/main/scala/rocket/DCache.scala 161:25]
    end else if (release_state == 4'h4) begin // @[src/main/scala/rocket/DCache.scala 825:44]
      s1_probe <= _GEN_416;
    end else begin
      s1_probe <= _s1_probe_T; // @[src/main/scala/rocket/DCache.scala 161:25]
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 311:25]
      s2_probe <= 1'h0; // @[src/main/scala/rocket/DCache.scala 311:25]
    end else begin
      s2_probe <= s1_probe; // @[src/main/scala/rocket/DCache.scala 311:25]
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 206:30]
      release_state <= 4'h0; // @[src/main/scala/rocket/DCache.scala 206:30]
    end else if (_T_297) begin // @[src/main/scala/rocket/DCache.scala 898:32]
      release_state <= 4'h0; // @[src/main/scala/rocket/DCache.scala 898:48]
    end else if (_T_293) begin // @[src/main/scala/rocket/DCache.scala 847:102]
      if (releaseDone) begin // @[src/main/scala/rocket/DCache.scala 862:26]
        release_state <= 4'h6; // @[src/main/scala/rocket/DCache.scala 862:42]
      end else begin
        release_state <= _GEN_443;
      end
    end else begin
      release_state <= _GEN_443;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 204:33]
      release_ack_wait <= 1'h0; // @[src/main/scala/rocket/DCache.scala 204:33]
    end else if (_T_293) begin // @[src/main/scala/rocket/DCache.scala 847:102]
      release_ack_wait <= _GEN_452;
    end else if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (!(grantIsCached)) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        release_ack_wait <= _GEN_326;
      end
    end
    if (_T_293) begin // @[src/main/scala/rocket/DCache.scala 847:102]
      if (_T_278 & c_first) begin // @[src/main/scala/rocket/DCache.scala 863:39]
        release_ack_addr <= probe_bits_address; // @[src/main/scala/rocket/DCache.scala 865:26]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 651:32]
      grantInProgress <= 1'h0; // @[src/main/scala/rocket/DCache.scala 651:32]
    end else if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        if (d_last) begin // @[src/main/scala/rocket/DCache.scala 662:20]
          grantInProgress <= 1'h0; // @[src/main/scala/rocket/DCache.scala 664:25]
        end else begin
          grantInProgress <= 1'h1; // @[src/main/scala/rocket/DCache.scala 660:23]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 309:25]
      s2_valid <= 1'h0; // @[src/main/scala/rocket/DCache.scala 309:25]
    end else begin
      s2_valid <= s1_valid_masked & ~s1_sfence; // @[src/main/scala/rocket/DCache.scala 309:25]
    end
    if (s2_want_victimize) begin // @[src/main/scala/rocket/DCache.scala 800:25]
      probe_bits_param <= 2'h0; // @[src/main/scala/rocket/DCache.scala 806:18]
    end else if (_s1_probe_T) begin // @[src/main/scala/rocket/DCache.scala 162:29]
      probe_bits_param <= auto_out_b_bits_param; // @[src/main/scala/rocket/DCache.scala 162:29]
    end
    if (s2_want_victimize) begin // @[src/main/scala/rocket/DCache.scala 800:25]
      probe_bits_size <= 3'h0; // @[src/main/scala/rocket/DCache.scala 806:18]
    end else if (_s1_probe_T) begin // @[src/main/scala/rocket/DCache.scala 162:29]
      probe_bits_size <= auto_out_b_bits_size; // @[src/main/scala/rocket/DCache.scala 162:29]
    end
    if (s2_want_victimize) begin // @[src/main/scala/rocket/DCache.scala 800:25]
      probe_bits_source <= 1'h0; // @[src/main/scala/rocket/DCache.scala 806:18]
    end else if (_s1_probe_T) begin // @[src/main/scala/rocket/DCache.scala 162:29]
      probe_bits_source <= auto_out_b_bits_source; // @[src/main/scala/rocket/DCache.scala 162:29]
    end
    if (s2_want_victimize) begin // @[src/main/scala/rocket/DCache.scala 800:25]
      probe_bits_address <= probe_bits_res_address; // @[src/main/scala/rocket/DCache.scala 806:18]
    end else if (_s1_probe_T) begin // @[src/main/scala/rocket/DCache.scala 162:29]
      probe_bits_address <= auto_out_b_bits_address; // @[src/main/scala/rocket/DCache.scala 162:29]
    end
    line_706_valid_reg <= _s1_probe_T;
    if (s1_probe) begin // @[src/main/scala/rocket/DCache.scala 362:33]
      if (_s1_meta_hit_way_T_1 & ~s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 297:41]
        s2_probe_state_state <= s1_meta_uncorrected_0_coh_state;
      end else begin
        s2_probe_state_state <= 2'h0;
      end
    end
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      counter_1 <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_T_278) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (c_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (beats1_opdata_1) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          counter_1 <= beats1_decode_1;
        end else begin
          counter_1 <= 2'h0;
        end
      end else begin
        counter_1 <= counter1_1;
      end
    end
    s2_release_data_valid <= s1_release_data_valid & ~releaseRejected; // @[src/main/scala/rocket/DCache.scala 786:61]
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_cmd <= io_cpu_req_bits_cmd; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        s2_req_cmd <= _GEN_176;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
          s2_req_cmd <= 5'h0; // @[src/main/scala/rocket/DCache.scala 679:22]
        end else begin
          s2_req_cmd <= _GEN_176;
        end
      end else begin
        s2_req_cmd <= _GEN_176;
      end
    end else begin
      s2_req_cmd <= _GEN_176;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 488:29]
      pstore1_held <= 1'h0; // @[src/main/scala/rocket/DCache.scala 488:29]
    end else begin
      pstore1_held <= pstore1_valid & pstore2_valid & ~pstore_drain; // @[src/main/scala/rocket/DCache.scala 505:16]
    end
    if (_pstore1_cmd_T) begin // @[src/main/scala/rocket/DCache.scala 477:31]
      pstore1_addr <= s1_vaddr; // @[src/main/scala/rocket/DCache.scala 477:31]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_addr <= s0_req_addr; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    if (_pstore1_cmd_T) begin // @[src/main/scala/rocket/DCache.scala 480:31]
      if (_s1_write_T_1) begin // @[src/main/scala/rocket/DCache.scala 305:20]
        pstore1_mask <= io_cpu_s1_data_mask;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_size <= io_cpu_req_bits_size; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 485:30]
      pstore2_valid <= 1'h0; // @[src/main/scala/rocket/DCache.scala 485:30]
    end else begin
      pstore2_valid <= pstore2_valid & _pstore1_held_T_9 | advance_pstore1; // @[src/main/scala/rocket/DCache.scala 507:17]
    end
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 508:31]
      pstore2_addr <= pstore1_addr; // @[src/main/scala/rocket/DCache.scala 508:31]
    end
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 516:45]
      pstore2_storegen_mask <= _pstore2_storegen_mask_mask_T_2; // @[src/main/scala/rocket/DCache.scala 518:12]
    end
    s2_not_nacked_in_s1 <= ~s1_nack; // @[src/main/scala/rocket/DCache.scala 313:37]
    if (_T_30) begin // @[src/main/scala/rocket/DCache.scala 364:31]
      if (_s1_meta_hit_way_T_1 & ~s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 297:41]
        s2_hit_state_state <= s1_meta_uncorrected_0_coh_state;
      end else begin
        s2_hit_state_state <= 2'h0;
      end
    end
    line_707_valid_reg <= _T;
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_tag <= io_cpu_req_bits_tag; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_signed <= io_cpu_req_bits_signed; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 174:25]
      s1_req_dprv <= io_cpu_req_bits_dprv; // @[src/main/scala/rocket/DCache.scala 174:25]
    end
    line_708_valid_reg <= s0_clk_en;
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 186:29]
      s1_tlb_req_vaddr <= s0_req_addr; // @[src/main/scala/rocket/DCache.scala 186:29]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 186:29]
      s1_tlb_req_passthrough <= s0_req_phys; // @[src/main/scala/rocket/DCache.scala 186:29]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 186:29]
      s1_tlb_req_size <= io_cpu_req_bits_size; // @[src/main/scala/rocket/DCache.scala 186:29]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 186:29]
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd; // @[src/main/scala/rocket/DCache.scala 186:29]
    end
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 186:29]
      s1_tlb_req_prv <= io_cpu_req_bits_dprv; // @[src/main/scala/rocket/DCache.scala 186:29]
    end
    line_709_valid_reg <= s0_clk_en;
    s1_flush_valid <= _s1_flush_valid_T & _s1_meta_hit_state_T_1 & _s2_cannot_victimize_T & _io_cpu_req_ready_T &
      _tl_out_a_valid_T_7; // @[src/main/scala/rocket/DCache.scala 1011:122]
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 201:34]
      cached_grant_wait <= 1'h0; // @[src/main/scala/rocket/DCache.scala 201:34]
    end else if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        if (d_last) begin // @[src/main/scala/rocket/DCache.scala 662:20]
          cached_grant_wait <= 1'h0; // @[src/main/scala/rocket/DCache.scala 663:27]
        end else begin
          cached_grant_wait <= _GEN_301;
        end
      end else begin
        cached_grant_wait <= _GEN_301;
      end
    end else begin
      cached_grant_wait <= _GEN_301;
    end
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 202:26]
      resetting <= 1'h0; // @[src/main/scala/rocket/DCache.scala 202:26]
    end else if (resetting) begin // @[src/main/scala/rocket/DCache.scala 1048:20]
      if (flushDone) begin // @[src/main/scala/rocket/DCache.scala 1050:22]
        resetting <= 1'h0; // @[src/main/scala/rocket/DCache.scala 1051:17]
      end else begin
        resetting <= _GEN_470;
      end
    end else begin
      resetting <= _GEN_470;
    end
    flushCounter <= _GEN_489[0]; // @[src/main/scala/rocket/DCache.scala 203:{29,29}]
    if (reset) begin // @[src/main/scala/rocket/DCache.scala 214:33]
      uncachedInFlight_0 <= 1'h0; // @[src/main/scala/rocket/DCache.scala 214:33]
    end else if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        uncachedInFlight_0 <= _GEN_288;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        uncachedInFlight_0 <= _GEN_309;
      end else begin
        uncachedInFlight_0 <= _GEN_288;
      end
    end else begin
      uncachedInFlight_0 <= _GEN_288;
    end
    if (_T_244) begin // @[src/main/scala/rocket/DCache.scala 615:24]
      if (s2_uncached) begin // @[src/main/scala/rocket/DCache.scala 616:24]
        if (a_sel) begin // @[src/main/scala/rocket/DCache.scala 618:18]
          uncachedReqs_0_addr <= s2_req_addr; // @[src/main/scala/rocket/DCache.scala 620:13]
        end
      end
    end
    if (_T_244) begin // @[src/main/scala/rocket/DCache.scala 615:24]
      if (s2_uncached) begin // @[src/main/scala/rocket/DCache.scala 616:24]
        if (a_sel) begin // @[src/main/scala/rocket/DCache.scala 618:18]
          uncachedReqs_0_tag <= s2_req_tag; // @[src/main/scala/rocket/DCache.scala 620:13]
        end
      end
    end
    if (_T_244) begin // @[src/main/scala/rocket/DCache.scala 615:24]
      if (s2_uncached) begin // @[src/main/scala/rocket/DCache.scala 616:24]
        if (a_sel) begin // @[src/main/scala/rocket/DCache.scala 618:18]
          uncachedReqs_0_size <= s2_req_size; // @[src/main/scala/rocket/DCache.scala 620:13]
        end
      end
    end
    if (_T_244) begin // @[src/main/scala/rocket/DCache.scala 615:24]
      if (s2_uncached) begin // @[src/main/scala/rocket/DCache.scala 616:24]
        if (a_sel) begin // @[src/main/scala/rocket/DCache.scala 618:18]
          uncachedReqs_0_signed <= s2_req_signed; // @[src/main/scala/rocket/DCache.scala 620:13]
        end
      end
    end
    line_710_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_711_valid_reg <= _dataArb_io_in_3_valid_T_57;
    line_712_valid_reg <= _T_4;
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 237:30]
      s1_did_read <= dataArb_io_in_3_ready & (io_cpu_req_valid & _dataArb_io_in_3_valid_T_52); // @[src/main/scala/rocket/DCache.scala 237:30]
    end
    line_713_valid_reg <= s0_clk_en;
    if (s0_clk_en) begin // @[src/main/scala/rocket/DCache.scala 238:31]
      s1_read_mask <= dataArb_io_in_3_bits_wordMask; // @[src/main/scala/rocket/DCache.scala 238:31]
    end
    line_714_valid_reg <= s0_clk_en;
    line_715_valid_reg <= _T;
    line_716_valid_reg <= _T_10;
    line_717_valid_reg <= _T_14;
    line_718_valid_reg <= _T_19;
    line_719_valid_reg <= s0_clk_en;
    line_720_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_721_valid_reg <= _T_29;
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        s2_req_addr <= _GEN_174;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
          s2_req_addr <= {{8'd0}, _s2_req_addr_T_1}; // @[src/main/scala/rocket/DCache.scala 683:23]
        end else begin
          s2_req_addr <= _GEN_174;
        end
      end else begin
        s2_req_addr <= _GEN_174;
      end
    end else begin
      s2_req_addr <= _GEN_174;
    end
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        s2_req_tag <= _GEN_175;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
          s2_req_tag <= uncachedReqs_0_tag; // @[src/main/scala/rocket/DCache.scala 682:22]
        end else begin
          s2_req_tag <= _GEN_175;
        end
      end else begin
        s2_req_tag <= _GEN_175;
      end
    end else begin
      s2_req_tag <= _GEN_175;
    end
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        s2_req_size <= _GEN_177;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
          s2_req_size <= uncachedReqs_0_size; // @[src/main/scala/rocket/DCache.scala 680:23]
        end else begin
          s2_req_size <= _GEN_177;
        end
      end else begin
        s2_req_size <= _GEN_177;
      end
    end else begin
      s2_req_size <= _GEN_177;
    end
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (grantIsCached) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        s2_req_signed <= _GEN_178;
      end else if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
        if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
          s2_req_signed <= uncachedReqs_0_signed; // @[src/main/scala/rocket/DCache.scala 681:25]
        end else begin
          s2_req_signed <= _GEN_178;
        end
      end else begin
        s2_req_signed <= _GEN_178;
      end
    end else begin
      s2_req_signed <= _GEN_178;
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_req_dprv <= s1_req_dprv; // @[src/main/scala/rocket/DCache.scala 324:12]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st; // @[src/main/scala/rocket/DCache.scala 326:17]
    end
    if (s1_valid_not_nacked | s1_flush_valid) begin // @[src/main/scala/rocket/DCache.scala 323:48]
      s2_pma_cacheable <= tlb_io_resp_cacheable; // @[src/main/scala/rocket/DCache.scala 327:12]
    end
    if (_T_252) begin // @[src/main/scala/rocket/DCache.scala 658:24]
      if (!(grantIsCached)) begin // @[src/main/scala/rocket/DCache.scala 659:26]
        if (grantIsUncached) begin // @[src/main/scala/rocket/DCache.scala 668:35]
          if (grantIsUncachedData) begin // @[src/main/scala/rocket/DCache.scala 675:34]
            s2_uncached_resp_addr <= uncachedReqs_0_addr; // @[src/main/scala/rocket/DCache.scala 688:33]
          end
        end
      end
    end
    line_722_valid_reg <= _T_30;
    if (_T_30) begin // @[src/main/scala/rocket/DCache.scala 329:31]
      s2_vaddr_r <= s1_vaddr; // @[src/main/scala/rocket/DCache.scala 329:31]
    end
    line_723_valid_reg <= _T_30;
    s2_flush_valid_pre_tag_ecc <= s1_flush_valid; // @[src/main/scala/rocket/DCache.scala 333:43]
    line_724_valid_reg <= s1_meta_clk_en;
    line_725_valid_reg <= s1_meta_clk_en;
    if (s1_meta_clk_en) begin // @[src/main/scala/rocket/DCache.scala 339:61]
      s2_meta_corrected_r <= tag_array_0_s1_meta_data; // @[src/main/scala/rocket/DCache.scala 339:61]
    end
    line_726_valid_reg <= s1_meta_clk_en;
    if (grantIsUncachedData & (blockUncachedGrant | s1_valid)) begin // @[src/main/scala/rocket/DCache.scala 736:68]
      if (auto_out_d_valid) begin // @[src/main/scala/rocket/DCache.scala 739:29]
        blockUncachedGrant <= _T_272; // @[src/main/scala/rocket/DCache.scala 743:28]
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid; // @[src/main/scala/rocket/DCache.scala 735:24]
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid; // @[src/main/scala/rocket/DCache.scala 735:24]
    end
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_T_252) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (d_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (beats1_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          counter <= beats1_decode;
        end else begin
          counter <= 2'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (s2_data_en) begin // @[src/main/scala/rocket/DCache.scala 357:18]
      s2_data <= _s2_data_T_6; // @[src/main/scala/rocket/DCache.scala 357:18]
    end
    line_727_valid_reg <= s2_data_en;
    line_728_valid_reg <= s1_probe;
    line_729_valid_reg <= s1_probe;
    line_730_valid_reg <= s1_valid_not_nacked;
    line_731_valid_reg <= _T_30;
    line_732_valid_reg <= s1_valid_not_nacked;
    line_733_valid_reg <= _T_30;
    line_734_valid_reg <= _T_223;
    if (s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_48 & _io_cpu_req_ready_T_1 | s2_valid_cached_miss) begin // @[src/main/scala/rocket/DCache.scala 456:99]
      lrscAddr <= s2_req_addr[39:5]; // @[src/main/scala/rocket/DCache.scala 458:14]
    end
    line_735_valid_reg <= _T_227;
    line_736_valid_reg <= _lrscBackingOff_T;
    line_737_valid_reg <= _T_231;
    line_738_valid_reg <= s1_probe;
    if (s1_valid_not_nacked & s1_write) begin // @[src/main/scala/rocket/DCache.scala 476:30]
      pstore1_cmd <= s1_req_cmd; // @[src/main/scala/rocket/DCache.scala 476:30]
    end
    line_739_valid_reg <= _pstore1_cmd_T;
    line_740_valid_reg <= _pstore1_cmd_T;
    if (_pstore1_cmd_T) begin // @[src/main/scala/rocket/DCache.scala 478:31]
      pstore1_data <= io_cpu_s1_data_data; // @[src/main/scala/rocket/DCache.scala 478:31]
    end
    line_741_valid_reg <= _pstore1_cmd_T;
    line_742_valid_reg <= _pstore1_cmd_T;
    line_743_valid_reg <= _pstore1_cmd_T;
    if (_pstore1_cmd_T) begin // @[src/main/scala/rocket/DCache.scala 482:44]
      pstore1_rmw_r <= _pstore1_rmw_T_52; // @[src/main/scala/rocket/DCache.scala 482:44]
    end
    line_744_valid_reg <= _pstore1_cmd_T;
    line_745_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_746_valid_reg <= _dataArb_io_in_3_valid_T_57;
    pstore_drain_on_miss_REG <= io_cpu_s2_nack; // @[src/main/scala/rocket/DCache.scala 487:56]
    line_747_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_748_valid_reg <= _T_240;
    line_749_valid_reg <= advance_pstore1;
    line_750_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r <= pstore1_storegen_data[7:0]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_751_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_1 <= pstore1_storegen_data[15:8]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_752_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_2 <= pstore1_storegen_data[23:16]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_753_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_3 <= pstore1_storegen_data[31:24]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_754_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_4 <= pstore1_storegen_data[39:32]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_755_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_5 <= pstore1_storegen_data[47:40]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_756_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_6 <= pstore1_storegen_data[55:48]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_757_valid_reg <= advance_pstore1;
    if (advance_pstore1) begin // @[src/main/scala/rocket/DCache.scala 512:22]
      pstore2_storegen_data_r_7 <= pstore1_storegen_data[63:56]; // @[src/main/scala/rocket/DCache.scala 512:22]
    end
    line_758_valid_reg <= advance_pstore1;
    line_759_valid_reg <= advance_pstore1;
    line_760_valid_reg <= _T_243;
    line_761_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_762_valid_reg <= _atomics_T_6;
    line_763_valid_reg <= _T_244;
    line_764_valid_reg <= s2_uncached;
    line_765_valid_reg <= a_sel;
    line_766_valid_reg <= s2_uncached;
    line_767_valid_reg <= _T_252;
    line_768_valid_reg <= _block_probe_for_core_progress_T;
    line_769_valid_reg <= _T_252;
    line_770_valid_reg <= grantIsCached;
    line_771_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_772_valid_reg <= _io_cpu_req_ready_T_1;
    line_773_valid_reg <= d_last;
    line_774_valid_reg <= grantIsCached;
    line_775_valid_reg <= grantIsUncached;
    line_776_valid_reg <= _T_257;
    line_777_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_778_valid_reg <= _a_source_T;
    line_779_valid_reg <= grantIsUncachedData;
    line_780_valid_reg <= grantIsUncached;
    line_781_valid_reg <= grantIsVoluntary;
    line_782_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_783_valid_reg <= _tl_out_a_valid_T_7;
    line_784_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_785_valid_reg <= _T_271;
    line_786_valid_reg <= _T_273;
    line_787_valid_reg <= _T_275;
    line_788_valid_reg <= auto_out_d_valid;
    line_789_valid_reg <= _T_278;
    s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    line_790_valid_reg <= s2_want_victimize;
    line_791_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_792_valid_reg <= _T_283;
    line_793_valid_reg <= s2_probe;
    line_794_valid_reg <= s2_prb_ack_data;
    line_795_valid_reg <= s2_prb_ack_data;
    line_796_valid_reg <= _T_284;
    line_797_valid_reg <= _T_284;
    line_798_valid_reg <= probeNack;
    line_799_valid_reg <= _T_285;
    line_800_valid_reg <= metaArb_io_in_6_ready;
    line_801_valid_reg <= _T_286;
    line_802_valid_reg <= releaseDone;
    line_803_valid_reg <= _T_287;
    line_804_valid_reg <= releaseDone;
    line_805_valid_reg <= _T_288;
    line_806_valid_reg <= releaseDone;
    line_807_valid_reg <= _T_293;
    line_808_valid_reg <= _T_291;
    line_809_valid_reg <= _T_291;
    line_810_valid_reg <= releaseDone;
    line_811_valid_reg <= _T_296;
    line_812_valid_reg <= _T_297;
    io_cpu_s2_xcpt_REG <= tlb_io_req_valid & _s1_valid_not_nacked_T; // @[src/main/scala/rocket/DCache.scala 915:65]
    line_813_valid_reg <= io_cpu_replay_next;
    doUncachedResp <= io_cpu_replay_next; // @[src/main/scala/rocket/DCache.scala 931:31]
    line_814_valid_reg <= doUncachedResp;
    line_815_valid_reg <= _dataArb_io_in_3_valid_T_56;
    line_816_valid_reg <= _T_303;
    REG <= reset; // @[src/main/scala/rocket/DCache.scala 1005:25]
    line_817_valid_reg <= REG;
    line_818_valid_reg <= resetting;
    line_819_valid_reg <= flushDone;
    line_820_valid_reg <= _T_244;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      io_cpu_perf_release_counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (_T_278) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (io_cpu_perf_release_first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (beats1_opdata_1) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          io_cpu_perf_release_counter <= beats1_decode_1;
        end else begin
          io_cpu_perf_release_counter <= 2'h0;
        end
      end else begin
        io_cpu_perf_release_counter <= io_cpu_perf_release_counter1;
      end
    end
    line_821_valid_reg <= _T_278;
    line_822_valid_reg <= _io_cpu_perf_blocked_near_end_of_refill_T_1;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_dataArb_io_in_3_valid_T_52 | dataArb_io_in_3_valid_res)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1183 assert(!needsRead(req) || res)\n"); // @[src/main/scala/rocket/DCache.scala 1183:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(~(s1_valid_masked & _s1_write_T_1) | &_T_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:307 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n"
            ); // @[src/main/scala/rocket/DCache.scala 307:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_dataArb_io_in_3_valid_T_52 | dataArb_io_in_3_valid_res)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1183 assert(!needsRead(req) || res)\n"); // @[src/main/scala/rocket/DCache.scala 1183:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(pstore1_rmw_r | _T_235 == pstore1_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:494 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"
            ); // @[src/main/scala/rocket/DCache.scala 494:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(~(tl_out_a_valid & s2_read & s2_write & s2_uncached))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:583 assert (!(tl_out_a.valid && s2_read && s2_write && s2_uncached))\n"
            ); // @[src/main/scala/rocket/DCache.scala 583:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_252 & grantIsCached & _dataArb_io_in_3_valid_T_56 & _io_cpu_req_ready_T_1) begin
          $fwrite(32'h80000002,
            "Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:661 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"
            ); // @[src/main/scala/rocket/DCache.scala 661:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_252 & _T_313 & grantIsUncached & _T_257 & _dataArb_io_in_3_valid_T_56 & _a_source_T) begin
          $fwrite(32'h80000002,
            "Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:671 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"
            ); // @[src/main/scala/rocket/DCache.scala 671:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_494 & _tl_d_data_encoded_T_11 & grantIsVoluntary & _dataArb_io_in_3_valid_T_56 & _tl_out_a_valid_T_7
          ) begin
          $fwrite(32'h80000002,
            "Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:692 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"
            ); // @[src/main/scala/rocket/DCache.scala 692:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_dataArb_io_in_3_valid_T_56 & ~(_T_264 == (_T_252 & d_first & grantIsCached))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:700 assert(tl_out.e.fire === (tl_out.d.fire && d_first && grantIsCached))\n"
            ); // @[src/main/scala/rocket/DCache.scala 700:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_want_victimize & _dataArb_io_in_3_valid_T_56 & ~(s2_valid_flush_line | s2_flush_valid_pre_tag_ecc |
          io_cpu_s2_nack)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at DCache.scala:801 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n"
            ); // @[src/main/scala/rocket/DCache.scala 801:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & _dataArb_io_in_3_valid_T_56 & ~_io_cpu_s2_nack_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:935 assert(!s2_valid_hit)\n"); // @[src/main/scala/rocket/DCache.scala 935:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[27:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_s1_meta_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_s1_meta_addr_pipe_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s1_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  lrscCount = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  s1_probe = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s2_probe = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  release_state = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  release_ack_wait = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  release_ack_addr = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  grantInProgress = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s2_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  probe_bits_param = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  probe_bits_size = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  probe_bits_source = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  probe_bits_address = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  line_706_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  counter_1 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s1_req_cmd = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  s2_req_cmd = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  pstore1_held = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  pstore1_addr = _RAND_24[39:0];
  _RAND_25 = {2{`RANDOM}};
  s1_req_addr = _RAND_25[39:0];
  _RAND_26 = {1{`RANDOM}};
  pstore1_mask = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  s1_req_size = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  pstore2_valid = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  pstore2_addr = _RAND_29[39:0];
  _RAND_30 = {1{`RANDOM}};
  pstore2_storegen_mask = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  line_707_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  s1_req_tag = _RAND_34[6:0];
  _RAND_35 = {1{`RANDOM}};
  s1_req_signed = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  s1_req_dprv = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  line_708_valid_reg = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_38[39:0];
  _RAND_39 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  s1_tlb_req_prv = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  line_709_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  s1_flush_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  cached_grant_wait = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  resetting = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  flushCounter = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_48[0:0];
  _RAND_49 = {2{`RANDOM}};
  uncachedReqs_0_addr = _RAND_49[39:0];
  _RAND_50 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_50[6:0];
  _RAND_51 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_710_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_711_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_712_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  s1_did_read = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_713_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  s1_read_mask = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_714_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_715_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_716_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_717_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_718_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_719_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_720_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_721_valid_reg = _RAND_66[0:0];
  _RAND_67 = {2{`RANDOM}};
  s2_req_addr = _RAND_67[39:0];
  _RAND_68 = {1{`RANDOM}};
  s2_req_tag = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  s2_req_size = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  s2_req_signed = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  s2_req_dprv = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_78[0:0];
  _RAND_79 = {2{`RANDOM}};
  s2_uncached_resp_addr = _RAND_79[39:0];
  _RAND_80 = {1{`RANDOM}};
  line_722_valid_reg = _RAND_80[0:0];
  _RAND_81 = {2{`RANDOM}};
  s2_vaddr_r = _RAND_81[39:0];
  _RAND_82 = {1{`RANDOM}};
  line_723_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  s2_flush_valid_pre_tag_ecc = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_724_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_725_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  s2_meta_corrected_r = _RAND_86[27:0];
  _RAND_87 = {1{`RANDOM}};
  line_726_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  counter = _RAND_89[1:0];
  _RAND_90 = {2{`RANDOM}};
  s2_data = _RAND_90[63:0];
  _RAND_91 = {1{`RANDOM}};
  line_727_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_728_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_729_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_730_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_731_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_732_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_733_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_734_valid_reg = _RAND_98[0:0];
  _RAND_99 = {2{`RANDOM}};
  lrscAddr = _RAND_99[34:0];
  _RAND_100 = {1{`RANDOM}};
  line_735_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_736_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_737_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_738_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  pstore1_cmd = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  line_739_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_740_valid_reg = _RAND_106[0:0];
  _RAND_107 = {2{`RANDOM}};
  pstore1_data = _RAND_107[63:0];
  _RAND_108 = {1{`RANDOM}};
  line_741_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_742_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_743_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  pstore1_rmw_r = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_744_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_745_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_746_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  pstore_drain_on_miss_REG = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_747_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_748_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_749_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_750_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  pstore2_storegen_data_r = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  line_751_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  pstore2_storegen_data_r_1 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  line_752_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  pstore2_storegen_data_r_2 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  line_753_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  pstore2_storegen_data_r_3 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  line_754_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  pstore2_storegen_data_r_4 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  line_755_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  pstore2_storegen_data_r_5 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  line_756_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  pstore2_storegen_data_r_6 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  line_757_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  pstore2_storegen_data_r_7 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  line_758_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_759_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_760_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_761_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_762_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_763_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_764_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_765_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_766_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_767_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_768_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_769_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_770_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_771_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_772_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_773_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_774_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_775_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_776_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_777_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_778_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_779_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_780_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_781_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_782_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_783_valid_reg = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  line_784_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  line_785_valid_reg = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  line_786_valid_reg = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  line_787_valid_reg = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  line_788_valid_reg = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  line_789_valid_reg = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  line_790_valid_reg = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  line_791_valid_reg = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  line_792_valid_reg = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  line_793_valid_reg = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  line_794_valid_reg = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  line_795_valid_reg = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  line_796_valid_reg = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  line_797_valid_reg = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  line_798_valid_reg = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  line_799_valid_reg = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  line_800_valid_reg = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  line_801_valid_reg = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  line_802_valid_reg = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  line_803_valid_reg = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  line_804_valid_reg = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  line_805_valid_reg = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  line_806_valid_reg = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  line_807_valid_reg = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  line_808_valid_reg = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  line_809_valid_reg = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  line_810_valid_reg = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  line_811_valid_reg = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  line_812_valid_reg = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  io_cpu_s2_xcpt_REG = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  line_813_valid_reg = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  doUncachedResp = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  line_814_valid_reg = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  line_815_valid_reg = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  line_816_valid_reg = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  REG = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  line_817_valid_reg = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  line_818_valid_reg = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  line_819_valid_reg = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  line_820_valid_reg = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  io_cpu_perf_release_counter = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  line_821_valid_reg = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  line_822_valid_reg = _RAND_204[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~_dataArb_io_in_3_valid_T_52 | dataArb_io_in_3_valid_res); // @[src/main/scala/rocket/DCache.scala 1183:11]
    end
    //
    if (_dataArb_io_in_3_valid_T_56) begin
      assert(~(s1_valid_masked & _s1_write_T_1) | &_T_24); // @[src/main/scala/rocket/DCache.scala 307:9]
    end
    //
    if (~reset) begin
      assert(~_dataArb_io_in_3_valid_T_52 | dataArb_io_in_3_valid_res); // @[src/main/scala/rocket/DCache.scala 1183:11]
    end
    //
    if (_dataArb_io_in_3_valid_T_56) begin
      assert(pstore1_rmw_r | _T_235 == pstore1_valid); // @[src/main/scala/rocket/DCache.scala 494:9]
    end
    //
    if (_dataArb_io_in_3_valid_T_56) begin
      assert(~(tl_out_a_valid & s2_read & s2_write & s2_uncached)); // @[src/main/scala/rocket/DCache.scala 583:12]
    end
    //
    if (_T_252 & grantIsCached & _dataArb_io_in_3_valid_T_56) begin
      assert(cached_grant_wait); // @[src/main/scala/rocket/DCache.scala 661:13]
    end
    //
    if (_T_252 & _T_313 & grantIsUncached & _T_257 & _dataArb_io_in_3_valid_T_56) begin
      assert(uncachedInFlight_0); // @[src/main/scala/rocket/DCache.scala 671:17]
    end
    //
    if (_GEN_494 & _tl_d_data_encoded_T_11 & grantIsVoluntary & _dataArb_io_in_3_valid_T_56) begin
      assert(release_ack_wait); // @[src/main/scala/rocket/DCache.scala 692:13]
    end
    //
    if (_dataArb_io_in_3_valid_T_56) begin
      assert(_T_264 == (_T_252 & d_first & grantIsCached)); // @[src/main/scala/rocket/DCache.scala 700:9]
    end
    //
    if (s2_want_victimize & _dataArb_io_in_3_valid_T_56) begin
      assert(s2_valid_flush_line | s2_flush_valid_pre_tag_ecc | io_cpu_s2_nack); // @[src/main/scala/rocket/DCache.scala 801:13]
    end
    //
    if (doUncachedResp & _dataArb_io_in_3_valid_T_56) begin
      assert(_io_cpu_s2_nack_T_4); // @[src/main/scala/rocket/DCache.scala 935:11]
    end
  end
endmodule
module ICache(
  input         clock,
  input         reset,
  input         auto_master_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_master_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_master_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_master_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_master_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_master_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_master_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_master_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        io_req_ready, // @[src/main/scala/rocket/ICache.scala 248:14]
  input         io_req_valid, // @[src/main/scala/rocket/ICache.scala 248:14]
  input  [38:0] io_req_bits_addr, // @[src/main/scala/rocket/ICache.scala 248:14]
  input  [31:0] io_s1_paddr, // @[src/main/scala/rocket/ICache.scala 248:14]
  input         io_s1_kill, // @[src/main/scala/rocket/ICache.scala 248:14]
  input         io_s2_kill, // @[src/main/scala/rocket/ICache.scala 248:14]
  output        io_resp_valid, // @[src/main/scala/rocket/ICache.scala 248:14]
  output [31:0] io_resp_bits_data, // @[src/main/scala/rocket/ICache.scala 248:14]
  output        io_resp_bits_ae, // @[src/main/scala/rocket/ICache.scala 248:14]
  input         io_invalidate // @[src/main/scala/rocket/ICache.scala 248:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] tag_array_0 [0:1]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_tag_rdata_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_tag_rdata_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [26:0] tag_array_0_tag_rdata_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [26:0] tag_array_0_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  tag_array_0_MPORT_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  tag_array_0_tag_rdata_en_pipe_0;
  reg  tag_array_0_tag_rdata_addr_pipe_0;
  reg [31:0] data_arrays_0_0 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_dout_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_0_dout_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [31:0] data_arrays_0_0_dout_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [31:0] data_arrays_0_0_MPORT_1_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_0_0_MPORT_1_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_MPORT_1_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_0_0_MPORT_1_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_0_0_dout_en_pipe_0;
  reg [2:0] data_arrays_0_0_dout_addr_pipe_0;
  reg [31:0] data_arrays_1_0 [0:7]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_1_0_dout_1_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_1_0_dout_1_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [31:0] data_arrays_1_0_dout_1_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [31:0] data_arrays_1_0_MPORT_2_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire [2:0] data_arrays_1_0_MPORT_2_addr; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_1_0_MPORT_2_mask; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  wire  data_arrays_1_0_MPORT_2_en; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  reg  data_arrays_1_0_dout_1_en_pipe_0;
  reg [2:0] data_arrays_1_0_dout_1_addr_pipe_0;
  wire  s0_valid = io_req_ready & io_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  s1_valid; // @[src/main/scala/rocket/ICache.scala 333:25]
  wire  line_823_clock;
  wire  line_823_reset;
  wire  line_823_valid;
  reg  line_823_valid_reg;
  reg [1:0] vb_array; // @[src/main/scala/rocket/ICache.scala 440:25]
  wire  s1_idx = io_s1_paddr[5]; // @[src/main/scala/rocket/ICache.scala 851:21]
  wire [1:0] _s1_vb_T = {1'h0,s1_idx}; // @[src/main/scala/rocket/ICache.scala 500:29]
  wire [1:0] _s1_vb_T_1 = vb_array >> _s1_vb_T; // @[src/main/scala/rocket/ICache.scala 500:25]
  wire  s1_vb = _s1_vb_T_1[0]; // @[src/main/scala/rocket/ICache.scala 500:25]
  wire [25:0] tag = tag_array_0_tag_rdata_data[25:0]; // @[src/main/scala/util/package.scala 155:13]
  wire [25:0] s1_tag = io_s1_paddr[31:6]; // @[src/main/scala/rocket/ICache.scala 485:30]
  wire  tagMatch = s1_vb & tag == s1_tag; // @[src/main/scala/rocket/ICache.scala 506:26]
  wire  _s1_tag_hit_0_T = tagMatch; // @[src/main/scala/rocket/ICache.scala 506:26]
  wire  s1_hit = tagMatch; // @[src/main/scala/rocket/ICache.scala 506:26]
  reg  s2_valid; // @[src/main/scala/rocket/ICache.scala 355:25]
  reg  s2_hit; // @[src/main/scala/rocket/ICache.scala 356:23]
  reg  invalidated; // @[src/main/scala/rocket/ICache.scala 359:24]
  reg  refill_valid; // @[src/main/scala/rocket/ICache.scala 360:29]
  wire  s2_miss = s2_valid & ~s2_hit & ~io_s2_kill; // @[src/main/scala/rocket/ICache.scala 370:37]
  reg  s2_request_refill_REG; // @[src/main/scala/rocket/ICache.scala 377:45]
  wire  s2_request_refill = s2_miss & s2_request_refill_REG; // @[src/main/scala/rocket/ICache.scala 377:35]
  wire  refill_fire = auto_master_out_a_ready & s2_request_refill; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  s1_can_request_refill = ~(s2_miss | refill_valid); // @[src/main/scala/rocket/ICache.scala 372:31]
  wire  _refill_paddr_T = s1_valid & s1_can_request_refill; // @[src/main/scala/rocket/ICache.scala 378:54]
  reg [31:0] refill_paddr; // @[src/main/scala/rocket/ICache.scala 378:31]
  wire  line_824_clock;
  wire  line_824_reset;
  wire  line_824_valid;
  reg  line_824_valid_reg;
  wire  line_825_clock;
  wire  line_825_reset;
  wire  line_825_valid;
  reg  line_825_valid_reg;
  wire [25:0] refill_tag = refill_paddr[31:6]; // @[src/main/scala/rocket/ICache.scala 380:33]
  wire  refill_idx = refill_paddr[5]; // @[src/main/scala/rocket/ICache.scala 851:21]
  wire  refill_one_beat_opdata = auto_master_out_d_bits_opcode[0]; // @[src/main/scala/tilelink/Edges.scala 106:36]
  wire  refill_one_beat = auto_master_out_d_valid & refill_one_beat_opdata; // @[src/main/scala/rocket/ICache.scala 383:39]
  wire [11:0] _beats1_decode_T_1 = 12'h1f << auto_master_out_d_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [4:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[4:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [1:0] beats1_decode = _beats1_decode_T_3[4:3]; // @[src/main/scala/tilelink/Edges.scala 220:59]
  wire [1:0] beats1 = refill_one_beat_opdata ? beats1_decode : 2'h0; // @[src/main/scala/tilelink/Edges.scala 221:14]
  reg [1:0] counter; // @[src/main/scala/tilelink/Edges.scala 229:27]
  wire [1:0] counter1 = counter - 2'h1; // @[src/main/scala/tilelink/Edges.scala 230:28]
  wire  first = counter == 2'h0; // @[src/main/scala/tilelink/Edges.scala 231:25]
  wire  last = counter == 2'h1 | beats1 == 2'h0; // @[src/main/scala/tilelink/Edges.scala 232:33]
  wire  d_done = last & auto_master_out_d_valid; // @[src/main/scala/tilelink/Edges.scala 233:22]
  wire [1:0] _count_T = ~counter1; // @[src/main/scala/tilelink/Edges.scala 234:27]
  wire [1:0] refill_cnt = beats1 & _count_T; // @[src/main/scala/tilelink/Edges.scala 234:25]
  wire  line_826_clock;
  wire  line_826_reset;
  wire  line_826_valid;
  reg  line_826_valid_reg;
  wire  refill_done = refill_one_beat & d_done; // @[src/main/scala/rocket/ICache.scala 391:37]
  wire  _tag_rdata_T_1 = ~refill_done; // @[src/main/scala/rocket/ICache.scala 418:70]
  wire  _tag_rdata_T_2 = ~refill_done & s0_valid; // @[src/main/scala/rocket/ICache.scala 418:83]
  wire  line_827_clock;
  wire  line_827_reset;
  wire  line_827_valid;
  reg  line_827_valid_reg;
  reg  accruedRefillError; // @[src/main/scala/rocket/ICache.scala 420:31]
  wire  refillError = auto_master_out_d_bits_corrupt | refill_cnt > 2'h0 & accruedRefillError; // @[src/main/scala/rocket/ICache.scala 422:43]
  wire  line_828_clock;
  wire  line_828_reset;
  wire  line_828_valid;
  reg  line_828_valid_reg;
  wire  line_829_clock;
  wire  line_829_reset;
  wire  line_829_valid;
  reg  line_829_valid_reg;
  wire [1:0] _vb_array_T = {1'h0,refill_idx}; // @[src/main/scala/rocket/ICache.scala 444:36]
  wire  _vb_array_T_1 = ~invalidated; // @[src/main/scala/rocket/ICache.scala 444:75]
  wire [3:0] _vb_array_T_3 = 4'h1 << _vb_array_T; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _GEN_82 = {{2'd0}, vb_array}; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _vb_array_T_4 = _GEN_82 | _vb_array_T_3; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [1:0] _vb_array_T_5 = ~vb_array; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _GEN_83 = {{2'd0}, _vb_array_T_5}; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _vb_array_T_6 = _GEN_83 | _vb_array_T_3; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _vb_array_T_7 = ~_vb_array_T_6; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _vb_array_T_8 = refill_done & ~invalidated ? _vb_array_T_4 : _vb_array_T_7; // @[src/main/scala/rocket/ICache.scala 444:32]
  wire [3:0] _GEN_46 = refill_one_beat ? _vb_array_T_8 : {{2'd0}, vb_array}; // @[src/main/scala/rocket/ICache.scala 441:26 444:14 440:25]
  wire  line_830_clock;
  wire  line_830_reset;
  wire  line_830_valid;
  reg  line_830_valid_reg;
  wire [3:0] _GEN_47 = io_invalidate ? 4'h0 : _GEN_46; // @[src/main/scala/rocket/ICache.scala 449:21 450:14]
  wire  _GEN_48 = io_invalidate | invalidated; // @[src/main/scala/rocket/ICache.scala 449:21 451:17 359:24]
  wire  tl_error = tag_array_0_tag_rdata_data[26]; // @[src/main/scala/util/package.scala 155:13]
  wire  s1_tl_error_0 = tagMatch & tl_error; // @[src/main/scala/rocket/ICache.scala 510:32]
  wire  _T_9 = ~reset; // @[src/main/scala/rocket/ICache.scala 513:9]
  wire  line_831_clock;
  wire  line_831_reset;
  wire  line_831_valid;
  reg  line_831_valid_reg;
  wire  _s0_ren_T_1 = ~io_req_bits_addr[2]; // @[src/main/scala/rocket/ICache.scala 556:111]
  wire  s0_ren = s0_valid & _s0_ren_T_1; // @[src/main/scala/rocket/ICache.scala 559:28]
  wire  wen = refill_one_beat & _vb_array_T_1; // @[src/main/scala/rocket/ICache.scala 562:32]
  wire [2:0] _mem_idx_T = {refill_idx, 2'h0}; // @[src/main/scala/rocket/ICache.scala 566:40]
  wire [2:0] _GEN_84 = {{1'd0}, refill_cnt}; // @[src/main/scala/rocket/ICache.scala 566:67]
  wire [2:0] _mem_idx_T_1 = _mem_idx_T | _GEN_84; // @[src/main/scala/rocket/ICache.scala 566:67]
  wire  line_832_clock;
  wire  line_832_reset;
  wire  line_832_valid;
  reg  line_832_valid_reg;
  wire  _dout_T = ~wen; // @[src/main/scala/rocket/ICache.scala 582:41]
  wire  _dout_T_1 = ~wen & s0_ren; // @[src/main/scala/rocket/ICache.scala 582:46]
  wire  line_833_clock;
  wire  line_833_reset;
  wire  line_833_valid;
  reg  line_833_valid_reg;
  wire  _T_14 = ~io_s1_paddr[2]; // @[src/main/scala/rocket/ICache.scala 556:111]
  wire  line_834_clock;
  wire  line_834_reset;
  wire  line_834_valid;
  reg  line_834_valid_reg;
  wire [31:0] _GEN_60 = data_arrays_0_0_dout_data; // @[src/main/scala/rocket/ICache.scala 584:71 585:15]
  wire  s0_ren_1 = s0_valid & io_req_bits_addr[2]; // @[src/main/scala/rocket/ICache.scala 559:28]
  wire  line_835_clock;
  wire  line_835_reset;
  wire  line_835_valid;
  reg  line_835_valid_reg;
  wire  _dout_T_5 = ~wen & s0_ren_1; // @[src/main/scala/rocket/ICache.scala 582:46]
  wire  line_836_clock;
  wire  line_836_reset;
  wire  line_836_valid;
  reg  line_836_valid_reg;
  wire  line_837_clock;
  wire  line_837_reset;
  wire  line_837_valid;
  reg  line_837_valid_reg;
  wire  line_838_clock;
  wire  line_838_reset;
  wire  line_838_valid;
  reg  line_838_valid_reg;
  reg [31:0] s2_dout_0; // @[src/main/scala/rocket/ICache.scala 604:26]
  wire  line_839_clock;
  wire  line_839_reset;
  wire  line_839_valid;
  reg  line_839_valid_reg;
  wire  line_840_clock;
  wire  line_840_reset;
  wire  line_840_valid;
  reg  line_840_valid_reg;
  reg  s2_tl_error; // @[src/main/scala/rocket/ICache.scala 607:30]
  wire  line_841_clock;
  wire  line_841_reset;
  wire  line_841_valid;
  reg  line_841_valid_reg;
  wire  line_842_clock;
  wire  line_842_reset;
  wire  line_842_valid;
  reg  line_842_valid_reg;
  wire  line_843_clock;
  wire  line_843_reset;
  wire  line_843_valid;
  reg  line_843_valid_reg;
  wire  _T_25 = ~refill_valid; // @[src/main/scala/rocket/ICache.scala 821:9]
  wire  line_844_clock;
  wire  line_844_reset;
  wire  line_844_valid;
  reg  line_844_valid_reg;
  wire  line_845_clock;
  wire  line_845_reset;
  wire  line_845_valid;
  reg  line_845_valid_reg;
  wire  _GEN_80 = refill_fire | refill_valid; // @[src/main/scala/rocket/ICache.scala 822:22 360:29 822:37]
  wire  line_846_clock;
  wire  line_846_reset;
  wire  line_846_valid;
  reg  line_846_valid_reg;
  wire [3:0] _GEN_86 = reset ? 4'h0 : _GEN_47; // @[src/main/scala/rocket/ICache.scala 440:{25,25}]
  GEN_w1_line #(.COVER_INDEX(823)) line_823 (
    .clock(line_823_clock),
    .reset(line_823_reset),
    .valid(line_823_valid)
  );
  GEN_w1_line #(.COVER_INDEX(824)) line_824 (
    .clock(line_824_clock),
    .reset(line_824_reset),
    .valid(line_824_valid)
  );
  GEN_w1_line #(.COVER_INDEX(825)) line_825 (
    .clock(line_825_clock),
    .reset(line_825_reset),
    .valid(line_825_valid)
  );
  GEN_w1_line #(.COVER_INDEX(826)) line_826 (
    .clock(line_826_clock),
    .reset(line_826_reset),
    .valid(line_826_valid)
  );
  GEN_w1_line #(.COVER_INDEX(827)) line_827 (
    .clock(line_827_clock),
    .reset(line_827_reset),
    .valid(line_827_valid)
  );
  GEN_w1_line #(.COVER_INDEX(828)) line_828 (
    .clock(line_828_clock),
    .reset(line_828_reset),
    .valid(line_828_valid)
  );
  GEN_w1_line #(.COVER_INDEX(829)) line_829 (
    .clock(line_829_clock),
    .reset(line_829_reset),
    .valid(line_829_valid)
  );
  GEN_w1_line #(.COVER_INDEX(830)) line_830 (
    .clock(line_830_clock),
    .reset(line_830_reset),
    .valid(line_830_valid)
  );
  GEN_w1_line #(.COVER_INDEX(831)) line_831 (
    .clock(line_831_clock),
    .reset(line_831_reset),
    .valid(line_831_valid)
  );
  GEN_w1_line #(.COVER_INDEX(832)) line_832 (
    .clock(line_832_clock),
    .reset(line_832_reset),
    .valid(line_832_valid)
  );
  GEN_w1_line #(.COVER_INDEX(833)) line_833 (
    .clock(line_833_clock),
    .reset(line_833_reset),
    .valid(line_833_valid)
  );
  GEN_w1_line #(.COVER_INDEX(834)) line_834 (
    .clock(line_834_clock),
    .reset(line_834_reset),
    .valid(line_834_valid)
  );
  GEN_w1_line #(.COVER_INDEX(835)) line_835 (
    .clock(line_835_clock),
    .reset(line_835_reset),
    .valid(line_835_valid)
  );
  GEN_w1_line #(.COVER_INDEX(836)) line_836 (
    .clock(line_836_clock),
    .reset(line_836_reset),
    .valid(line_836_valid)
  );
  GEN_w1_line #(.COVER_INDEX(837)) line_837 (
    .clock(line_837_clock),
    .reset(line_837_reset),
    .valid(line_837_valid)
  );
  GEN_w1_line #(.COVER_INDEX(838)) line_838 (
    .clock(line_838_clock),
    .reset(line_838_reset),
    .valid(line_838_valid)
  );
  GEN_w1_line #(.COVER_INDEX(839)) line_839 (
    .clock(line_839_clock),
    .reset(line_839_reset),
    .valid(line_839_valid)
  );
  GEN_w1_line #(.COVER_INDEX(840)) line_840 (
    .clock(line_840_clock),
    .reset(line_840_reset),
    .valid(line_840_valid)
  );
  GEN_w1_line #(.COVER_INDEX(841)) line_841 (
    .clock(line_841_clock),
    .reset(line_841_reset),
    .valid(line_841_valid)
  );
  GEN_w1_line #(.COVER_INDEX(842)) line_842 (
    .clock(line_842_clock),
    .reset(line_842_reset),
    .valid(line_842_valid)
  );
  GEN_w1_line #(.COVER_INDEX(843)) line_843 (
    .clock(line_843_clock),
    .reset(line_843_reset),
    .valid(line_843_valid)
  );
  GEN_w1_line #(.COVER_INDEX(844)) line_844 (
    .clock(line_844_clock),
    .reset(line_844_reset),
    .valid(line_844_valid)
  );
  GEN_w1_line #(.COVER_INDEX(845)) line_845 (
    .clock(line_845_clock),
    .reset(line_845_reset),
    .valid(line_845_valid)
  );
  GEN_w1_line #(.COVER_INDEX(846)) line_846 (
    .clock(line_846_clock),
    .reset(line_846_reset),
    .valid(line_846_valid)
  );
  assign tag_array_0_tag_rdata_en = tag_array_0_tag_rdata_en_pipe_0;
  assign tag_array_0_tag_rdata_addr = tag_array_0_tag_rdata_addr_pipe_0;
  assign tag_array_0_tag_rdata_data = tag_array_0[tag_array_0_tag_rdata_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign tag_array_0_MPORT_data = {refillError,refill_tag};
  assign tag_array_0_MPORT_addr = refill_paddr[5];
  assign tag_array_0_MPORT_mask = 1'h1;
  assign tag_array_0_MPORT_en = refill_one_beat & d_done;
  assign data_arrays_0_0_dout_en = data_arrays_0_0_dout_en_pipe_0;
  assign data_arrays_0_0_dout_addr = data_arrays_0_0_dout_addr_pipe_0;
  assign data_arrays_0_0_dout_data = data_arrays_0_0[data_arrays_0_0_dout_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_0_0_MPORT_1_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_0_MPORT_1_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[5:3];
  assign data_arrays_0_0_MPORT_1_mask = 1'h1;
  assign data_arrays_0_0_MPORT_1_en = refill_one_beat & _vb_array_T_1;
  assign data_arrays_1_0_dout_1_en = data_arrays_1_0_dout_1_en_pipe_0;
  assign data_arrays_1_0_dout_1_addr = data_arrays_1_0_dout_1_addr_pipe_0;
  assign data_arrays_1_0_dout_1_data = data_arrays_1_0[data_arrays_1_0_dout_1_addr]; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
  assign data_arrays_1_0_MPORT_2_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_0_MPORT_2_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[5:3];
  assign data_arrays_1_0_MPORT_2_mask = 1'h1;
  assign data_arrays_1_0_MPORT_2_en = refill_one_beat & _vb_array_T_1;
  assign line_823_clock = clock;
  assign line_823_reset = reset;
  assign line_823_valid = s0_valid ^ line_823_valid_reg;
  assign line_824_clock = clock;
  assign line_824_reset = reset;
  assign line_824_valid = _refill_paddr_T ^ line_824_valid_reg;
  assign line_825_clock = clock;
  assign line_825_reset = reset;
  assign line_825_valid = _refill_paddr_T ^ line_825_valid_reg;
  assign line_826_clock = clock;
  assign line_826_reset = reset;
  assign line_826_valid = auto_master_out_d_valid ^ line_826_valid_reg;
  assign line_827_clock = clock;
  assign line_827_reset = reset;
  assign line_827_valid = _tag_rdata_T_2 ^ line_827_valid_reg;
  assign line_828_clock = clock;
  assign line_828_reset = reset;
  assign line_828_valid = refill_done ^ line_828_valid_reg;
  assign line_829_clock = clock;
  assign line_829_reset = reset;
  assign line_829_valid = refill_one_beat ^ line_829_valid_reg;
  assign line_830_clock = clock;
  assign line_830_reset = reset;
  assign line_830_valid = io_invalidate ^ line_830_valid_reg;
  assign line_831_clock = clock;
  assign line_831_reset = reset;
  assign line_831_valid = _T_9 ^ line_831_valid_reg;
  assign line_832_clock = clock;
  assign line_832_reset = reset;
  assign line_832_valid = wen ^ line_832_valid_reg;
  assign line_833_clock = clock;
  assign line_833_reset = reset;
  assign line_833_valid = _dout_T_1 ^ line_833_valid_reg;
  assign line_834_clock = clock;
  assign line_834_reset = reset;
  assign line_834_valid = _T_14 ^ line_834_valid_reg;
  assign line_835_clock = clock;
  assign line_835_reset = reset;
  assign line_835_valid = wen ^ line_835_valid_reg;
  assign line_836_clock = clock;
  assign line_836_reset = reset;
  assign line_836_valid = _dout_T_5 ^ line_836_valid_reg;
  assign line_837_clock = clock;
  assign line_837_reset = reset;
  assign line_837_valid = io_s1_paddr[2] ^ line_837_valid_reg;
  assign line_838_clock = clock;
  assign line_838_reset = reset;
  assign line_838_valid = s1_valid ^ line_838_valid_reg;
  assign line_839_clock = clock;
  assign line_839_reset = reset;
  assign line_839_valid = s1_valid ^ line_839_valid_reg;
  assign line_840_clock = clock;
  assign line_840_reset = reset;
  assign line_840_valid = s1_valid ^ line_840_valid_reg;
  assign line_841_clock = clock;
  assign line_841_reset = reset;
  assign line_841_valid = s1_valid ^ line_841_valid_reg;
  assign line_842_clock = clock;
  assign line_842_reset = reset;
  assign line_842_valid = s1_valid ^ line_842_valid_reg;
  assign line_843_clock = clock;
  assign line_843_reset = reset;
  assign line_843_valid = _T_9 ^ line_843_valid_reg;
  assign line_844_clock = clock;
  assign line_844_reset = reset;
  assign line_844_valid = _T_25 ^ line_844_valid_reg;
  assign line_845_clock = clock;
  assign line_845_reset = reset;
  assign line_845_valid = refill_fire ^ line_845_valid_reg;
  assign line_846_clock = clock;
  assign line_846_reset = reset;
  assign line_846_valid = refill_done ^ line_846_valid_reg;
  assign auto_master_out_a_valid = s2_miss & s2_request_refill_REG; // @[src/main/scala/rocket/ICache.scala 377:35]
  assign auto_master_out_a_bits_address = {refill_paddr[31:5], 5'h0}; // @[src/main/scala/rocket/ICache.scala 761:64]
  assign io_req_ready = ~refill_one_beat; // @[src/main/scala/rocket/ICache.scala 386:19]
  assign io_resp_valid = s2_valid & s2_hit; // @[src/main/scala/rocket/ICache.scala 651:33]
  assign io_resp_bits_data = s2_dout_0; // @[src/main/scala/rocket/ICache.scala 648:25]
  assign io_resp_bits_ae = s2_tl_error; // @[src/main/scala/rocket/ICache.scala 649:23]
  always @(posedge clock) begin
    if (tag_array_0_MPORT_en & tag_array_0_MPORT_mask) begin
      tag_array_0[tag_array_0_MPORT_addr] <= tag_array_0_MPORT_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    tag_array_0_tag_rdata_en_pipe_0 <= _tag_rdata_T_1 & s0_valid;
    if (_tag_rdata_T_1 & s0_valid) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= io_req_bits_addr[5];
    end
    if (data_arrays_0_0_MPORT_1_en & data_arrays_0_0_MPORT_1_mask) begin
      data_arrays_0_0[data_arrays_0_0_MPORT_1_addr] <= data_arrays_0_0_MPORT_1_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_0_0_dout_en_pipe_0 <= _dout_T & s0_ren;
    if (_dout_T & s0_ren) begin
      if (refill_one_beat) begin
        data_arrays_0_0_dout_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_0_0_dout_addr_pipe_0 <= io_req_bits_addr[5:3];
      end
    end
    if (data_arrays_1_0_MPORT_2_en & data_arrays_1_0_MPORT_2_mask) begin
      data_arrays_1_0[data_arrays_1_0_MPORT_2_addr] <= data_arrays_1_0_MPORT_2_data; // @[src/main/scala/util/DescribedSRAM.scala 17:26]
    end
    data_arrays_1_0_dout_1_en_pipe_0 <= _dout_T & s0_ren_1;
    if (_dout_T & s0_ren_1) begin
      if (refill_one_beat) begin
        data_arrays_1_0_dout_1_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_1_0_dout_1_addr_pipe_0 <= io_req_bits_addr[5:3];
      end
    end
    if (reset) begin // @[src/main/scala/rocket/ICache.scala 333:25]
      s1_valid <= 1'h0; // @[src/main/scala/rocket/ICache.scala 333:25]
    end else begin
      s1_valid <= s0_valid; // @[src/main/scala/rocket/ICache.scala 387:12]
    end
    line_823_valid_reg <= s0_valid;
    vb_array <= _GEN_86[1:0]; // @[src/main/scala/rocket/ICache.scala 440:{25,25}]
    if (reset) begin // @[src/main/scala/rocket/ICache.scala 355:25]
      s2_valid <= 1'h0; // @[src/main/scala/rocket/ICache.scala 355:25]
    end else begin
      s2_valid <= s1_valid & ~io_s1_kill; // @[src/main/scala/rocket/ICache.scala 355:25]
    end
    s2_hit <= _s1_tag_hit_0_T; // @[src/main/scala/rocket/ICache.scala 356:23]
    if (~refill_valid) begin // @[src/main/scala/rocket/ICache.scala 821:24]
      invalidated <= 1'h0; // @[src/main/scala/rocket/ICache.scala 821:38]
    end else begin
      invalidated <= _GEN_48;
    end
    if (reset) begin // @[src/main/scala/rocket/ICache.scala 360:29]
      refill_valid <= 1'h0; // @[src/main/scala/rocket/ICache.scala 360:29]
    end else if (refill_done) begin // @[src/main/scala/rocket/ICache.scala 823:22]
      refill_valid <= 1'h0; // @[src/main/scala/rocket/ICache.scala 823:37]
    end else begin
      refill_valid <= _GEN_80;
    end
    s2_request_refill_REG <= ~(s2_miss | refill_valid); // @[src/main/scala/rocket/ICache.scala 372:31]
    if (s1_valid & s1_can_request_refill) begin // @[src/main/scala/rocket/ICache.scala 378:31]
      refill_paddr <= io_s1_paddr; // @[src/main/scala/rocket/ICache.scala 378:31]
    end
    line_824_valid_reg <= _refill_paddr_T;
    line_825_valid_reg <= _refill_paddr_T;
    if (reset) begin // @[src/main/scala/tilelink/Edges.scala 229:27]
      counter <= 2'h0; // @[src/main/scala/tilelink/Edges.scala 229:27]
    end else if (auto_master_out_d_valid) begin // @[src/main/scala/tilelink/Edges.scala 235:17]
      if (first) begin // @[src/main/scala/tilelink/Edges.scala 236:21]
        if (refill_one_beat_opdata) begin // @[src/main/scala/tilelink/Edges.scala 221:14]
          counter <= beats1_decode;
        end else begin
          counter <= 2'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    line_826_valid_reg <= auto_master_out_d_valid;
    line_827_valid_reg <= _tag_rdata_T_2;
    if (refill_one_beat) begin // @[src/main/scala/rocket/ICache.scala 441:26]
      accruedRefillError <= refillError; // @[src/main/scala/rocket/ICache.scala 442:24]
    end
    line_828_valid_reg <= refill_done;
    line_829_valid_reg <= refill_one_beat;
    line_830_valid_reg <= io_invalidate;
    line_831_valid_reg <= _T_9;
    line_832_valid_reg <= wen;
    line_833_valid_reg <= _dout_T_1;
    line_834_valid_reg <= _T_14;
    line_835_valid_reg <= wen;
    line_836_valid_reg <= _dout_T_5;
    line_837_valid_reg <= io_s1_paddr[2];
    line_838_valid_reg <= s1_valid;
    if (s1_valid) begin // @[src/main/scala/rocket/ICache.scala 604:26]
      if (io_s1_paddr[2]) begin // @[src/main/scala/rocket/ICache.scala 584:71]
        s2_dout_0 <= data_arrays_1_0_dout_1_data; // @[src/main/scala/rocket/ICache.scala 585:15]
      end else begin
        s2_dout_0 <= _GEN_60;
      end
    end
    line_839_valid_reg <= s1_valid;
    line_840_valid_reg <= s1_valid;
    if (s1_valid) begin // @[src/main/scala/rocket/ICache.scala 607:30]
      s2_tl_error <= |s1_tl_error_0; // @[src/main/scala/rocket/ICache.scala 607:30]
    end
    line_841_valid_reg <= s1_valid;
    line_842_valid_reg <= s1_valid;
    line_843_valid_reg <= _T_9;
    line_844_valid_reg <= _T_25;
    line_845_valid_reg <= refill_fire;
    line_846_valid_reg <= refill_done;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[26:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_3[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    data_arrays_1_0[initvar] = _RAND_6[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_tag_rdata_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_tag_rdata_addr_pipe_0 = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  data_arrays_0_0_dout_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data_arrays_0_0_dout_addr_pipe_0 = _RAND_5[2:0];
  _RAND_7 = {1{`RANDOM}};
  data_arrays_1_0_dout_1_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  data_arrays_1_0_dout_1_addr_pipe_0 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  s1_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_823_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vb_array = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  s2_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  s2_hit = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  invalidated = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  refill_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  s2_request_refill_REG = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  refill_paddr = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  line_824_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_825_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  counter = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  line_826_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  line_827_valid_reg = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  accruedRefillError = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_828_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_829_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  line_830_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  line_831_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  line_832_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  line_833_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_834_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_835_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_836_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_837_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_838_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  s2_dout_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  line_839_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_840_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  s2_tl_error = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_841_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_842_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_843_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_844_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_845_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_846_valid_reg = _RAND_44[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/rocket/ICache.scala 513:9]
    end
    //
    if (_T_9) begin
      assert(1'h1); // @[src/main/scala/rocket/ICache.scala 818:9]
    end
  end
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input         io_enq_valid, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input  [39:0] io_enq_bits_pc, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input  [31:0] io_enq_bits_data, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input         io_enq_bits_xcpt_pf_inst, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input         io_enq_bits_xcpt_ae_inst, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input         io_enq_bits_replay, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  input         io_deq_ready, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output        io_deq_valid, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output [39:0] io_deq_bits_pc, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output [31:0] io_deq_bits_data, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output        io_deq_bits_xcpt_pf_inst, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output        io_deq_bits_xcpt_ae_inst, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output        io_deq_bits_replay, // @[src/main/scala/util/ShiftQueue.scala 17:14]
  output [4:0]  io_mask // @[src/main/scala/util/ShiftQueue.scala 17:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  reg  valid_0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
  reg  valid_1; // @[src/main/scala/util/ShiftQueue.scala 21:30]
  reg  valid_2; // @[src/main/scala/util/ShiftQueue.scala 21:30]
  reg  valid_3; // @[src/main/scala/util/ShiftQueue.scala 21:30]
  reg  valid_4; // @[src/main/scala/util/ShiftQueue.scala 21:30]
  reg [39:0] elts_0_pc; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [31:0] elts_0_data; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_0_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_0_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_0_replay; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [39:0] elts_1_pc; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [31:0] elts_1_data; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_1_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_1_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_1_replay; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [39:0] elts_2_pc; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [31:0] elts_2_data; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_2_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_2_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_2_replay; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [39:0] elts_3_pc; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [31:0] elts_3_data; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_3_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_3_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_3_replay; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [39:0] elts_4_pc; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg [31:0] elts_4_data; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_4_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_4_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  reg  elts_4_replay; // @[src/main/scala/util/ShiftQueue.scala 22:25]
  wire  _wen_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _wen_T_2 = _wen_T & valid_0; // @[src/main/scala/util/ShiftQueue.scala 30:43]
  wire  _wen_T_3 = valid_1 | _wen_T & valid_0; // @[src/main/scala/util/ShiftQueue.scala 30:28]
  wire  _wen_T_6 = ~valid_0; // @[src/main/scala/util/ShiftQueue.scala 31:46]
  wire  _wen_T_7 = _wen_T & ~valid_0; // @[src/main/scala/util/ShiftQueue.scala 31:43]
  wire  wen = io_deq_ready ? _wen_T_3 : _wen_T_7; // @[src/main/scala/util/ShiftQueue.scala 29:10]
  wire  line_847_clock;
  wire  line_847_reset;
  wire  line_847_valid;
  reg  line_847_valid_reg;
  wire  _valid_0_T_6 = _wen_T | valid_0; // @[src/main/scala/util/ShiftQueue.scala 37:43]
  wire  _wen_T_10 = _wen_T & valid_1; // @[src/main/scala/util/ShiftQueue.scala 30:43]
  wire  _wen_T_11 = valid_2 | _wen_T & valid_1; // @[src/main/scala/util/ShiftQueue.scala 30:28]
  wire  _wen_T_15 = _wen_T_2 & ~valid_1; // @[src/main/scala/util/ShiftQueue.scala 31:43]
  wire  wen_1 = io_deq_ready ? _wen_T_11 : _wen_T_15; // @[src/main/scala/util/ShiftQueue.scala 29:10]
  wire  line_848_clock;
  wire  line_848_reset;
  wire  line_848_valid;
  reg  line_848_valid_reg;
  wire  _valid_1_T_6 = _wen_T_2 | valid_1; // @[src/main/scala/util/ShiftQueue.scala 37:43]
  wire  _wen_T_18 = _wen_T & valid_2; // @[src/main/scala/util/ShiftQueue.scala 30:43]
  wire  _wen_T_19 = valid_3 | _wen_T & valid_2; // @[src/main/scala/util/ShiftQueue.scala 30:28]
  wire  _wen_T_23 = _wen_T_10 & ~valid_2; // @[src/main/scala/util/ShiftQueue.scala 31:43]
  wire  wen_2 = io_deq_ready ? _wen_T_19 : _wen_T_23; // @[src/main/scala/util/ShiftQueue.scala 29:10]
  wire  line_849_clock;
  wire  line_849_reset;
  wire  line_849_valid;
  reg  line_849_valid_reg;
  wire  _valid_2_T_6 = _wen_T_10 | valid_2; // @[src/main/scala/util/ShiftQueue.scala 37:43]
  wire  _wen_T_26 = _wen_T & valid_3; // @[src/main/scala/util/ShiftQueue.scala 30:43]
  wire  _wen_T_27 = valid_4 | _wen_T & valid_3; // @[src/main/scala/util/ShiftQueue.scala 30:28]
  wire  _wen_T_31 = _wen_T_18 & ~valid_3; // @[src/main/scala/util/ShiftQueue.scala 31:43]
  wire  wen_3 = io_deq_ready ? _wen_T_27 : _wen_T_31; // @[src/main/scala/util/ShiftQueue.scala 29:10]
  wire  line_850_clock;
  wire  line_850_reset;
  wire  line_850_valid;
  reg  line_850_valid_reg;
  wire  _valid_3_T_6 = _wen_T_18 | valid_3; // @[src/main/scala/util/ShiftQueue.scala 37:43]
  wire  _wen_T_34 = _wen_T & valid_4; // @[src/main/scala/util/ShiftQueue.scala 30:43]
  wire  _wen_T_39 = _wen_T_26 & ~valid_4; // @[src/main/scala/util/ShiftQueue.scala 31:43]
  wire  wen_4 = io_deq_ready ? _wen_T_34 : _wen_T_39; // @[src/main/scala/util/ShiftQueue.scala 29:10]
  wire  line_851_clock;
  wire  line_851_reset;
  wire  line_851_valid;
  reg  line_851_valid_reg;
  wire  _valid_4_T_6 = _wen_T_26 | valid_4; // @[src/main/scala/util/ShiftQueue.scala 37:43]
  wire  line_852_clock;
  wire  line_852_reset;
  wire  line_852_valid;
  reg  line_852_valid_reg;
  wire  line_853_clock;
  wire  line_853_reset;
  wire  line_853_valid;
  reg  line_853_valid_reg;
  wire [1:0] io_mask_lo = {valid_1,valid_0}; // @[src/main/scala/util/ShiftQueue.scala 53:20]
  wire [2:0] io_mask_hi = {valid_4,valid_3,valid_2}; // @[src/main/scala/util/ShiftQueue.scala 53:20]
  GEN_w1_line #(.COVER_INDEX(847)) line_847 (
    .clock(line_847_clock),
    .reset(line_847_reset),
    .valid(line_847_valid)
  );
  GEN_w1_line #(.COVER_INDEX(848)) line_848 (
    .clock(line_848_clock),
    .reset(line_848_reset),
    .valid(line_848_valid)
  );
  GEN_w1_line #(.COVER_INDEX(849)) line_849 (
    .clock(line_849_clock),
    .reset(line_849_reset),
    .valid(line_849_valid)
  );
  GEN_w1_line #(.COVER_INDEX(850)) line_850 (
    .clock(line_850_clock),
    .reset(line_850_reset),
    .valid(line_850_valid)
  );
  GEN_w1_line #(.COVER_INDEX(851)) line_851 (
    .clock(line_851_clock),
    .reset(line_851_reset),
    .valid(line_851_valid)
  );
  GEN_w1_line #(.COVER_INDEX(852)) line_852 (
    .clock(line_852_clock),
    .reset(line_852_reset),
    .valid(line_852_valid)
  );
  GEN_w1_line #(.COVER_INDEX(853)) line_853 (
    .clock(line_853_clock),
    .reset(line_853_reset),
    .valid(line_853_valid)
  );
  assign line_847_clock = clock;
  assign line_847_reset = reset;
  assign line_847_valid = wen ^ line_847_valid_reg;
  assign line_848_clock = clock;
  assign line_848_reset = reset;
  assign line_848_valid = wen_1 ^ line_848_valid_reg;
  assign line_849_clock = clock;
  assign line_849_reset = reset;
  assign line_849_valid = wen_2 ^ line_849_valid_reg;
  assign line_850_clock = clock;
  assign line_850_reset = reset;
  assign line_850_valid = wen_3 ^ line_850_valid_reg;
  assign line_851_clock = clock;
  assign line_851_reset = reset;
  assign line_851_valid = wen_4 ^ line_851_valid_reg;
  assign line_852_clock = clock;
  assign line_852_reset = reset;
  assign line_852_valid = io_enq_valid ^ line_852_valid_reg;
  assign line_853_clock = clock;
  assign line_853_reset = reset;
  assign line_853_valid = _wen_T_6 ^ line_853_valid_reg;
  assign io_enq_ready = ~valid_4; // @[src/main/scala/util/ShiftQueue.scala 40:19]
  assign io_deq_valid = io_enq_valid | valid_0; // @[src/main/scala/util/ShiftQueue.scala 41:16 45:{25,40}]
  assign io_deq_bits_pc = _wen_T_6 ? io_enq_bits_pc : elts_0_pc; // @[src/main/scala/util/ShiftQueue.scala 42:15 46:{22,36}]
  assign io_deq_bits_data = _wen_T_6 ? io_enq_bits_data : elts_0_data; // @[src/main/scala/util/ShiftQueue.scala 42:15 46:{22,36}]
  assign io_deq_bits_xcpt_pf_inst = _wen_T_6 ? io_enq_bits_xcpt_pf_inst : elts_0_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 42:15 46:{22,36}]
  assign io_deq_bits_xcpt_ae_inst = _wen_T_6 ? io_enq_bits_xcpt_ae_inst : elts_0_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 42:15 46:{22,36}]
  assign io_deq_bits_replay = _wen_T_6 ? io_enq_bits_replay : elts_0_replay; // @[src/main/scala/util/ShiftQueue.scala 42:15 46:{22,36}]
  assign io_mask = {io_mask_hi,io_mask_lo}; // @[src/main/scala/util/ShiftQueue.scala 53:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/util/ShiftQueue.scala 21:30]
      valid_0 <= 1'h0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 35:10]
      valid_0 <= _wen_T_3;
    end else begin
      valid_0 <= _valid_0_T_6;
    end
    if (reset) begin // @[src/main/scala/util/ShiftQueue.scala 21:30]
      valid_1 <= 1'h0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 35:10]
      valid_1 <= _wen_T_11;
    end else begin
      valid_1 <= _valid_1_T_6;
    end
    if (reset) begin // @[src/main/scala/util/ShiftQueue.scala 21:30]
      valid_2 <= 1'h0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 35:10]
      valid_2 <= _wen_T_19;
    end else begin
      valid_2 <= _valid_2_T_6;
    end
    if (reset) begin // @[src/main/scala/util/ShiftQueue.scala 21:30]
      valid_3 <= 1'h0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 35:10]
      valid_3 <= _wen_T_27;
    end else begin
      valid_3 <= _valid_3_T_6;
    end
    if (reset) begin // @[src/main/scala/util/ShiftQueue.scala 21:30]
      valid_4 <= 1'h0; // @[src/main/scala/util/ShiftQueue.scala 21:30]
    end else if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 35:10]
      valid_4 <= _wen_T_34;
    end else begin
      valid_4 <= _valid_4_T_6;
    end
    if (wen) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_1) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_0_pc <= elts_1_pc;
      end else begin
        elts_0_pc <= io_enq_bits_pc;
      end
    end
    if (wen) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_1) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_0_data <= elts_1_data;
      end else begin
        elts_0_data <= io_enq_bits_data;
      end
    end
    if (wen) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_1) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_0_xcpt_pf_inst <= elts_1_xcpt_pf_inst;
      end else begin
        elts_0_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (wen) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_1) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_0_xcpt_ae_inst <= elts_1_xcpt_ae_inst;
      end else begin
        elts_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (wen) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_1) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_0_replay <= elts_1_replay;
      end else begin
        elts_0_replay <= io_enq_bits_replay;
      end
    end
    if (wen_1) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_2) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_1_pc <= elts_2_pc;
      end else begin
        elts_1_pc <= io_enq_bits_pc;
      end
    end
    if (wen_1) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_2) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_1_data <= elts_2_data;
      end else begin
        elts_1_data <= io_enq_bits_data;
      end
    end
    if (wen_1) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_2) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_1_xcpt_pf_inst <= elts_2_xcpt_pf_inst;
      end else begin
        elts_1_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (wen_1) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_2) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_1_xcpt_ae_inst <= elts_2_xcpt_ae_inst;
      end else begin
        elts_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (wen_1) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_2) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_1_replay <= elts_2_replay;
      end else begin
        elts_1_replay <= io_enq_bits_replay;
      end
    end
    if (wen_2) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_3) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_2_pc <= elts_3_pc;
      end else begin
        elts_2_pc <= io_enq_bits_pc;
      end
    end
    if (wen_2) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_3) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_2_data <= elts_3_data;
      end else begin
        elts_2_data <= io_enq_bits_data;
      end
    end
    if (wen_2) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_3) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_2_xcpt_pf_inst <= elts_3_xcpt_pf_inst;
      end else begin
        elts_2_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (wen_2) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_3) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_2_xcpt_ae_inst <= elts_3_xcpt_ae_inst;
      end else begin
        elts_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (wen_2) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_3) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_2_replay <= elts_3_replay;
      end else begin
        elts_2_replay <= io_enq_bits_replay;
      end
    end
    if (wen_3) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_4) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_3_pc <= elts_4_pc;
      end else begin
        elts_3_pc <= io_enq_bits_pc;
      end
    end
    if (wen_3) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_4) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_3_data <= elts_4_data;
      end else begin
        elts_3_data <= io_enq_bits_data;
      end
    end
    if (wen_3) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_4) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_3_xcpt_pf_inst <= elts_4_xcpt_pf_inst;
      end else begin
        elts_3_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (wen_3) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_4) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_3_xcpt_ae_inst <= elts_4_xcpt_ae_inst;
      end else begin
        elts_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (wen_3) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      if (valid_4) begin // @[src/main/scala/util/ShiftQueue.scala 27:57]
        elts_3_replay <= elts_4_replay;
      end else begin
        elts_3_replay <= io_enq_bits_replay;
      end
    end
    if (wen_4) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      elts_4_pc <= io_enq_bits_pc; // @[src/main/scala/util/ShiftQueue.scala 32:26]
    end
    if (wen_4) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      elts_4_data <= io_enq_bits_data; // @[src/main/scala/util/ShiftQueue.scala 32:26]
    end
    if (wen_4) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      elts_4_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst; // @[src/main/scala/util/ShiftQueue.scala 32:26]
    end
    if (wen_4) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      elts_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst; // @[src/main/scala/util/ShiftQueue.scala 32:26]
    end
    if (wen_4) begin // @[src/main/scala/util/ShiftQueue.scala 32:16]
      elts_4_replay <= io_enq_bits_replay; // @[src/main/scala/util/ShiftQueue.scala 32:26]
    end
    if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 29:10]
      line_847_valid_reg <= _wen_T_3;
    end else begin
      line_847_valid_reg <= _wen_T_7;
    end
    if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 29:10]
      line_848_valid_reg <= _wen_T_11;
    end else begin
      line_848_valid_reg <= _wen_T_15;
    end
    if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 29:10]
      line_849_valid_reg <= _wen_T_19;
    end else begin
      line_849_valid_reg <= _wen_T_23;
    end
    if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 29:10]
      line_850_valid_reg <= _wen_T_27;
    end else begin
      line_850_valid_reg <= _wen_T_31;
    end
    if (io_deq_ready) begin // @[src/main/scala/util/ShiftQueue.scala 29:10]
      line_851_valid_reg <= _wen_T_34;
    end else begin
      line_851_valid_reg <= _wen_T_39;
    end
    line_852_valid_reg <= io_enq_valid;
    line_853_valid_reg <= _wen_T_6;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_4 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  elts_0_pc = _RAND_5[39:0];
  _RAND_6 = {1{`RANDOM}};
  elts_0_data = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  elts_0_xcpt_pf_inst = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  elts_0_xcpt_ae_inst = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  elts_0_replay = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  elts_1_pc = _RAND_10[39:0];
  _RAND_11 = {1{`RANDOM}};
  elts_1_data = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  elts_1_xcpt_pf_inst = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  elts_1_xcpt_ae_inst = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  elts_1_replay = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  elts_2_pc = _RAND_15[39:0];
  _RAND_16 = {1{`RANDOM}};
  elts_2_data = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  elts_2_xcpt_pf_inst = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  elts_2_xcpt_ae_inst = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  elts_2_replay = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  elts_3_pc = _RAND_20[39:0];
  _RAND_21 = {1{`RANDOM}};
  elts_3_data = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  elts_3_xcpt_pf_inst = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  elts_3_xcpt_ae_inst = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  elts_3_replay = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  elts_4_pc = _RAND_25[39:0];
  _RAND_26 = {1{`RANDOM}};
  elts_4_data = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  elts_4_xcpt_pf_inst = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  elts_4_xcpt_ae_inst = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  elts_4_replay = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  line_847_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  line_848_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  line_849_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_850_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_851_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_852_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_853_valid_reg = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OptimizationBarrier_12(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
endmodule
module PMPChecker_2(
  input   clock,
  input   reset
);
endmodule
module OptimizationBarrier_13(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_px, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_px, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_px = io_x_px; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_14(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_px, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_px, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_px = io_x_px; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_15(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_px, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_px, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_px = io_x_px; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_16(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_px, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_c, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_px, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_c // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_px = io_x_px; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_c = io_x_c; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_17(
  input         clock,
  input         reset,
  input  [19:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_ae_final, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_pf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_gf, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_sx, // @[src/main/scala/util/package.scala 260:18]
  output [19:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_ptw, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_ae_final, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_pf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_gf, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_sx // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_ptw = io_x_ae_ptw; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_ae_final = io_x_ae_final; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_pf = io_x_pf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_gf = io_x_gf; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_sx = io_x_sx; // @[src/main/scala/util/package.scala 264:12]
endmodule
module TLB_1(
  input         clock,
  input         reset,
  output        io_req_ready, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_req_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [39:0] io_req_bits_vaddr, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [1:0]  io_req_bits_prv, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_miss, // @[src/main/scala/rocket/TLB.scala 309:14]
  output [31:0] io_resp_paddr, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_pf_inst, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_ae_inst, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_resp_cacheable, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_bits_rs1, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_sfence_bits_rs2, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [38:0] io_sfence_bits_addr, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_req_ready, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_bits_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  output [26:0] io_ptw_req_bits_bits_addr, // @[src/main/scala/rocket/TLB.scala 309:14]
  output        io_ptw_req_bits_bits_need_gpa, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_valid, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_ae_ptw, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_ae_final, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pf, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [43:0] io_ptw_resp_bits_pte_ppn, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_d, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_a, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_g, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_u, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_x, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_w, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_r, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_pte_v, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [1:0]  io_ptw_resp_bits_level, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_ptw_resp_bits_homogeneous, // @[src/main/scala/rocket/TLB.scala 309:14]
  input  [3:0]  io_ptw_ptbr_mode, // @[src/main/scala/rocket/TLB.scala 309:14]
  input         io_kill // @[src/main/scala/rocket/TLB.scala 309:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
`endif // RANDOMIZE_REG_INIT
  wire  mpu_ppn_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  mpu_ppn_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] mpu_ppn_barrier_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] mpu_ppn_barrier_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  pmp_clock; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  pmp_reset; // @[src/main/scala/rocket/TLB.scala 405:19]
  wire  entries_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_1_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_1_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_1_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_2_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_2_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_2_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_3_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_x_c; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_3_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_px; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_3_io_y_c; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_4_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_x_sx; // @[src/main/scala/util/package.scala 259:25]
  wire [19:0] entries_barrier_4_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_ae_ptw; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_ae_final; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_pf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_gf; // @[src/main/scala/util/package.scala 259:25]
  wire  entries_barrier_4_io_y_sx; // @[src/main/scala/util/package.scala 259:25]
  wire [26:0] vpn = io_req_bits_vaddr[38:12]; // @[src/main/scala/rocket/TLB.scala 324:30]
  reg [26:0] sectored_entries_0_0_tag_vpn; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_0_data_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [26:0] sectored_entries_0_1_tag_vpn; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [41:0] sectored_entries_0_1_data_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg  sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29]
  reg [1:0] superpage_entries_0_level; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [26:0] superpage_entries_0_tag_vpn; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [41:0] superpage_entries_0_data_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg  superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [1:0] superpage_entries_1_level; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [26:0] superpage_entries_1_tag_vpn; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [41:0] superpage_entries_1_data_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg  superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30]
  reg [1:0] special_entry_level; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [26:0] special_entry_tag_vpn; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [41:0] special_entry_data_0; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg  special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 335:56]
  reg [1:0] state; // @[src/main/scala/rocket/TLB.scala 341:22]
  reg [26:0] r_refill_tag; // @[src/main/scala/rocket/TLB.scala 343:25]
  reg  r_superpage_repl_addr; // @[src/main/scala/rocket/TLB.scala 344:34]
  reg  r_sectored_repl_addr; // @[src/main/scala/rocket/TLB.scala 345:33]
  reg  r_sectored_hit_valid; // @[src/main/scala/rocket/TLB.scala 346:27]
  reg  r_sectored_hit_bits; // @[src/main/scala/rocket/TLB.scala 346:27]
  reg  r_need_gpa; // @[src/main/scala/rocket/TLB.scala 350:23]
  wire  priv_s = io_req_bits_prv[0]; // @[src/main/scala/rocket/TLB.scala 359:20]
  wire  priv_uses_vm = io_req_bits_prv <= 2'h1; // @[src/main/scala/rocket/TLB.scala 361:27]
  wire  stage1_en = io_ptw_ptbr_mode[3]; // @[src/main/scala/rocket/TLB.scala 363:41]
  wire  vm_enabled = stage1_en & priv_uses_vm; // @[src/main/scala/rocket/TLB.scala 388:45]
  wire [19:0] refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[src/main/scala/rocket/TLB.scala 395:44]
  wire  _invalidate_refill_T = state == 2'h1; // @[src/main/scala/util/package.scala 16:47]
  wire  _invalidate_refill_T_1 = state == 2'h3; // @[src/main/scala/util/package.scala 16:47]
  wire  _invalidate_refill_T_2 = _invalidate_refill_T | _invalidate_refill_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  invalidate_refill = _invalidate_refill_T_2 | io_sfence_valid; // @[src/main/scala/rocket/TLB.scala 399:88]
  wire [1:0] mpu_ppn_res = mpu_ppn_barrier_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire  mpu_ppn_ignore = special_entry_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 187:28]
  wire [26:0] _mpu_ppn_T_24 = mpu_ppn_ignore ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_488 = {{7'd0}, mpu_ppn_barrier_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _mpu_ppn_T_25 = _mpu_ppn_T_24 | _GEN_488; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire  mpu_ppn_ignore_1 = special_entry_level < 2'h2; // @[src/main/scala/rocket/TLB.scala 187:28]
  wire [26:0] _mpu_ppn_T_28 = mpu_ppn_ignore_1 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _mpu_ppn_T_29 = _mpu_ppn_T_28 | _GEN_488; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _mpu_ppn_T_31 = {mpu_ppn_res,_mpu_ppn_T_25[17:9],_mpu_ppn_T_29[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [27:0] _mpu_ppn_T_33 = vm_enabled ? {{8'd0}, _mpu_ppn_T_31} : io_req_bits_vaddr[39:12]; // @[src/main/scala/rocket/TLB.scala 402:20]
  wire [27:0] mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _mpu_ppn_T_33; // @[src/main/scala/rocket/TLB.scala 401:20]
  wire [39:0] mpu_physaddr = {mpu_ppn,io_req_bits_vaddr[11:0]}; // @[src/main/scala/rocket/TLB.scala 403:25]
  wire [39:0] _legal_address_T = mpu_physaddr ^ 40'h10000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [40:0] _legal_address_T_1 = {1'b0,$signed(_legal_address_T)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [40:0] _legal_address_T_3 = $signed(_legal_address_T_1) & -41'sh10000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _legal_address_T_4 = $signed(_legal_address_T_3) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire [39:0] _legal_address_T_5 = mpu_physaddr ^ 40'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [40:0] _legal_address_T_6 = {1'b0,$signed(_legal_address_T_5)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [40:0] _legal_address_T_8 = $signed(_legal_address_T_6) & -41'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _legal_address_T_9 = $signed(_legal_address_T_8) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire  legal_address = _legal_address_T_4 | _legal_address_T_9; // @[src/main/scala/rocket/TLB.scala 412:67]
  wire [40:0] _cacheable_T_8 = $signed(_legal_address_T_6) & 41'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _cacheable_T_9 = $signed(_cacheable_T_8) == 41'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire  cacheable = legal_address & _cacheable_T_9; // @[src/main/scala/rocket/TLB.scala 415:19]
  wire  _sector_hits_T_2 = sectored_entries_0_0_valid_0 | sectored_entries_0_0_valid_1 | sectored_entries_0_0_valid_2 |
    sectored_entries_0_0_valid_3; // @[src/main/scala/util/package.scala 73:59]
  wire [26:0] _sector_hits_T_3 = sectored_entries_0_0_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 164:61]
  wire  _sector_hits_T_5 = _sector_hits_T_3[26:2] == 25'h0; // @[src/main/scala/rocket/TLB.scala 164:86]
  wire  sector_hits_0 = _sector_hits_T_2 & _sector_hits_T_5; // @[src/main/scala/rocket/TLB.scala 162:55]
  wire  _sector_hits_T_10 = sectored_entries_0_1_valid_0 | sectored_entries_0_1_valid_1 | sectored_entries_0_1_valid_2
     | sectored_entries_0_1_valid_3; // @[src/main/scala/util/package.scala 73:59]
  wire [26:0] _sector_hits_T_11 = sectored_entries_0_1_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 164:61]
  wire  _sector_hits_T_13 = _sector_hits_T_11[26:2] == 25'h0; // @[src/main/scala/rocket/TLB.scala 164:86]
  wire  sector_hits_1 = _sector_hits_T_10 & _sector_hits_T_13; // @[src/main/scala/rocket/TLB.scala 162:55]
  wire [26:0] _superpage_hits_T = superpage_entries_0_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  superpage_hits_ignore_1 = superpage_entries_0_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 172:28]
  wire  superpage_hits_0 = superpage_entries_0_valid_0 & _superpage_hits_T[26:18] == 9'h0 & (superpage_hits_ignore_1 |
    _superpage_hits_T[17:9] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire [26:0] _superpage_hits_T_14 = superpage_entries_1_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  superpage_hits_ignore_4 = superpage_entries_1_level < 2'h1; // @[src/main/scala/rocket/TLB.scala 172:28]
  wire  superpage_hits_1 = superpage_entries_1_valid_0 & _superpage_hits_T_14[26:18] == 9'h0 & (superpage_hits_ignore_4
     | _superpage_hits_T_14[17:9] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire [1:0] hitsVec_idx = vpn[1:0]; // @[src/main/scala/util/package.scala 155:13]
  wire  _GEN_0 = 2'h0 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_854_clock;
  wire  line_854_reset;
  wire  line_854_valid;
  reg  line_854_valid_reg;
  wire  _GEN_1 = 2'h1 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_855_clock;
  wire  line_855_reset;
  wire  line_855_valid;
  reg  line_855_valid_reg;
  wire  _GEN_146 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_valid_1 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _GEN_2 = 2'h2 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_856_clock;
  wire  line_856_reset;
  wire  line_856_valid;
  reg  line_856_valid_reg;
  wire  _GEN_147 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_valid_2 : _GEN_146; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _GEN_3 = 2'h3 == hitsVec_idx; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  line_857_clock;
  wire  line_857_reset;
  wire  line_857_valid;
  reg  line_857_valid_reg;
  wire  _GEN_148 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_valid_3 : _GEN_147; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _hitsVec_T_5 = _GEN_148 & _sector_hits_T_5; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  hitsVec_0 = vm_enabled & _hitsVec_T_5; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  line_858_clock;
  wire  line_858_reset;
  wire  line_858_valid;
  reg  line_858_valid_reg;
  wire  line_859_clock;
  wire  line_859_reset;
  wire  line_859_valid;
  reg  line_859_valid_reg;
  wire  _GEN_150 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_valid_1 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  line_860_clock;
  wire  line_860_reset;
  wire  line_860_valid;
  reg  line_860_valid_reg;
  wire  _GEN_151 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_valid_2 : _GEN_150; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  line_861_clock;
  wire  line_861_reset;
  wire  line_861_valid;
  reg  line_861_valid_reg;
  wire  _GEN_152 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_valid_3 : _GEN_151; // @[src/main/scala/rocket/TLB.scala 178:{18,18}]
  wire  _hitsVec_T_11 = _GEN_152 & _sector_hits_T_13; // @[src/main/scala/rocket/TLB.scala 178:18]
  wire  hitsVec_1 = vm_enabled & _hitsVec_T_11; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  hitsVec_2 = vm_enabled & superpage_hits_0; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire  hitsVec_3 = vm_enabled & superpage_hits_1; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire [26:0] _hitsVec_T_42 = special_entry_tag_vpn ^ vpn; // @[src/main/scala/rocket/TLB.scala 173:52]
  wire  _hitsVec_T_56 = special_entry_valid_0 & _hitsVec_T_42[26:18] == 9'h0 & (mpu_ppn_ignore | _hitsVec_T_42[17:9] == 9'h0
    ) & (mpu_ppn_ignore_1 | _hitsVec_T_42[8:0] == 9'h0); // @[src/main/scala/rocket/TLB.scala 173:29]
  wire  hitsVec_4 = vm_enabled & _hitsVec_T_56; // @[src/main/scala/rocket/TLB.scala 432:44]
  wire [4:0] real_hits = {hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[src/main/scala/util/package.scala 37:27]
  wire  _hits_T = ~vm_enabled; // @[src/main/scala/rocket/TLB.scala 434:18]
  wire [5:0] hits = {_hits_T,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[src/main/scala/rocket/TLB.scala 434:17]
  wire  line_862_clock;
  wire  line_862_reset;
  wire  line_862_valid;
  reg  line_862_valid_reg;
  wire  newEntry_g = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/TLB.scala 445:25]
  wire  _newEntry_sr_T_4 = io_ptw_resp_bits_pte_v & (io_ptw_resp_bits_pte_r | io_ptw_resp_bits_pte_x & ~
    io_ptw_resp_bits_pte_w) & io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/PTW.scala 141:52]
  wire  newEntry_sr = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/PTW.scala 149:35]
  wire  newEntry_sw = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_w & io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/PTW.scala 151:40]
  wire  newEntry_sx = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/PTW.scala 153:35]
  wire  _T = ~io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/TLB.scala 466:39]
  wire  line_863_clock;
  wire  line_863_reset;
  wire  line_863_valid;
  reg  line_863_valid_reg;
  wire [10:0] special_entry_data_0_lo = {2'h3,cacheable,legal_address,legal_address,cacheable,3'h0,cacheable,1'h0}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire [5:0] special_entry_data_0_hi_lo = {io_ptw_resp_bits_pf,1'h0,newEntry_sw,newEntry_sx,newEntry_sr,1'h1}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire [41:0] _special_entry_data_0_T = {refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae_ptw,
    io_ptw_resp_bits_ae_final,1'h0,special_entry_data_0_hi_lo,special_entry_data_0_lo}; // @[src/main/scala/rocket/TLB.scala 207:24]
  wire  line_864_clock;
  wire  line_864_reset;
  wire  line_864_valid;
  reg  line_864_valid_reg;
  wire  _T_2 = io_ptw_resp_bits_level < 2'h2; // @[src/main/scala/rocket/TLB.scala 468:40]
  wire  line_865_clock;
  wire  line_865_reset;
  wire  line_865_valid;
  reg  line_865_valid_reg;
  wire  _T_3 = ~r_superpage_repl_addr; // @[src/main/scala/rocket/TLB.scala 470:82]
  wire  line_866_clock;
  wire  line_866_reset;
  wire  line_866_valid;
  reg  line_866_valid_reg;
  wire  line_867_clock;
  wire  line_867_reset;
  wire  line_867_valid;
  reg  line_867_valid_reg;
  wire  _GEN_153 = invalidate_refill ? 1'h0 : 1'h1; // @[src/main/scala/rocket/TLB.scala 206:16 472:34 210:46]
  wire  _GEN_157 = ~r_superpage_repl_addr ? _GEN_153 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 470:91]
  wire  line_868_clock;
  wire  line_868_reset;
  wire  line_868_valid;
  reg  line_868_valid_reg;
  wire  line_869_clock;
  wire  line_869_reset;
  wire  line_869_valid;
  reg  line_869_valid_reg;
  wire  _GEN_162 = r_superpage_repl_addr ? _GEN_153 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 470:91]
  wire  line_870_clock;
  wire  line_870_reset;
  wire  line_870_valid;
  reg  line_870_valid_reg;
  wire  waddr_1 = r_sectored_hit_valid ? r_sectored_hit_bits : r_sectored_repl_addr; // @[src/main/scala/rocket/TLB.scala 477:22]
  wire  _T_5 = ~waddr_1; // @[src/main/scala/rocket/TLB.scala 478:75]
  wire  line_871_clock;
  wire  line_871_reset;
  wire  line_871_valid;
  reg  line_871_valid_reg;
  wire  _T_6 = ~r_sectored_hit_valid; // @[src/main/scala/rocket/TLB.scala 479:15]
  wire  line_872_clock;
  wire  line_872_reset;
  wire  line_872_valid;
  reg  line_872_valid_reg;
  wire  _GEN_164 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_165 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_166 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_167 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire [1:0] idx = r_refill_tag[1:0]; // @[src/main/scala/util/package.scala 155:13]
  wire  line_873_clock;
  wire  line_873_reset;
  wire  line_873_valid;
  reg  line_873_valid_reg;
  wire  _GEN_168 = 2'h0 == idx | _GEN_164; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_874_clock;
  wire  line_874_reset;
  wire  line_874_valid;
  reg  line_874_valid_reg;
  wire  _GEN_169 = 2'h1 == idx | _GEN_165; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_875_clock;
  wire  line_875_reset;
  wire  line_875_valid;
  reg  line_875_valid_reg;
  wire  _GEN_170 = 2'h2 == idx | _GEN_166; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_876_clock;
  wire  line_876_reset;
  wire  line_876_valid;
  reg  line_876_valid_reg;
  wire  _GEN_171 = 2'h3 == idx | _GEN_167; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_877_clock;
  wire  line_877_reset;
  wire  line_877_valid;
  reg  line_877_valid_reg;
  wire [41:0] _GEN_172 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_878_clock;
  wire  line_878_reset;
  wire  line_878_valid;
  reg  line_878_valid_reg;
  wire [41:0] _GEN_173 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_1; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_879_clock;
  wire  line_879_reset;
  wire  line_879_valid;
  reg  line_879_valid_reg;
  wire [41:0] _GEN_174 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_2; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_880_clock;
  wire  line_880_reset;
  wire  line_880_valid;
  reg  line_880_valid_reg;
  wire [41:0] _GEN_175 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_0_0_data_3; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_881_clock;
  wire  line_881_reset;
  wire  line_881_valid;
  reg  line_881_valid_reg;
  wire  _GEN_176 = invalidate_refill ? 1'h0 : _GEN_168; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_177 = invalidate_refill ? 1'h0 : _GEN_169; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_178 = invalidate_refill ? 1'h0 : _GEN_170; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_179 = invalidate_refill ? 1'h0 : _GEN_171; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_180 = ~waddr_1 ? _GEN_176 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_181 = ~waddr_1 ? _GEN_177 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_182 = ~waddr_1 ? _GEN_178 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_183 = ~waddr_1 ? _GEN_179 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  line_882_clock;
  wire  line_882_reset;
  wire  line_882_valid;
  reg  line_882_valid_reg;
  wire  line_883_clock;
  wire  line_883_reset;
  wire  line_883_valid;
  reg  line_883_valid_reg;
  wire  _GEN_191 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_192 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_193 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  _GEN_194 = ~r_sectored_hit_valid ? 1'h0 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 479:38 210:46 328:29]
  wire  line_884_clock;
  wire  line_884_reset;
  wire  line_884_valid;
  reg  line_884_valid_reg;
  wire  _GEN_195 = 2'h0 == idx | _GEN_191; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_885_clock;
  wire  line_885_reset;
  wire  line_885_valid;
  reg  line_885_valid_reg;
  wire  _GEN_196 = 2'h1 == idx | _GEN_192; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_886_clock;
  wire  line_886_reset;
  wire  line_886_valid;
  reg  line_886_valid_reg;
  wire  _GEN_197 = 2'h2 == idx | _GEN_193; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_887_clock;
  wire  line_887_reset;
  wire  line_887_valid;
  reg  line_887_valid_reg;
  wire  _GEN_198 = 2'h3 == idx | _GEN_194; // @[src/main/scala/rocket/TLB.scala 206:{16,16}]
  wire  line_888_clock;
  wire  line_888_reset;
  wire  line_888_valid;
  reg  line_888_valid_reg;
  wire [41:0] _GEN_199 = 2'h0 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_889_clock;
  wire  line_889_reset;
  wire  line_889_valid;
  reg  line_889_valid_reg;
  wire [41:0] _GEN_200 = 2'h1 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_1; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_890_clock;
  wire  line_890_reset;
  wire  line_890_valid;
  reg  line_890_valid_reg;
  wire [41:0] _GEN_201 = 2'h2 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_2; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_891_clock;
  wire  line_891_reset;
  wire  line_891_valid;
  reg  line_891_valid_reg;
  wire [41:0] _GEN_202 = 2'h3 == idx ? _special_entry_data_0_T : sectored_entries_0_1_data_3; // @[src/main/scala/rocket/TLB.scala 207:{15,15} 328:29]
  wire  line_892_clock;
  wire  line_892_reset;
  wire  line_892_valid;
  reg  line_892_valid_reg;
  wire  _GEN_203 = invalidate_refill ? 1'h0 : _GEN_195; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_204 = invalidate_refill ? 1'h0 : _GEN_196; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_205 = invalidate_refill ? 1'h0 : _GEN_197; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_206 = invalidate_refill ? 1'h0 : _GEN_198; // @[src/main/scala/rocket/TLB.scala 481:34 210:46]
  wire  _GEN_207 = waddr_1 ? _GEN_203 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_208 = waddr_1 ? _GEN_204 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_209 = waddr_1 ? _GEN_205 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_210 = waddr_1 ? _GEN_206 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 328:29 478:84]
  wire  _GEN_221 = io_ptw_resp_bits_level < 2'h2 ? _GEN_157 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 468:58]
  wire  _GEN_226 = io_ptw_resp_bits_level < 2'h2 ? _GEN_162 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 330:30 468:58]
  wire  _GEN_228 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_0 : _GEN_180; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_229 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_1 : _GEN_181; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_230 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_2 : _GEN_182; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_231 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_0_valid_3 : _GEN_183; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_239 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_0 : _GEN_207; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_240 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_1 : _GEN_208; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_241 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_2 : _GEN_209; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_242 = io_ptw_resp_bits_level < 2'h2 ? sectored_entries_0_1_valid_3 : _GEN_210; // @[src/main/scala/rocket/TLB.scala 328:29 468:58]
  wire  _GEN_253 = ~io_ptw_resp_bits_homogeneous | special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 206:16 335:56 466:70]
  wire  _GEN_258 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_0_valid_0 : _GEN_221; // @[src/main/scala/rocket/TLB.scala 330:30 466:70]
  wire  _GEN_263 = ~io_ptw_resp_bits_homogeneous ? superpage_entries_1_valid_0 : _GEN_226; // @[src/main/scala/rocket/TLB.scala 330:30 466:70]
  wire  _GEN_265 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_0 : _GEN_228; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_266 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_1 : _GEN_229; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_267 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_2 : _GEN_230; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_268 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_0_valid_3 : _GEN_231; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_276 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_0 : _GEN_239; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_277 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_1 : _GEN_240; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_278 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_2 : _GEN_241; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_279 = ~io_ptw_resp_bits_homogeneous ? sectored_entries_0_1_valid_3 : _GEN_242; // @[src/main/scala/rocket/TLB.scala 328:29 466:70]
  wire  _GEN_290 = io_ptw_resp_valid ? _GEN_253 : special_entry_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 335:56]
  wire  _GEN_295 = io_ptw_resp_valid ? _GEN_258 : superpage_entries_0_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 330:30]
  wire  _GEN_300 = io_ptw_resp_valid ? _GEN_263 : superpage_entries_1_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 330:30]
  wire  _GEN_302 = io_ptw_resp_valid ? _GEN_265 : sectored_entries_0_0_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_303 = io_ptw_resp_valid ? _GEN_266 : sectored_entries_0_0_valid_1; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_304 = io_ptw_resp_valid ? _GEN_267 : sectored_entries_0_0_valid_2; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_305 = io_ptw_resp_valid ? _GEN_268 : sectored_entries_0_0_valid_3; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_313 = io_ptw_resp_valid ? _GEN_276 : sectored_entries_0_1_valid_0; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_314 = io_ptw_resp_valid ? _GEN_277 : sectored_entries_0_1_valid_1; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_315 = io_ptw_resp_valid ? _GEN_278 : sectored_entries_0_1_valid_2; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  _GEN_316 = io_ptw_resp_valid ? _GEN_279 : sectored_entries_0_1_valid_3; // @[src/main/scala/rocket/TLB.scala 438:20 328:29]
  wire  line_893_clock;
  wire  line_893_reset;
  wire  line_893_valid;
  reg  line_893_valid_reg;
  wire  line_894_clock;
  wire  line_894_reset;
  wire  line_894_valid;
  reg  line_894_valid_reg;
  wire [41:0] _GEN_328 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_data_1 : sectored_entries_0_0_data_0; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_895_clock;
  wire  line_895_reset;
  wire  line_895_valid;
  reg  line_895_valid_reg;
  wire [41:0] _GEN_329 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_data_2 : _GEN_328; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_896_clock;
  wire  line_896_reset;
  wire  line_896_valid;
  reg  line_896_valid_reg;
  wire [41:0] _GEN_330 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_data_3 : _GEN_329; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_897_clock;
  wire  line_897_reset;
  wire  line_897_valid;
  reg  line_897_valid_reg;
  wire  line_898_clock;
  wire  line_898_reset;
  wire  line_898_valid;
  reg  line_898_valid_reg;
  wire [41:0] _GEN_332 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_data_1 : sectored_entries_0_1_data_0; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_899_clock;
  wire  line_899_reset;
  wire  line_899_valid;
  reg  line_899_valid_reg;
  wire [41:0] _GEN_333 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_data_2 : _GEN_332; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire  line_900_clock;
  wire  line_900_reset;
  wire  line_900_valid;
  reg  line_900_valid_reg;
  wire [41:0] _GEN_334 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_data_3 : _GEN_333; // @[src/main/scala/rocket/TLB.scala 160:{77,77}]
  wire [1:0] ppn_res = entries_barrier_2_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _ppn_T_1 = superpage_hits_ignore_1 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_498 = {{7'd0}, entries_barrier_2_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_2 = _ppn_T_1 | _GEN_498; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_6 = vpn | _GEN_498; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_8 = {ppn_res,_ppn_T_2[17:9],_ppn_T_6[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [1:0] ppn_res_1 = entries_barrier_3_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _ppn_T_9 = superpage_hits_ignore_4 ? vpn : 27'h0; // @[src/main/scala/rocket/TLB.scala 188:28]
  wire [26:0] _GEN_500 = {{7'd0}, entries_barrier_3_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_10 = _ppn_T_9 | _GEN_500; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_14 = vpn | _GEN_500; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_16 = {ppn_res_1,_ppn_T_10[17:9],_ppn_T_14[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [1:0] ppn_res_2 = entries_barrier_4_io_y_ppn[19:18]; // @[src/main/scala/rocket/TLB.scala 185:26]
  wire [26:0] _GEN_502 = {{7'd0}, entries_barrier_4_io_y_ppn}; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_18 = _mpu_ppn_T_24 | _GEN_502; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [26:0] _ppn_T_22 = _mpu_ppn_T_28 | _GEN_502; // @[src/main/scala/rocket/TLB.scala 188:47]
  wire [19:0] _ppn_T_24 = {ppn_res_2,_ppn_T_18[17:9],_ppn_T_22[8:0]}; // @[src/main/scala/rocket/TLB.scala 188:18]
  wire [19:0] _ppn_T_26 = hitsVec_0 ? entries_barrier_io_y_ppn : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_27 = hitsVec_1 ? entries_barrier_1_io_y_ppn : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_28 = hitsVec_2 ? _ppn_T_8 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_29 = hitsVec_3 ? _ppn_T_16 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_30 = hitsVec_4 ? _ppn_T_24 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_31 = _hits_T ? vpn[19:0] : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_32 = _ppn_T_26 | _ppn_T_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_33 = _ppn_T_32 | _ppn_T_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_34 = _ppn_T_33 | _ppn_T_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _ppn_T_35 = _ppn_T_34 | _ppn_T_30; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] ppn = _ppn_T_35 | _ppn_T_31; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [5:0] ptw_ae_array = {1'h0,entries_barrier_4_io_y_ae_ptw,entries_barrier_3_io_y_ae_ptw,
    entries_barrier_2_io_y_ae_ptw,entries_barrier_1_io_y_ae_ptw,entries_barrier_io_y_ae_ptw}; // @[src/main/scala/rocket/TLB.scala 498:25]
  wire [5:0] final_ae_array = {1'h0,entries_barrier_4_io_y_ae_final,entries_barrier_3_io_y_ae_final,
    entries_barrier_2_io_y_ae_final,entries_barrier_1_io_y_ae_final,entries_barrier_io_y_ae_final}; // @[src/main/scala/rocket/TLB.scala 499:27]
  wire [5:0] ptw_pf_array = {1'h0,entries_barrier_4_io_y_pf,entries_barrier_3_io_y_pf,entries_barrier_2_io_y_pf,
    entries_barrier_1_io_y_pf,entries_barrier_io_y_pf}; // @[src/main/scala/rocket/TLB.scala 500:25]
  wire [5:0] ptw_gf_array = {1'h0,entries_barrier_4_io_y_gf,entries_barrier_3_io_y_gf,entries_barrier_2_io_y_gf,
    entries_barrier_1_io_y_gf,entries_barrier_io_y_gf}; // @[src/main/scala/rocket/TLB.scala 501:25]
  wire [4:0] _priv_rw_ok_T_2 = {entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,
    entries_barrier_1_io_y_u,entries_barrier_io_y_u}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _priv_rw_ok_T_5 = ~_priv_rw_ok_T_2; // @[src/main/scala/rocket/TLB.scala 505:84]
  wire [4:0] priv_x_ok = priv_s ? _priv_rw_ok_T_5 : _priv_rw_ok_T_2; // @[src/main/scala/rocket/TLB.scala 508:22]
  wire [4:0] _r_array_T_1 = {entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,
    entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; // @[src/main/scala/util/package.scala 37:27]
  wire [4:0] _x_array_T_1 = priv_x_ok & _r_array_T_1; // @[src/main/scala/rocket/TLB.scala 514:40]
  wire [5:0] x_array = {1'h1,_x_array_T_1}; // @[src/main/scala/rocket/TLB.scala 514:20]
  wire [1:0] _pr_array_T = legal_address ? 2'h3 : 2'h0; // @[src/main/scala/rocket/TLB.scala 521:26]
  wire [5:0] _pr_array_T_3 = ptw_ae_array | final_ae_array; // @[src/main/scala/rocket/TLB.scala 521:104]
  wire [5:0] _pr_array_T_4 = ~_pr_array_T_3; // @[src/main/scala/rocket/TLB.scala 521:89]
  wire [1:0] _pw_array_T = cacheable ? 2'h3 : 2'h0; // @[src/main/scala/rocket/TLB.scala 523:26]
  wire [5:0] _px_array_T_2 = {_pr_array_T,entries_barrier_3_io_y_px,entries_barrier_2_io_y_px,entries_barrier_1_io_y_px,
    entries_barrier_io_y_px}; // @[src/main/scala/rocket/TLB.scala 525:21]
  wire [5:0] px_array = _px_array_T_2 & _pr_array_T_4; // @[src/main/scala/rocket/TLB.scala 525:87]
  wire [5:0] c_array = {_pw_array_T,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,
    entries_barrier_io_y_c}; // @[src/main/scala/rocket/TLB.scala 529:20]
  wire [39:0] bad_va_maskedVAddr = io_req_bits_vaddr & 40'hc000000000; // @[src/main/scala/rocket/TLB.scala 551:43]
  wire  _bad_va_T_6 = ~(bad_va_maskedVAddr == 40'h0 | bad_va_maskedVAddr == 40'hc000000000); // @[src/main/scala/rocket/TLB.scala 552:37]
  wire  bad_va = vm_enabled & stage1_en & _bad_va_T_6; // @[src/main/scala/rocket/TLB.scala 560:34]
  wire [5:0] _pf_ld_array_T_2 = ~ptw_ae_array; // @[src/main/scala/rocket/TLB.scala 589:73]
  wire [5:0] _pf_ld_array_T_5 = ~ptw_gf_array; // @[src/main/scala/rocket/TLB.scala 589:106]
  wire [5:0] _pf_inst_array_T = ~x_array; // @[src/main/scala/rocket/TLB.scala 591:25]
  wire [5:0] _pf_inst_array_T_2 = _pf_inst_array_T & _pf_ld_array_T_2; // @[src/main/scala/rocket/TLB.scala 591:34]
  wire [5:0] _pf_inst_array_T_3 = _pf_inst_array_T_2 | ptw_pf_array; // @[src/main/scala/rocket/TLB.scala 591:51]
  wire [5:0] pf_inst_array = _pf_inst_array_T_3 & _pf_ld_array_T_5; // @[src/main/scala/rocket/TLB.scala 591:67]
  wire  tlb_hit_if_not_gpa_miss = |real_hits; // @[src/main/scala/rocket/TLB.scala 602:43]
  wire  tlb_miss = vm_enabled & ~bad_va & ~tlb_hit_if_not_gpa_miss; // @[src/main/scala/rocket/TLB.scala 605:64]
  reg  state_vec_0; // @[src/main/scala/util/Replacement.scala 374:17]
  reg  state_reg_1; // @[src/main/scala/util/Replacement.scala 168:72]
  wire  _T_9 = io_req_valid & vm_enabled; // @[src/main/scala/rocket/TLB.scala 609:22]
  wire  line_901_clock;
  wire  line_901_reset;
  wire  line_901_valid;
  reg  line_901_valid_reg;
  wire  _T_10 = sector_hits_0 | sector_hits_1; // @[src/main/scala/util/package.scala 73:59]
  wire  line_902_clock;
  wire  line_902_reset;
  wire  line_902_valid;
  reg  line_902_valid_reg;
  wire [1:0] _T_11 = {sector_hits_1,sector_hits_0}; // @[src/main/scala/chisel3/util/OneHot.scala 21:45]
  wire  state_vec_0_touch_way_sized = _T_11[1]; // @[src/main/scala/chisel3/util/CircuitMath.scala 28:8]
  wire  _state_vec_0_T_1 = ~state_vec_0_touch_way_sized; // @[src/main/scala/util/Replacement.scala 218:7]
  wire  _T_13 = superpage_hits_0 | superpage_hits_1; // @[src/main/scala/util/package.scala 73:59]
  wire  line_903_clock;
  wire  line_903_reset;
  wire  line_903_valid;
  reg  line_903_valid_reg;
  wire [1:0] _T_14 = {superpage_hits_1,superpage_hits_0}; // @[src/main/scala/chisel3/util/OneHot.scala 21:45]
  wire  state_reg_touch_way_sized = _T_14[1]; // @[src/main/scala/chisel3/util/CircuitMath.scala 28:8]
  wire  _state_reg_T_1 = ~state_reg_touch_way_sized; // @[src/main/scala/util/Replacement.scala 218:7]
  wire  multipleHits_leftOne = real_hits[0]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_rightOne = real_hits[1]; // @[src/main/scala/util/Misc.scala 182:39]
  wire  multipleHits_leftOne_1 = multipleHits_leftOne | multipleHits_rightOne; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_leftTwo = multipleHits_leftOne & multipleHits_rightOne; // @[src/main/scala/util/Misc.scala 183:61]
  wire  multipleHits_leftOne_2 = real_hits[2]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_leftOne_3 = real_hits[3]; // @[src/main/scala/util/Misc.scala 181:37]
  wire  multipleHits_rightOne_1 = real_hits[4]; // @[src/main/scala/util/Misc.scala 182:39]
  wire  multipleHits_rightOne_2 = multipleHits_leftOne_3 | multipleHits_rightOne_1; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_rightTwo = multipleHits_leftOne_3 & multipleHits_rightOne_1; // @[src/main/scala/util/Misc.scala 183:61]
  wire  multipleHits_rightOne_3 = multipleHits_leftOne_2 | multipleHits_rightOne_2; // @[src/main/scala/util/Misc.scala 183:16]
  wire  multipleHits_rightTwo_1 = multipleHits_rightTwo | multipleHits_leftOne_2 & multipleHits_rightOne_2; // @[src/main/scala/util/Misc.scala 183:49]
  wire  multipleHits = multipleHits_leftTwo | multipleHits_rightTwo_1 | multipleHits_leftOne_1 & multipleHits_rightOne_3
    ; // @[src/main/scala/util/Misc.scala 183:49]
  wire [5:0] _io_resp_pf_inst_T = pf_inst_array & hits; // @[src/main/scala/rocket/TLB.scala 627:47]
  wire [5:0] _io_resp_ae_inst_T = ~px_array; // @[src/main/scala/rocket/TLB.scala 635:23]
  wire [5:0] _io_resp_ae_inst_T_1 = _io_resp_ae_inst_T & hits; // @[src/main/scala/rocket/TLB.scala 635:33]
  wire [5:0] _io_resp_cacheable_T = c_array & hits; // @[src/main/scala/rocket/TLB.scala 640:33]
  wire  _T_16 = io_ptw_req_ready & io_ptw_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_17 = _T_16 & io_ptw_req_bits_valid; // @[src/main/scala/rocket/TLB.scala 660:26]
  wire  line_904_clock;
  wire  line_904_reset;
  wire  line_904_valid;
  reg  line_904_valid_reg;
  wire  _T_18 = io_req_ready & io_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_19 = _T_18 & tlb_miss; // @[src/main/scala/rocket/TLB.scala 669:23]
  wire  line_905_clock;
  wire  line_905_reset;
  wire  line_905_valid;
  reg  line_905_valid_reg;
  wire [1:0] r_superpage_repl_addr_valids = {superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[src/main/scala/util/package.scala 37:27]
  wire [1:0] _r_superpage_repl_addr_T_2 = ~r_superpage_repl_addr_valids; // @[src/main/scala/rocket/TLB.scala 747:43]
  wire [1:0] r_sectored_repl_addr_valids = {_sector_hits_T_10,_sector_hits_T_2}; // @[src/main/scala/util/package.scala 37:27]
  wire [1:0] _r_sectored_repl_addr_T_2 = ~r_sectored_repl_addr_valids; // @[src/main/scala/rocket/TLB.scala 747:43]
  wire [1:0] _GEN_341 = _T_18 & tlb_miss ? 2'h1 : state; // @[src/main/scala/rocket/TLB.scala 669:36 670:13 341:22]
  wire  line_906_clock;
  wire  line_906_reset;
  wire  line_906_valid;
  reg  line_906_valid_reg;
  wire  line_907_clock;
  wire  line_907_reset;
  wire  line_907_valid;
  reg  line_907_valid_reg;
  wire [1:0] _GEN_352 = io_sfence_valid ? 2'h0 : _GEN_341; // @[src/main/scala/rocket/TLB.scala 691:{21,29}]
  wire  line_908_clock;
  wire  line_908_reset;
  wire  line_908_valid;
  reg  line_908_valid_reg;
  wire [1:0] _state_T = io_sfence_valid ? 2'h3 : 2'h2; // @[src/main/scala/rocket/TLB.scala 694:45]
  wire [1:0] _GEN_353 = io_ptw_req_ready ? _state_T : _GEN_352; // @[src/main/scala/rocket/TLB.scala 694:{31,39}]
  wire  line_909_clock;
  wire  line_909_reset;
  wire  line_909_valid;
  reg  line_909_valid_reg;
  wire [1:0] _GEN_354 = io_kill ? 2'h0 : _GEN_353; // @[src/main/scala/rocket/TLB.scala 696:{22,30}]
  wire  _T_22 = state == 2'h2 & io_sfence_valid; // @[src/main/scala/rocket/TLB.scala 699:28]
  wire  line_910_clock;
  wire  line_910_reset;
  wire  line_910_valid;
  reg  line_910_valid_reg;
  wire  line_911_clock;
  wire  line_911_reset;
  wire  line_911_valid;
  reg  line_911_valid_reg;
  wire  line_912_clock;
  wire  line_912_reset;
  wire  line_912_valid;
  reg  line_912_valid_reg;
  wire  _T_28 = ~reset; // @[src/main/scala/rocket/TLB.scala 709:13]
  wire  line_913_clock;
  wire  line_913_reset;
  wire  line_913_valid;
  reg  line_913_valid_reg;
  wire  _T_29 = ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn); // @[src/main/scala/rocket/TLB.scala 709:13]
  wire  line_914_clock;
  wire  line_914_reset;
  wire  line_914_valid;
  reg  line_914_valid_reg;
  wire  line_915_clock;
  wire  line_915_reset;
  wire  line_915_valid;
  reg  line_915_valid_reg;
  wire  line_916_clock;
  wire  line_916_reset;
  wire  line_916_valid;
  reg  line_916_valid_reg;
  wire  line_917_clock;
  wire  line_917_reset;
  wire  line_917_valid;
  reg  line_917_valid_reg;
  wire  _GEN_358 = _GEN_0 ? 1'h0 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_918_clock;
  wire  line_918_reset;
  wire  line_918_valid;
  reg  line_918_valid_reg;
  wire  _GEN_359 = _GEN_1 ? 1'h0 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_919_clock;
  wire  line_919_reset;
  wire  line_919_valid;
  reg  line_919_valid_reg;
  wire  _GEN_360 = _GEN_2 ? 1'h0 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_920_clock;
  wire  line_920_reset;
  wire  line_920_valid;
  reg  line_920_valid_reg;
  wire  _GEN_361 = _GEN_3 ? 1'h0 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  _GEN_362 = _sector_hits_T_5 ? _GEN_358 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_363 = _sector_hits_T_5 ? _GEN_359 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_364 = _sector_hits_T_5 ? _GEN_360 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_365 = _sector_hits_T_5 ? _GEN_361 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _T_147 = _sector_hits_T_3[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_921_clock;
  wire  line_921_reset;
  wire  line_921_valid;
  reg  line_921_valid_reg;
  wire  line_922_clock;
  wire  line_922_reset;
  wire  line_922_valid;
  reg  line_922_valid_reg;
  wire  _GEN_366 = sectored_entries_0_0_data_0[0] ? 1'h0 : _GEN_362; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_923_clock;
  wire  line_923_reset;
  wire  line_923_valid;
  reg  line_923_valid_reg;
  wire  _GEN_367 = sectored_entries_0_0_data_1[0] ? 1'h0 : _GEN_363; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_924_clock;
  wire  line_924_reset;
  wire  line_924_valid;
  reg  line_924_valid_reg;
  wire  _GEN_368 = sectored_entries_0_0_data_2[0] ? 1'h0 : _GEN_364; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_925_clock;
  wire  line_925_reset;
  wire  line_925_valid;
  reg  line_925_valid_reg;
  wire  _GEN_369 = sectored_entries_0_0_data_3[0] ? 1'h0 : _GEN_365; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_926_clock;
  wire  line_926_reset;
  wire  line_926_valid;
  reg  line_926_valid_reg;
  wire  line_927_clock;
  wire  line_927_reset;
  wire  line_927_valid;
  reg  line_927_valid_reg;
  wire  _T_343 = ~sectored_entries_0_0_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_928_clock;
  wire  line_928_reset;
  wire  line_928_valid;
  reg  line_928_valid_reg;
  wire  _GEN_374 = ~sectored_entries_0_0_data_0[20] ? 1'h0 : _GEN_302; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_346 = ~sectored_entries_0_0_data_1[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_929_clock;
  wire  line_929_reset;
  wire  line_929_valid;
  reg  line_929_valid_reg;
  wire  _GEN_375 = ~sectored_entries_0_0_data_1[20] ? 1'h0 : _GEN_303; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_349 = ~sectored_entries_0_0_data_2[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_930_clock;
  wire  line_930_reset;
  wire  line_930_valid;
  reg  line_930_valid_reg;
  wire  _GEN_376 = ~sectored_entries_0_0_data_2[20] ? 1'h0 : _GEN_304; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_352 = ~sectored_entries_0_0_data_3[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_931_clock;
  wire  line_931_reset;
  wire  line_931_valid;
  reg  line_931_valid_reg;
  wire  _GEN_377 = ~sectored_entries_0_0_data_3[20] ? 1'h0 : _GEN_305; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_932_clock;
  wire  line_932_reset;
  wire  line_932_valid;
  reg  line_932_valid_reg;
  wire  _GEN_382 = io_sfence_bits_rs2 & _GEN_374; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_383 = io_sfence_bits_rs2 & _GEN_375; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_384 = io_sfence_bits_rs2 & _GEN_376; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_385 = io_sfence_bits_rs2 & _GEN_377; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_933_clock;
  wire  line_933_reset;
  wire  line_933_valid;
  reg  line_933_valid_reg;
  wire  line_934_clock;
  wire  line_934_reset;
  wire  line_934_valid;
  reg  line_934_valid_reg;
  wire  line_935_clock;
  wire  line_935_reset;
  wire  line_935_valid;
  reg  line_935_valid_reg;
  wire  _GEN_390 = _GEN_0 ? 1'h0 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_936_clock;
  wire  line_936_reset;
  wire  line_936_valid;
  reg  line_936_valid_reg;
  wire  _GEN_391 = _GEN_1 ? 1'h0 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_937_clock;
  wire  line_937_reset;
  wire  line_937_valid;
  reg  line_937_valid_reg;
  wire  _GEN_392 = _GEN_2 ? 1'h0 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  line_938_clock;
  wire  line_938_reset;
  wire  line_938_valid;
  reg  line_938_valid_reg;
  wire  _GEN_393 = _GEN_3 ? 1'h0 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 221:{62,66}]
  wire  _GEN_394 = _sector_hits_T_13 ? _GEN_390 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_395 = _sector_hits_T_13 ? _GEN_391 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_396 = _sector_hits_T_13 ? _GEN_392 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _GEN_397 = _sector_hits_T_13 ? _GEN_393 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 219:43]
  wire  _T_568 = _sector_hits_T_11[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_939_clock;
  wire  line_939_reset;
  wire  line_939_valid;
  reg  line_939_valid_reg;
  wire  line_940_clock;
  wire  line_940_reset;
  wire  line_940_valid;
  reg  line_940_valid_reg;
  wire  _GEN_398 = sectored_entries_0_1_data_0[0] ? 1'h0 : _GEN_394; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_941_clock;
  wire  line_941_reset;
  wire  line_941_valid;
  reg  line_941_valid_reg;
  wire  _GEN_399 = sectored_entries_0_1_data_1[0] ? 1'h0 : _GEN_395; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_942_clock;
  wire  line_942_reset;
  wire  line_942_valid;
  reg  line_942_valid_reg;
  wire  _GEN_400 = sectored_entries_0_1_data_2[0] ? 1'h0 : _GEN_396; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_943_clock;
  wire  line_943_reset;
  wire  line_943_valid;
  reg  line_943_valid_reg;
  wire  _GEN_401 = sectored_entries_0_1_data_3[0] ? 1'h0 : _GEN_397; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_944_clock;
  wire  line_944_reset;
  wire  line_944_valid;
  reg  line_944_valid_reg;
  wire  line_945_clock;
  wire  line_945_reset;
  wire  line_945_valid;
  reg  line_945_valid_reg;
  wire  _T_764 = ~sectored_entries_0_1_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_946_clock;
  wire  line_946_reset;
  wire  line_946_valid;
  reg  line_946_valid_reg;
  wire  _GEN_406 = ~sectored_entries_0_1_data_0[20] ? 1'h0 : _GEN_313; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_767 = ~sectored_entries_0_1_data_1[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_947_clock;
  wire  line_947_reset;
  wire  line_947_valid;
  reg  line_947_valid_reg;
  wire  _GEN_407 = ~sectored_entries_0_1_data_1[20] ? 1'h0 : _GEN_314; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_770 = ~sectored_entries_0_1_data_2[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_948_clock;
  wire  line_948_reset;
  wire  line_948_valid;
  reg  line_948_valid_reg;
  wire  _GEN_408 = ~sectored_entries_0_1_data_2[20] ? 1'h0 : _GEN_315; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  _T_773 = ~sectored_entries_0_1_data_3[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_949_clock;
  wire  line_949_reset;
  wire  line_949_valid;
  reg  line_949_valid_reg;
  wire  _GEN_409 = ~sectored_entries_0_1_data_3[20] ? 1'h0 : _GEN_316; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_950_clock;
  wire  line_950_reset;
  wire  line_950_valid;
  reg  line_950_valid_reg;
  wire  _GEN_414 = io_sfence_bits_rs2 & _GEN_406; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_415 = io_sfence_bits_rs2 & _GEN_407; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_416 = io_sfence_bits_rs2 & _GEN_408; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _GEN_417 = io_sfence_bits_rs2 & _GEN_409; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_951_clock;
  wire  line_951_reset;
  wire  line_951_valid;
  reg  line_951_valid_reg;
  wire  line_952_clock;
  wire  line_952_reset;
  wire  line_952_valid;
  reg  line_952_valid_reg;
  wire  _GEN_422 = superpage_hits_0 ? 1'h0 : _GEN_295; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_891 = _superpage_hits_T[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_953_clock;
  wire  line_953_reset;
  wire  line_953_valid;
  reg  line_953_valid_reg;
  wire  line_954_clock;
  wire  line_954_reset;
  wire  line_954_valid;
  reg  line_954_valid_reg;
  wire  _GEN_423 = superpage_entries_0_data_0[0] ? 1'h0 : _GEN_422; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_955_clock;
  wire  line_955_reset;
  wire  line_955_valid;
  reg  line_955_valid_reg;
  wire  line_956_clock;
  wire  line_956_reset;
  wire  line_956_valid;
  reg  line_956_valid_reg;
  wire  _T_943 = ~superpage_entries_0_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_957_clock;
  wire  line_957_reset;
  wire  line_957_valid;
  reg  line_957_valid_reg;
  wire  _GEN_425 = ~superpage_entries_0_data_0[20] ? 1'h0 : _GEN_295; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_958_clock;
  wire  line_958_reset;
  wire  line_958_valid;
  reg  line_958_valid_reg;
  wire  _GEN_427 = io_sfence_bits_rs2 & _GEN_425; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_959_clock;
  wire  line_959_reset;
  wire  line_959_valid;
  reg  line_959_valid_reg;
  wire  line_960_clock;
  wire  line_960_reset;
  wire  line_960_valid;
  reg  line_960_valid_reg;
  wire  _GEN_429 = superpage_hits_1 ? 1'h0 : _GEN_300; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_989 = _superpage_hits_T_14[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_961_clock;
  wire  line_961_reset;
  wire  line_961_valid;
  reg  line_961_valid_reg;
  wire  line_962_clock;
  wire  line_962_reset;
  wire  line_962_valid;
  reg  line_962_valid_reg;
  wire  _GEN_430 = superpage_entries_1_data_0[0] ? 1'h0 : _GEN_429; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_963_clock;
  wire  line_963_reset;
  wire  line_963_valid;
  reg  line_963_valid_reg;
  wire  line_964_clock;
  wire  line_964_reset;
  wire  line_964_valid;
  reg  line_964_valid_reg;
  wire  _T_1041 = ~superpage_entries_1_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_965_clock;
  wire  line_965_reset;
  wire  line_965_valid;
  reg  line_965_valid_reg;
  wire  _GEN_432 = ~superpage_entries_1_data_0[20] ? 1'h0 : _GEN_300; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_966_clock;
  wire  line_966_reset;
  wire  line_966_valid;
  reg  line_966_valid_reg;
  wire  _GEN_434 = io_sfence_bits_rs2 & _GEN_432; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  line_967_clock;
  wire  line_967_reset;
  wire  line_967_valid;
  reg  line_967_valid_reg;
  wire  line_968_clock;
  wire  line_968_reset;
  wire  line_968_valid;
  reg  line_968_valid_reg;
  wire  _GEN_436 = _hitsVec_T_56 ? 1'h0 : _GEN_290; // @[src/main/scala/rocket/TLB.scala 217:32 210:46]
  wire  _T_1087 = _hitsVec_T_42[26:18] == 9'h0; // @[src/main/scala/rocket/TLB.scala 226:63]
  wire  line_969_clock;
  wire  line_969_reset;
  wire  line_969_valid;
  reg  line_969_valid_reg;
  wire  line_970_clock;
  wire  line_970_reset;
  wire  line_970_valid;
  reg  line_970_valid_reg;
  wire  _GEN_437 = special_entry_data_0[0] ? 1'h0 : _GEN_436; // @[src/main/scala/rocket/TLB.scala 228:{60,64}]
  wire  line_971_clock;
  wire  line_971_reset;
  wire  line_971_valid;
  reg  line_971_valid_reg;
  wire  line_972_clock;
  wire  line_972_reset;
  wire  line_972_valid;
  reg  line_972_valid_reg;
  wire  _T_1139 = ~special_entry_data_0[20]; // @[src/main/scala/rocket/TLB.scala 233:34]
  wire  line_973_clock;
  wire  line_973_reset;
  wire  line_973_valid;
  reg  line_973_valid_reg;
  wire  _GEN_439 = ~special_entry_data_0[20] ? 1'h0 : _GEN_290; // @[src/main/scala/rocket/TLB.scala 233:{40,44}]
  wire  line_974_clock;
  wire  line_974_reset;
  wire  line_974_valid;
  reg  line_974_valid_reg;
  wire  _GEN_441 = io_sfence_bits_rs2 & _GEN_439; // @[src/main/scala/rocket/TLB.scala 714:47]
  wire  _T_1433 = multipleHits | reset; // @[src/main/scala/rocket/TLB.scala 722:24]
  wire  line_975_clock;
  wire  line_975_reset;
  wire  line_975_valid;
  reg  line_975_valid_reg;
  OptimizationBarrier_12 mpu_ppn_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(mpu_ppn_barrier_clock),
    .reset(mpu_ppn_barrier_reset),
    .io_x_ppn(mpu_ppn_barrier_io_x_ppn),
    .io_y_ppn(mpu_ppn_barrier_io_y_ppn)
  );
  PMPChecker_2 pmp ( // @[src/main/scala/rocket/TLB.scala 405:19]
    .clock(pmp_clock),
    .reset(pmp_reset)
  );
  OptimizationBarrier_13 entries_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_clock),
    .reset(entries_barrier_reset),
    .io_x_ppn(entries_barrier_io_x_ppn),
    .io_x_u(entries_barrier_io_x_u),
    .io_x_ae_ptw(entries_barrier_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_io_x_ae_final),
    .io_x_pf(entries_barrier_io_x_pf),
    .io_x_gf(entries_barrier_io_x_gf),
    .io_x_sx(entries_barrier_io_x_sx),
    .io_x_px(entries_barrier_io_x_px),
    .io_x_c(entries_barrier_io_x_c),
    .io_y_ppn(entries_barrier_io_y_ppn),
    .io_y_u(entries_barrier_io_y_u),
    .io_y_ae_ptw(entries_barrier_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_io_y_ae_final),
    .io_y_pf(entries_barrier_io_y_pf),
    .io_y_gf(entries_barrier_io_y_gf),
    .io_y_sx(entries_barrier_io_y_sx),
    .io_y_px(entries_barrier_io_y_px),
    .io_y_c(entries_barrier_io_y_c)
  );
  OptimizationBarrier_14 entries_barrier_1 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_1_clock),
    .reset(entries_barrier_1_reset),
    .io_x_ppn(entries_barrier_1_io_x_ppn),
    .io_x_u(entries_barrier_1_io_x_u),
    .io_x_ae_ptw(entries_barrier_1_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_1_io_x_ae_final),
    .io_x_pf(entries_barrier_1_io_x_pf),
    .io_x_gf(entries_barrier_1_io_x_gf),
    .io_x_sx(entries_barrier_1_io_x_sx),
    .io_x_px(entries_barrier_1_io_x_px),
    .io_x_c(entries_barrier_1_io_x_c),
    .io_y_ppn(entries_barrier_1_io_y_ppn),
    .io_y_u(entries_barrier_1_io_y_u),
    .io_y_ae_ptw(entries_barrier_1_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_1_io_y_ae_final),
    .io_y_pf(entries_barrier_1_io_y_pf),
    .io_y_gf(entries_barrier_1_io_y_gf),
    .io_y_sx(entries_barrier_1_io_y_sx),
    .io_y_px(entries_barrier_1_io_y_px),
    .io_y_c(entries_barrier_1_io_y_c)
  );
  OptimizationBarrier_15 entries_barrier_2 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_2_clock),
    .reset(entries_barrier_2_reset),
    .io_x_ppn(entries_barrier_2_io_x_ppn),
    .io_x_u(entries_barrier_2_io_x_u),
    .io_x_ae_ptw(entries_barrier_2_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_2_io_x_ae_final),
    .io_x_pf(entries_barrier_2_io_x_pf),
    .io_x_gf(entries_barrier_2_io_x_gf),
    .io_x_sx(entries_barrier_2_io_x_sx),
    .io_x_px(entries_barrier_2_io_x_px),
    .io_x_c(entries_barrier_2_io_x_c),
    .io_y_ppn(entries_barrier_2_io_y_ppn),
    .io_y_u(entries_barrier_2_io_y_u),
    .io_y_ae_ptw(entries_barrier_2_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_2_io_y_ae_final),
    .io_y_pf(entries_barrier_2_io_y_pf),
    .io_y_gf(entries_barrier_2_io_y_gf),
    .io_y_sx(entries_barrier_2_io_y_sx),
    .io_y_px(entries_barrier_2_io_y_px),
    .io_y_c(entries_barrier_2_io_y_c)
  );
  OptimizationBarrier_16 entries_barrier_3 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_3_clock),
    .reset(entries_barrier_3_reset),
    .io_x_ppn(entries_barrier_3_io_x_ppn),
    .io_x_u(entries_barrier_3_io_x_u),
    .io_x_ae_ptw(entries_barrier_3_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_3_io_x_ae_final),
    .io_x_pf(entries_barrier_3_io_x_pf),
    .io_x_gf(entries_barrier_3_io_x_gf),
    .io_x_sx(entries_barrier_3_io_x_sx),
    .io_x_px(entries_barrier_3_io_x_px),
    .io_x_c(entries_barrier_3_io_x_c),
    .io_y_ppn(entries_barrier_3_io_y_ppn),
    .io_y_u(entries_barrier_3_io_y_u),
    .io_y_ae_ptw(entries_barrier_3_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_3_io_y_ae_final),
    .io_y_pf(entries_barrier_3_io_y_pf),
    .io_y_gf(entries_barrier_3_io_y_gf),
    .io_y_sx(entries_barrier_3_io_y_sx),
    .io_y_px(entries_barrier_3_io_y_px),
    .io_y_c(entries_barrier_3_io_y_c)
  );
  OptimizationBarrier_17 entries_barrier_4 ( // @[src/main/scala/util/package.scala 259:25]
    .clock(entries_barrier_4_clock),
    .reset(entries_barrier_4_reset),
    .io_x_ppn(entries_barrier_4_io_x_ppn),
    .io_x_u(entries_barrier_4_io_x_u),
    .io_x_ae_ptw(entries_barrier_4_io_x_ae_ptw),
    .io_x_ae_final(entries_barrier_4_io_x_ae_final),
    .io_x_pf(entries_barrier_4_io_x_pf),
    .io_x_gf(entries_barrier_4_io_x_gf),
    .io_x_sx(entries_barrier_4_io_x_sx),
    .io_y_ppn(entries_barrier_4_io_y_ppn),
    .io_y_u(entries_barrier_4_io_y_u),
    .io_y_ae_ptw(entries_barrier_4_io_y_ae_ptw),
    .io_y_ae_final(entries_barrier_4_io_y_ae_final),
    .io_y_pf(entries_barrier_4_io_y_pf),
    .io_y_gf(entries_barrier_4_io_y_gf),
    .io_y_sx(entries_barrier_4_io_y_sx)
  );
  GEN_w1_line #(.COVER_INDEX(854)) line_854 (
    .clock(line_854_clock),
    .reset(line_854_reset),
    .valid(line_854_valid)
  );
  GEN_w1_line #(.COVER_INDEX(855)) line_855 (
    .clock(line_855_clock),
    .reset(line_855_reset),
    .valid(line_855_valid)
  );
  GEN_w1_line #(.COVER_INDEX(856)) line_856 (
    .clock(line_856_clock),
    .reset(line_856_reset),
    .valid(line_856_valid)
  );
  GEN_w1_line #(.COVER_INDEX(857)) line_857 (
    .clock(line_857_clock),
    .reset(line_857_reset),
    .valid(line_857_valid)
  );
  GEN_w1_line #(.COVER_INDEX(858)) line_858 (
    .clock(line_858_clock),
    .reset(line_858_reset),
    .valid(line_858_valid)
  );
  GEN_w1_line #(.COVER_INDEX(859)) line_859 (
    .clock(line_859_clock),
    .reset(line_859_reset),
    .valid(line_859_valid)
  );
  GEN_w1_line #(.COVER_INDEX(860)) line_860 (
    .clock(line_860_clock),
    .reset(line_860_reset),
    .valid(line_860_valid)
  );
  GEN_w1_line #(.COVER_INDEX(861)) line_861 (
    .clock(line_861_clock),
    .reset(line_861_reset),
    .valid(line_861_valid)
  );
  GEN_w1_line #(.COVER_INDEX(862)) line_862 (
    .clock(line_862_clock),
    .reset(line_862_reset),
    .valid(line_862_valid)
  );
  GEN_w1_line #(.COVER_INDEX(863)) line_863 (
    .clock(line_863_clock),
    .reset(line_863_reset),
    .valid(line_863_valid)
  );
  GEN_w1_line #(.COVER_INDEX(864)) line_864 (
    .clock(line_864_clock),
    .reset(line_864_reset),
    .valid(line_864_valid)
  );
  GEN_w1_line #(.COVER_INDEX(865)) line_865 (
    .clock(line_865_clock),
    .reset(line_865_reset),
    .valid(line_865_valid)
  );
  GEN_w1_line #(.COVER_INDEX(866)) line_866 (
    .clock(line_866_clock),
    .reset(line_866_reset),
    .valid(line_866_valid)
  );
  GEN_w1_line #(.COVER_INDEX(867)) line_867 (
    .clock(line_867_clock),
    .reset(line_867_reset),
    .valid(line_867_valid)
  );
  GEN_w1_line #(.COVER_INDEX(868)) line_868 (
    .clock(line_868_clock),
    .reset(line_868_reset),
    .valid(line_868_valid)
  );
  GEN_w1_line #(.COVER_INDEX(869)) line_869 (
    .clock(line_869_clock),
    .reset(line_869_reset),
    .valid(line_869_valid)
  );
  GEN_w1_line #(.COVER_INDEX(870)) line_870 (
    .clock(line_870_clock),
    .reset(line_870_reset),
    .valid(line_870_valid)
  );
  GEN_w1_line #(.COVER_INDEX(871)) line_871 (
    .clock(line_871_clock),
    .reset(line_871_reset),
    .valid(line_871_valid)
  );
  GEN_w1_line #(.COVER_INDEX(872)) line_872 (
    .clock(line_872_clock),
    .reset(line_872_reset),
    .valid(line_872_valid)
  );
  GEN_w1_line #(.COVER_INDEX(873)) line_873 (
    .clock(line_873_clock),
    .reset(line_873_reset),
    .valid(line_873_valid)
  );
  GEN_w1_line #(.COVER_INDEX(874)) line_874 (
    .clock(line_874_clock),
    .reset(line_874_reset),
    .valid(line_874_valid)
  );
  GEN_w1_line #(.COVER_INDEX(875)) line_875 (
    .clock(line_875_clock),
    .reset(line_875_reset),
    .valid(line_875_valid)
  );
  GEN_w1_line #(.COVER_INDEX(876)) line_876 (
    .clock(line_876_clock),
    .reset(line_876_reset),
    .valid(line_876_valid)
  );
  GEN_w1_line #(.COVER_INDEX(877)) line_877 (
    .clock(line_877_clock),
    .reset(line_877_reset),
    .valid(line_877_valid)
  );
  GEN_w1_line #(.COVER_INDEX(878)) line_878 (
    .clock(line_878_clock),
    .reset(line_878_reset),
    .valid(line_878_valid)
  );
  GEN_w1_line #(.COVER_INDEX(879)) line_879 (
    .clock(line_879_clock),
    .reset(line_879_reset),
    .valid(line_879_valid)
  );
  GEN_w1_line #(.COVER_INDEX(880)) line_880 (
    .clock(line_880_clock),
    .reset(line_880_reset),
    .valid(line_880_valid)
  );
  GEN_w1_line #(.COVER_INDEX(881)) line_881 (
    .clock(line_881_clock),
    .reset(line_881_reset),
    .valid(line_881_valid)
  );
  GEN_w1_line #(.COVER_INDEX(882)) line_882 (
    .clock(line_882_clock),
    .reset(line_882_reset),
    .valid(line_882_valid)
  );
  GEN_w1_line #(.COVER_INDEX(883)) line_883 (
    .clock(line_883_clock),
    .reset(line_883_reset),
    .valid(line_883_valid)
  );
  GEN_w1_line #(.COVER_INDEX(884)) line_884 (
    .clock(line_884_clock),
    .reset(line_884_reset),
    .valid(line_884_valid)
  );
  GEN_w1_line #(.COVER_INDEX(885)) line_885 (
    .clock(line_885_clock),
    .reset(line_885_reset),
    .valid(line_885_valid)
  );
  GEN_w1_line #(.COVER_INDEX(886)) line_886 (
    .clock(line_886_clock),
    .reset(line_886_reset),
    .valid(line_886_valid)
  );
  GEN_w1_line #(.COVER_INDEX(887)) line_887 (
    .clock(line_887_clock),
    .reset(line_887_reset),
    .valid(line_887_valid)
  );
  GEN_w1_line #(.COVER_INDEX(888)) line_888 (
    .clock(line_888_clock),
    .reset(line_888_reset),
    .valid(line_888_valid)
  );
  GEN_w1_line #(.COVER_INDEX(889)) line_889 (
    .clock(line_889_clock),
    .reset(line_889_reset),
    .valid(line_889_valid)
  );
  GEN_w1_line #(.COVER_INDEX(890)) line_890 (
    .clock(line_890_clock),
    .reset(line_890_reset),
    .valid(line_890_valid)
  );
  GEN_w1_line #(.COVER_INDEX(891)) line_891 (
    .clock(line_891_clock),
    .reset(line_891_reset),
    .valid(line_891_valid)
  );
  GEN_w1_line #(.COVER_INDEX(892)) line_892 (
    .clock(line_892_clock),
    .reset(line_892_reset),
    .valid(line_892_valid)
  );
  GEN_w1_line #(.COVER_INDEX(893)) line_893 (
    .clock(line_893_clock),
    .reset(line_893_reset),
    .valid(line_893_valid)
  );
  GEN_w1_line #(.COVER_INDEX(894)) line_894 (
    .clock(line_894_clock),
    .reset(line_894_reset),
    .valid(line_894_valid)
  );
  GEN_w1_line #(.COVER_INDEX(895)) line_895 (
    .clock(line_895_clock),
    .reset(line_895_reset),
    .valid(line_895_valid)
  );
  GEN_w1_line #(.COVER_INDEX(896)) line_896 (
    .clock(line_896_clock),
    .reset(line_896_reset),
    .valid(line_896_valid)
  );
  GEN_w1_line #(.COVER_INDEX(897)) line_897 (
    .clock(line_897_clock),
    .reset(line_897_reset),
    .valid(line_897_valid)
  );
  GEN_w1_line #(.COVER_INDEX(898)) line_898 (
    .clock(line_898_clock),
    .reset(line_898_reset),
    .valid(line_898_valid)
  );
  GEN_w1_line #(.COVER_INDEX(899)) line_899 (
    .clock(line_899_clock),
    .reset(line_899_reset),
    .valid(line_899_valid)
  );
  GEN_w1_line #(.COVER_INDEX(900)) line_900 (
    .clock(line_900_clock),
    .reset(line_900_reset),
    .valid(line_900_valid)
  );
  GEN_w1_line #(.COVER_INDEX(901)) line_901 (
    .clock(line_901_clock),
    .reset(line_901_reset),
    .valid(line_901_valid)
  );
  GEN_w1_line #(.COVER_INDEX(902)) line_902 (
    .clock(line_902_clock),
    .reset(line_902_reset),
    .valid(line_902_valid)
  );
  GEN_w1_line #(.COVER_INDEX(903)) line_903 (
    .clock(line_903_clock),
    .reset(line_903_reset),
    .valid(line_903_valid)
  );
  GEN_w1_line #(.COVER_INDEX(904)) line_904 (
    .clock(line_904_clock),
    .reset(line_904_reset),
    .valid(line_904_valid)
  );
  GEN_w1_line #(.COVER_INDEX(905)) line_905 (
    .clock(line_905_clock),
    .reset(line_905_reset),
    .valid(line_905_valid)
  );
  GEN_w1_line #(.COVER_INDEX(906)) line_906 (
    .clock(line_906_clock),
    .reset(line_906_reset),
    .valid(line_906_valid)
  );
  GEN_w1_line #(.COVER_INDEX(907)) line_907 (
    .clock(line_907_clock),
    .reset(line_907_reset),
    .valid(line_907_valid)
  );
  GEN_w1_line #(.COVER_INDEX(908)) line_908 (
    .clock(line_908_clock),
    .reset(line_908_reset),
    .valid(line_908_valid)
  );
  GEN_w1_line #(.COVER_INDEX(909)) line_909 (
    .clock(line_909_clock),
    .reset(line_909_reset),
    .valid(line_909_valid)
  );
  GEN_w1_line #(.COVER_INDEX(910)) line_910 (
    .clock(line_910_clock),
    .reset(line_910_reset),
    .valid(line_910_valid)
  );
  GEN_w1_line #(.COVER_INDEX(911)) line_911 (
    .clock(line_911_clock),
    .reset(line_911_reset),
    .valid(line_911_valid)
  );
  GEN_w1_line #(.COVER_INDEX(912)) line_912 (
    .clock(line_912_clock),
    .reset(line_912_reset),
    .valid(line_912_valid)
  );
  GEN_w1_line #(.COVER_INDEX(913)) line_913 (
    .clock(line_913_clock),
    .reset(line_913_reset),
    .valid(line_913_valid)
  );
  GEN_w1_line #(.COVER_INDEX(914)) line_914 (
    .clock(line_914_clock),
    .reset(line_914_reset),
    .valid(line_914_valid)
  );
  GEN_w1_line #(.COVER_INDEX(915)) line_915 (
    .clock(line_915_clock),
    .reset(line_915_reset),
    .valid(line_915_valid)
  );
  GEN_w1_line #(.COVER_INDEX(916)) line_916 (
    .clock(line_916_clock),
    .reset(line_916_reset),
    .valid(line_916_valid)
  );
  GEN_w1_line #(.COVER_INDEX(917)) line_917 (
    .clock(line_917_clock),
    .reset(line_917_reset),
    .valid(line_917_valid)
  );
  GEN_w1_line #(.COVER_INDEX(918)) line_918 (
    .clock(line_918_clock),
    .reset(line_918_reset),
    .valid(line_918_valid)
  );
  GEN_w1_line #(.COVER_INDEX(919)) line_919 (
    .clock(line_919_clock),
    .reset(line_919_reset),
    .valid(line_919_valid)
  );
  GEN_w1_line #(.COVER_INDEX(920)) line_920 (
    .clock(line_920_clock),
    .reset(line_920_reset),
    .valid(line_920_valid)
  );
  GEN_w1_line #(.COVER_INDEX(921)) line_921 (
    .clock(line_921_clock),
    .reset(line_921_reset),
    .valid(line_921_valid)
  );
  GEN_w1_line #(.COVER_INDEX(922)) line_922 (
    .clock(line_922_clock),
    .reset(line_922_reset),
    .valid(line_922_valid)
  );
  GEN_w1_line #(.COVER_INDEX(923)) line_923 (
    .clock(line_923_clock),
    .reset(line_923_reset),
    .valid(line_923_valid)
  );
  GEN_w1_line #(.COVER_INDEX(924)) line_924 (
    .clock(line_924_clock),
    .reset(line_924_reset),
    .valid(line_924_valid)
  );
  GEN_w1_line #(.COVER_INDEX(925)) line_925 (
    .clock(line_925_clock),
    .reset(line_925_reset),
    .valid(line_925_valid)
  );
  GEN_w1_line #(.COVER_INDEX(926)) line_926 (
    .clock(line_926_clock),
    .reset(line_926_reset),
    .valid(line_926_valid)
  );
  GEN_w1_line #(.COVER_INDEX(927)) line_927 (
    .clock(line_927_clock),
    .reset(line_927_reset),
    .valid(line_927_valid)
  );
  GEN_w1_line #(.COVER_INDEX(928)) line_928 (
    .clock(line_928_clock),
    .reset(line_928_reset),
    .valid(line_928_valid)
  );
  GEN_w1_line #(.COVER_INDEX(929)) line_929 (
    .clock(line_929_clock),
    .reset(line_929_reset),
    .valid(line_929_valid)
  );
  GEN_w1_line #(.COVER_INDEX(930)) line_930 (
    .clock(line_930_clock),
    .reset(line_930_reset),
    .valid(line_930_valid)
  );
  GEN_w1_line #(.COVER_INDEX(931)) line_931 (
    .clock(line_931_clock),
    .reset(line_931_reset),
    .valid(line_931_valid)
  );
  GEN_w1_line #(.COVER_INDEX(932)) line_932 (
    .clock(line_932_clock),
    .reset(line_932_reset),
    .valid(line_932_valid)
  );
  GEN_w1_line #(.COVER_INDEX(933)) line_933 (
    .clock(line_933_clock),
    .reset(line_933_reset),
    .valid(line_933_valid)
  );
  GEN_w1_line #(.COVER_INDEX(934)) line_934 (
    .clock(line_934_clock),
    .reset(line_934_reset),
    .valid(line_934_valid)
  );
  GEN_w1_line #(.COVER_INDEX(935)) line_935 (
    .clock(line_935_clock),
    .reset(line_935_reset),
    .valid(line_935_valid)
  );
  GEN_w1_line #(.COVER_INDEX(936)) line_936 (
    .clock(line_936_clock),
    .reset(line_936_reset),
    .valid(line_936_valid)
  );
  GEN_w1_line #(.COVER_INDEX(937)) line_937 (
    .clock(line_937_clock),
    .reset(line_937_reset),
    .valid(line_937_valid)
  );
  GEN_w1_line #(.COVER_INDEX(938)) line_938 (
    .clock(line_938_clock),
    .reset(line_938_reset),
    .valid(line_938_valid)
  );
  GEN_w1_line #(.COVER_INDEX(939)) line_939 (
    .clock(line_939_clock),
    .reset(line_939_reset),
    .valid(line_939_valid)
  );
  GEN_w1_line #(.COVER_INDEX(940)) line_940 (
    .clock(line_940_clock),
    .reset(line_940_reset),
    .valid(line_940_valid)
  );
  GEN_w1_line #(.COVER_INDEX(941)) line_941 (
    .clock(line_941_clock),
    .reset(line_941_reset),
    .valid(line_941_valid)
  );
  GEN_w1_line #(.COVER_INDEX(942)) line_942 (
    .clock(line_942_clock),
    .reset(line_942_reset),
    .valid(line_942_valid)
  );
  GEN_w1_line #(.COVER_INDEX(943)) line_943 (
    .clock(line_943_clock),
    .reset(line_943_reset),
    .valid(line_943_valid)
  );
  GEN_w1_line #(.COVER_INDEX(944)) line_944 (
    .clock(line_944_clock),
    .reset(line_944_reset),
    .valid(line_944_valid)
  );
  GEN_w1_line #(.COVER_INDEX(945)) line_945 (
    .clock(line_945_clock),
    .reset(line_945_reset),
    .valid(line_945_valid)
  );
  GEN_w1_line #(.COVER_INDEX(946)) line_946 (
    .clock(line_946_clock),
    .reset(line_946_reset),
    .valid(line_946_valid)
  );
  GEN_w1_line #(.COVER_INDEX(947)) line_947 (
    .clock(line_947_clock),
    .reset(line_947_reset),
    .valid(line_947_valid)
  );
  GEN_w1_line #(.COVER_INDEX(948)) line_948 (
    .clock(line_948_clock),
    .reset(line_948_reset),
    .valid(line_948_valid)
  );
  GEN_w1_line #(.COVER_INDEX(949)) line_949 (
    .clock(line_949_clock),
    .reset(line_949_reset),
    .valid(line_949_valid)
  );
  GEN_w1_line #(.COVER_INDEX(950)) line_950 (
    .clock(line_950_clock),
    .reset(line_950_reset),
    .valid(line_950_valid)
  );
  GEN_w1_line #(.COVER_INDEX(951)) line_951 (
    .clock(line_951_clock),
    .reset(line_951_reset),
    .valid(line_951_valid)
  );
  GEN_w1_line #(.COVER_INDEX(952)) line_952 (
    .clock(line_952_clock),
    .reset(line_952_reset),
    .valid(line_952_valid)
  );
  GEN_w1_line #(.COVER_INDEX(953)) line_953 (
    .clock(line_953_clock),
    .reset(line_953_reset),
    .valid(line_953_valid)
  );
  GEN_w1_line #(.COVER_INDEX(954)) line_954 (
    .clock(line_954_clock),
    .reset(line_954_reset),
    .valid(line_954_valid)
  );
  GEN_w1_line #(.COVER_INDEX(955)) line_955 (
    .clock(line_955_clock),
    .reset(line_955_reset),
    .valid(line_955_valid)
  );
  GEN_w1_line #(.COVER_INDEX(956)) line_956 (
    .clock(line_956_clock),
    .reset(line_956_reset),
    .valid(line_956_valid)
  );
  GEN_w1_line #(.COVER_INDEX(957)) line_957 (
    .clock(line_957_clock),
    .reset(line_957_reset),
    .valid(line_957_valid)
  );
  GEN_w1_line #(.COVER_INDEX(958)) line_958 (
    .clock(line_958_clock),
    .reset(line_958_reset),
    .valid(line_958_valid)
  );
  GEN_w1_line #(.COVER_INDEX(959)) line_959 (
    .clock(line_959_clock),
    .reset(line_959_reset),
    .valid(line_959_valid)
  );
  GEN_w1_line #(.COVER_INDEX(960)) line_960 (
    .clock(line_960_clock),
    .reset(line_960_reset),
    .valid(line_960_valid)
  );
  GEN_w1_line #(.COVER_INDEX(961)) line_961 (
    .clock(line_961_clock),
    .reset(line_961_reset),
    .valid(line_961_valid)
  );
  GEN_w1_line #(.COVER_INDEX(962)) line_962 (
    .clock(line_962_clock),
    .reset(line_962_reset),
    .valid(line_962_valid)
  );
  GEN_w1_line #(.COVER_INDEX(963)) line_963 (
    .clock(line_963_clock),
    .reset(line_963_reset),
    .valid(line_963_valid)
  );
  GEN_w1_line #(.COVER_INDEX(964)) line_964 (
    .clock(line_964_clock),
    .reset(line_964_reset),
    .valid(line_964_valid)
  );
  GEN_w1_line #(.COVER_INDEX(965)) line_965 (
    .clock(line_965_clock),
    .reset(line_965_reset),
    .valid(line_965_valid)
  );
  GEN_w1_line #(.COVER_INDEX(966)) line_966 (
    .clock(line_966_clock),
    .reset(line_966_reset),
    .valid(line_966_valid)
  );
  GEN_w1_line #(.COVER_INDEX(967)) line_967 (
    .clock(line_967_clock),
    .reset(line_967_reset),
    .valid(line_967_valid)
  );
  GEN_w1_line #(.COVER_INDEX(968)) line_968 (
    .clock(line_968_clock),
    .reset(line_968_reset),
    .valid(line_968_valid)
  );
  GEN_w1_line #(.COVER_INDEX(969)) line_969 (
    .clock(line_969_clock),
    .reset(line_969_reset),
    .valid(line_969_valid)
  );
  GEN_w1_line #(.COVER_INDEX(970)) line_970 (
    .clock(line_970_clock),
    .reset(line_970_reset),
    .valid(line_970_valid)
  );
  GEN_w1_line #(.COVER_INDEX(971)) line_971 (
    .clock(line_971_clock),
    .reset(line_971_reset),
    .valid(line_971_valid)
  );
  GEN_w1_line #(.COVER_INDEX(972)) line_972 (
    .clock(line_972_clock),
    .reset(line_972_reset),
    .valid(line_972_valid)
  );
  GEN_w1_line #(.COVER_INDEX(973)) line_973 (
    .clock(line_973_clock),
    .reset(line_973_reset),
    .valid(line_973_valid)
  );
  GEN_w1_line #(.COVER_INDEX(974)) line_974 (
    .clock(line_974_clock),
    .reset(line_974_reset),
    .valid(line_974_valid)
  );
  GEN_w1_line #(.COVER_INDEX(975)) line_975 (
    .clock(line_975_clock),
    .reset(line_975_reset),
    .valid(line_975_valid)
  );
  assign line_854_clock = clock;
  assign line_854_reset = reset;
  assign line_854_valid = 2'h0 == hitsVec_idx ^ line_854_valid_reg;
  assign line_855_clock = clock;
  assign line_855_reset = reset;
  assign line_855_valid = 2'h1 == hitsVec_idx ^ line_855_valid_reg;
  assign line_856_clock = clock;
  assign line_856_reset = reset;
  assign line_856_valid = 2'h2 == hitsVec_idx ^ line_856_valid_reg;
  assign line_857_clock = clock;
  assign line_857_reset = reset;
  assign line_857_valid = 2'h3 == hitsVec_idx ^ line_857_valid_reg;
  assign line_858_clock = clock;
  assign line_858_reset = reset;
  assign line_858_valid = 2'h0 == hitsVec_idx ^ line_858_valid_reg;
  assign line_859_clock = clock;
  assign line_859_reset = reset;
  assign line_859_valid = 2'h1 == hitsVec_idx ^ line_859_valid_reg;
  assign line_860_clock = clock;
  assign line_860_reset = reset;
  assign line_860_valid = 2'h2 == hitsVec_idx ^ line_860_valid_reg;
  assign line_861_clock = clock;
  assign line_861_reset = reset;
  assign line_861_valid = 2'h3 == hitsVec_idx ^ line_861_valid_reg;
  assign line_862_clock = clock;
  assign line_862_reset = reset;
  assign line_862_valid = io_ptw_resp_valid ^ line_862_valid_reg;
  assign line_863_clock = clock;
  assign line_863_reset = reset;
  assign line_863_valid = _T ^ line_863_valid_reg;
  assign line_864_clock = clock;
  assign line_864_reset = reset;
  assign line_864_valid = _T ^ line_864_valid_reg;
  assign line_865_clock = clock;
  assign line_865_reset = reset;
  assign line_865_valid = _T_2 ^ line_865_valid_reg;
  assign line_866_clock = clock;
  assign line_866_reset = reset;
  assign line_866_valid = _T_3 ^ line_866_valid_reg;
  assign line_867_clock = clock;
  assign line_867_reset = reset;
  assign line_867_valid = invalidate_refill ^ line_867_valid_reg;
  assign line_868_clock = clock;
  assign line_868_reset = reset;
  assign line_868_valid = r_superpage_repl_addr ^ line_868_valid_reg;
  assign line_869_clock = clock;
  assign line_869_reset = reset;
  assign line_869_valid = invalidate_refill ^ line_869_valid_reg;
  assign line_870_clock = clock;
  assign line_870_reset = reset;
  assign line_870_valid = _T_2 ^ line_870_valid_reg;
  assign line_871_clock = clock;
  assign line_871_reset = reset;
  assign line_871_valid = _T_5 ^ line_871_valid_reg;
  assign line_872_clock = clock;
  assign line_872_reset = reset;
  assign line_872_valid = _T_6 ^ line_872_valid_reg;
  assign line_873_clock = clock;
  assign line_873_reset = reset;
  assign line_873_valid = 2'h0 == idx ^ line_873_valid_reg;
  assign line_874_clock = clock;
  assign line_874_reset = reset;
  assign line_874_valid = 2'h1 == idx ^ line_874_valid_reg;
  assign line_875_clock = clock;
  assign line_875_reset = reset;
  assign line_875_valid = 2'h2 == idx ^ line_875_valid_reg;
  assign line_876_clock = clock;
  assign line_876_reset = reset;
  assign line_876_valid = 2'h3 == idx ^ line_876_valid_reg;
  assign line_877_clock = clock;
  assign line_877_reset = reset;
  assign line_877_valid = 2'h0 == idx ^ line_877_valid_reg;
  assign line_878_clock = clock;
  assign line_878_reset = reset;
  assign line_878_valid = 2'h1 == idx ^ line_878_valid_reg;
  assign line_879_clock = clock;
  assign line_879_reset = reset;
  assign line_879_valid = 2'h2 == idx ^ line_879_valid_reg;
  assign line_880_clock = clock;
  assign line_880_reset = reset;
  assign line_880_valid = 2'h3 == idx ^ line_880_valid_reg;
  assign line_881_clock = clock;
  assign line_881_reset = reset;
  assign line_881_valid = invalidate_refill ^ line_881_valid_reg;
  assign line_882_clock = clock;
  assign line_882_reset = reset;
  assign line_882_valid = waddr_1 ^ line_882_valid_reg;
  assign line_883_clock = clock;
  assign line_883_reset = reset;
  assign line_883_valid = _T_6 ^ line_883_valid_reg;
  assign line_884_clock = clock;
  assign line_884_reset = reset;
  assign line_884_valid = 2'h0 == idx ^ line_884_valid_reg;
  assign line_885_clock = clock;
  assign line_885_reset = reset;
  assign line_885_valid = 2'h1 == idx ^ line_885_valid_reg;
  assign line_886_clock = clock;
  assign line_886_reset = reset;
  assign line_886_valid = 2'h2 == idx ^ line_886_valid_reg;
  assign line_887_clock = clock;
  assign line_887_reset = reset;
  assign line_887_valid = 2'h3 == idx ^ line_887_valid_reg;
  assign line_888_clock = clock;
  assign line_888_reset = reset;
  assign line_888_valid = 2'h0 == idx ^ line_888_valid_reg;
  assign line_889_clock = clock;
  assign line_889_reset = reset;
  assign line_889_valid = 2'h1 == idx ^ line_889_valid_reg;
  assign line_890_clock = clock;
  assign line_890_reset = reset;
  assign line_890_valid = 2'h2 == idx ^ line_890_valid_reg;
  assign line_891_clock = clock;
  assign line_891_reset = reset;
  assign line_891_valid = 2'h3 == idx ^ line_891_valid_reg;
  assign line_892_clock = clock;
  assign line_892_reset = reset;
  assign line_892_valid = invalidate_refill ^ line_892_valid_reg;
  assign line_893_clock = clock;
  assign line_893_reset = reset;
  assign line_893_valid = 2'h0 == hitsVec_idx ^ line_893_valid_reg;
  assign line_894_clock = clock;
  assign line_894_reset = reset;
  assign line_894_valid = 2'h1 == hitsVec_idx ^ line_894_valid_reg;
  assign line_895_clock = clock;
  assign line_895_reset = reset;
  assign line_895_valid = 2'h2 == hitsVec_idx ^ line_895_valid_reg;
  assign line_896_clock = clock;
  assign line_896_reset = reset;
  assign line_896_valid = 2'h3 == hitsVec_idx ^ line_896_valid_reg;
  assign line_897_clock = clock;
  assign line_897_reset = reset;
  assign line_897_valid = 2'h0 == hitsVec_idx ^ line_897_valid_reg;
  assign line_898_clock = clock;
  assign line_898_reset = reset;
  assign line_898_valid = 2'h1 == hitsVec_idx ^ line_898_valid_reg;
  assign line_899_clock = clock;
  assign line_899_reset = reset;
  assign line_899_valid = 2'h2 == hitsVec_idx ^ line_899_valid_reg;
  assign line_900_clock = clock;
  assign line_900_reset = reset;
  assign line_900_valid = 2'h3 == hitsVec_idx ^ line_900_valid_reg;
  assign line_901_clock = clock;
  assign line_901_reset = reset;
  assign line_901_valid = _T_9 ^ line_901_valid_reg;
  assign line_902_clock = clock;
  assign line_902_reset = reset;
  assign line_902_valid = _T_10 ^ line_902_valid_reg;
  assign line_903_clock = clock;
  assign line_903_reset = reset;
  assign line_903_valid = _T_13 ^ line_903_valid_reg;
  assign line_904_clock = clock;
  assign line_904_reset = reset;
  assign line_904_valid = _T_17 ^ line_904_valid_reg;
  assign line_905_clock = clock;
  assign line_905_reset = reset;
  assign line_905_valid = _T_19 ^ line_905_valid_reg;
  assign line_906_clock = clock;
  assign line_906_reset = reset;
  assign line_906_valid = _invalidate_refill_T ^ line_906_valid_reg;
  assign line_907_clock = clock;
  assign line_907_reset = reset;
  assign line_907_valid = io_sfence_valid ^ line_907_valid_reg;
  assign line_908_clock = clock;
  assign line_908_reset = reset;
  assign line_908_valid = io_ptw_req_ready ^ line_908_valid_reg;
  assign line_909_clock = clock;
  assign line_909_reset = reset;
  assign line_909_valid = io_kill ^ line_909_valid_reg;
  assign line_910_clock = clock;
  assign line_910_reset = reset;
  assign line_910_valid = _T_22 ^ line_910_valid_reg;
  assign line_911_clock = clock;
  assign line_911_reset = reset;
  assign line_911_valid = io_ptw_resp_valid ^ line_911_valid_reg;
  assign line_912_clock = clock;
  assign line_912_reset = reset;
  assign line_912_valid = io_sfence_valid ^ line_912_valid_reg;
  assign line_913_clock = clock;
  assign line_913_reset = reset;
  assign line_913_valid = _T_28 ^ line_913_valid_reg;
  assign line_914_clock = clock;
  assign line_914_reset = reset;
  assign line_914_valid = _T_29 ^ line_914_valid_reg;
  assign line_915_clock = clock;
  assign line_915_reset = reset;
  assign line_915_valid = io_sfence_bits_rs1 ^ line_915_valid_reg;
  assign line_916_clock = clock;
  assign line_916_reset = reset;
  assign line_916_valid = _sector_hits_T_5 ^ line_916_valid_reg;
  assign line_917_clock = clock;
  assign line_917_reset = reset;
  assign line_917_valid = _GEN_0 ^ line_917_valid_reg;
  assign line_918_clock = clock;
  assign line_918_reset = reset;
  assign line_918_valid = _GEN_1 ^ line_918_valid_reg;
  assign line_919_clock = clock;
  assign line_919_reset = reset;
  assign line_919_valid = _GEN_2 ^ line_919_valid_reg;
  assign line_920_clock = clock;
  assign line_920_reset = reset;
  assign line_920_valid = _GEN_3 ^ line_920_valid_reg;
  assign line_921_clock = clock;
  assign line_921_reset = reset;
  assign line_921_valid = _T_147 ^ line_921_valid_reg;
  assign line_922_clock = clock;
  assign line_922_reset = reset;
  assign line_922_valid = sectored_entries_0_0_data_0[0] ^ line_922_valid_reg;
  assign line_923_clock = clock;
  assign line_923_reset = reset;
  assign line_923_valid = sectored_entries_0_0_data_1[0] ^ line_923_valid_reg;
  assign line_924_clock = clock;
  assign line_924_reset = reset;
  assign line_924_valid = sectored_entries_0_0_data_2[0] ^ line_924_valid_reg;
  assign line_925_clock = clock;
  assign line_925_reset = reset;
  assign line_925_valid = sectored_entries_0_0_data_3[0] ^ line_925_valid_reg;
  assign line_926_clock = clock;
  assign line_926_reset = reset;
  assign line_926_valid = io_sfence_bits_rs1 ^ line_926_valid_reg;
  assign line_927_clock = clock;
  assign line_927_reset = reset;
  assign line_927_valid = io_sfence_bits_rs2 ^ line_927_valid_reg;
  assign line_928_clock = clock;
  assign line_928_reset = reset;
  assign line_928_valid = _T_343 ^ line_928_valid_reg;
  assign line_929_clock = clock;
  assign line_929_reset = reset;
  assign line_929_valid = _T_346 ^ line_929_valid_reg;
  assign line_930_clock = clock;
  assign line_930_reset = reset;
  assign line_930_valid = _T_349 ^ line_930_valid_reg;
  assign line_931_clock = clock;
  assign line_931_reset = reset;
  assign line_931_valid = _T_352 ^ line_931_valid_reg;
  assign line_932_clock = clock;
  assign line_932_reset = reset;
  assign line_932_valid = io_sfence_bits_rs2 ^ line_932_valid_reg;
  assign line_933_clock = clock;
  assign line_933_reset = reset;
  assign line_933_valid = io_sfence_bits_rs1 ^ line_933_valid_reg;
  assign line_934_clock = clock;
  assign line_934_reset = reset;
  assign line_934_valid = _sector_hits_T_13 ^ line_934_valid_reg;
  assign line_935_clock = clock;
  assign line_935_reset = reset;
  assign line_935_valid = _GEN_0 ^ line_935_valid_reg;
  assign line_936_clock = clock;
  assign line_936_reset = reset;
  assign line_936_valid = _GEN_1 ^ line_936_valid_reg;
  assign line_937_clock = clock;
  assign line_937_reset = reset;
  assign line_937_valid = _GEN_2 ^ line_937_valid_reg;
  assign line_938_clock = clock;
  assign line_938_reset = reset;
  assign line_938_valid = _GEN_3 ^ line_938_valid_reg;
  assign line_939_clock = clock;
  assign line_939_reset = reset;
  assign line_939_valid = _T_568 ^ line_939_valid_reg;
  assign line_940_clock = clock;
  assign line_940_reset = reset;
  assign line_940_valid = sectored_entries_0_1_data_0[0] ^ line_940_valid_reg;
  assign line_941_clock = clock;
  assign line_941_reset = reset;
  assign line_941_valid = sectored_entries_0_1_data_1[0] ^ line_941_valid_reg;
  assign line_942_clock = clock;
  assign line_942_reset = reset;
  assign line_942_valid = sectored_entries_0_1_data_2[0] ^ line_942_valid_reg;
  assign line_943_clock = clock;
  assign line_943_reset = reset;
  assign line_943_valid = sectored_entries_0_1_data_3[0] ^ line_943_valid_reg;
  assign line_944_clock = clock;
  assign line_944_reset = reset;
  assign line_944_valid = io_sfence_bits_rs1 ^ line_944_valid_reg;
  assign line_945_clock = clock;
  assign line_945_reset = reset;
  assign line_945_valid = io_sfence_bits_rs2 ^ line_945_valid_reg;
  assign line_946_clock = clock;
  assign line_946_reset = reset;
  assign line_946_valid = _T_764 ^ line_946_valid_reg;
  assign line_947_clock = clock;
  assign line_947_reset = reset;
  assign line_947_valid = _T_767 ^ line_947_valid_reg;
  assign line_948_clock = clock;
  assign line_948_reset = reset;
  assign line_948_valid = _T_770 ^ line_948_valid_reg;
  assign line_949_clock = clock;
  assign line_949_reset = reset;
  assign line_949_valid = _T_773 ^ line_949_valid_reg;
  assign line_950_clock = clock;
  assign line_950_reset = reset;
  assign line_950_valid = io_sfence_bits_rs2 ^ line_950_valid_reg;
  assign line_951_clock = clock;
  assign line_951_reset = reset;
  assign line_951_valid = io_sfence_bits_rs1 ^ line_951_valid_reg;
  assign line_952_clock = clock;
  assign line_952_reset = reset;
  assign line_952_valid = superpage_hits_0 ^ line_952_valid_reg;
  assign line_953_clock = clock;
  assign line_953_reset = reset;
  assign line_953_valid = _T_891 ^ line_953_valid_reg;
  assign line_954_clock = clock;
  assign line_954_reset = reset;
  assign line_954_valid = superpage_entries_0_data_0[0] ^ line_954_valid_reg;
  assign line_955_clock = clock;
  assign line_955_reset = reset;
  assign line_955_valid = io_sfence_bits_rs1 ^ line_955_valid_reg;
  assign line_956_clock = clock;
  assign line_956_reset = reset;
  assign line_956_valid = io_sfence_bits_rs2 ^ line_956_valid_reg;
  assign line_957_clock = clock;
  assign line_957_reset = reset;
  assign line_957_valid = _T_943 ^ line_957_valid_reg;
  assign line_958_clock = clock;
  assign line_958_reset = reset;
  assign line_958_valid = io_sfence_bits_rs2 ^ line_958_valid_reg;
  assign line_959_clock = clock;
  assign line_959_reset = reset;
  assign line_959_valid = io_sfence_bits_rs1 ^ line_959_valid_reg;
  assign line_960_clock = clock;
  assign line_960_reset = reset;
  assign line_960_valid = superpage_hits_1 ^ line_960_valid_reg;
  assign line_961_clock = clock;
  assign line_961_reset = reset;
  assign line_961_valid = _T_989 ^ line_961_valid_reg;
  assign line_962_clock = clock;
  assign line_962_reset = reset;
  assign line_962_valid = superpage_entries_1_data_0[0] ^ line_962_valid_reg;
  assign line_963_clock = clock;
  assign line_963_reset = reset;
  assign line_963_valid = io_sfence_bits_rs1 ^ line_963_valid_reg;
  assign line_964_clock = clock;
  assign line_964_reset = reset;
  assign line_964_valid = io_sfence_bits_rs2 ^ line_964_valid_reg;
  assign line_965_clock = clock;
  assign line_965_reset = reset;
  assign line_965_valid = _T_1041 ^ line_965_valid_reg;
  assign line_966_clock = clock;
  assign line_966_reset = reset;
  assign line_966_valid = io_sfence_bits_rs2 ^ line_966_valid_reg;
  assign line_967_clock = clock;
  assign line_967_reset = reset;
  assign line_967_valid = io_sfence_bits_rs1 ^ line_967_valid_reg;
  assign line_968_clock = clock;
  assign line_968_reset = reset;
  assign line_968_valid = _hitsVec_T_56 ^ line_968_valid_reg;
  assign line_969_clock = clock;
  assign line_969_reset = reset;
  assign line_969_valid = _T_1087 ^ line_969_valid_reg;
  assign line_970_clock = clock;
  assign line_970_reset = reset;
  assign line_970_valid = special_entry_data_0[0] ^ line_970_valid_reg;
  assign line_971_clock = clock;
  assign line_971_reset = reset;
  assign line_971_valid = io_sfence_bits_rs1 ^ line_971_valid_reg;
  assign line_972_clock = clock;
  assign line_972_reset = reset;
  assign line_972_valid = io_sfence_bits_rs2 ^ line_972_valid_reg;
  assign line_973_clock = clock;
  assign line_973_reset = reset;
  assign line_973_valid = _T_1139 ^ line_973_valid_reg;
  assign line_974_clock = clock;
  assign line_974_reset = reset;
  assign line_974_valid = io_sfence_bits_rs2 ^ line_974_valid_reg;
  assign line_975_clock = clock;
  assign line_975_reset = reset;
  assign line_975_valid = _T_1433 ^ line_975_valid_reg;
  assign io_req_ready = state == 2'h0; // @[src/main/scala/rocket/TLB.scala 623:25]
  assign io_resp_miss = io_ptw_resp_valid | tlb_miss | multipleHits; // @[src/main/scala/rocket/TLB.scala 643:64]
  assign io_resp_paddr = {ppn,io_req_bits_vaddr[11:0]}; // @[src/main/scala/rocket/TLB.scala 644:23]
  assign io_resp_pf_inst = bad_va | |_io_resp_pf_inst_T; // @[src/main/scala/rocket/TLB.scala 627:29]
  assign io_resp_ae_inst = |_io_resp_ae_inst_T_1; // @[src/main/scala/rocket/TLB.scala 635:41]
  assign io_resp_cacheable = |_io_resp_cacheable_T; // @[src/main/scala/rocket/TLB.scala 640:41]
  assign io_ptw_req_valid = state == 2'h1; // @[src/main/scala/rocket/TLB.scala 652:29]
  assign io_ptw_req_bits_valid = ~io_kill; // @[src/main/scala/rocket/TLB.scala 653:28]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[src/main/scala/rocket/TLB.scala 654:29]
  assign io_ptw_req_bits_bits_need_gpa = r_need_gpa; // @[src/main/scala/rocket/TLB.scala 657:33]
  assign mpu_ppn_barrier_clock = clock;
  assign mpu_ppn_barrier_reset = reset;
  assign mpu_ppn_barrier_io_x_ppn = special_entry_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign entries_barrier_clock = clock;
  assign entries_barrier_reset = reset;
  assign entries_barrier_io_x_ppn = _GEN_330[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_u = _GEN_330[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_ae_ptw = _GEN_330[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_ae_final = _GEN_330[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_pf = _GEN_330[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_gf = _GEN_330[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_sx = _GEN_330[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_px = _GEN_330[7]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_io_x_c = _GEN_330[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_clock = clock;
  assign entries_barrier_1_reset = reset;
  assign entries_barrier_1_io_x_ppn = _GEN_334[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_u = _GEN_334[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_ae_ptw = _GEN_334[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_ae_final = _GEN_334[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_pf = _GEN_334[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_gf = _GEN_334[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_sx = _GEN_334[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_px = _GEN_334[7]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_1_io_x_c = _GEN_334[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_clock = clock;
  assign entries_barrier_2_reset = reset;
  assign entries_barrier_2_io_x_ppn = superpage_entries_0_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_u = superpage_entries_0_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_ae_ptw = superpage_entries_0_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_ae_final = superpage_entries_0_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_pf = superpage_entries_0_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_gf = superpage_entries_0_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_sx = superpage_entries_0_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_px = superpage_entries_0_data_0[7]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_2_io_x_c = superpage_entries_0_data_0[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_clock = clock;
  assign entries_barrier_3_reset = reset;
  assign entries_barrier_3_io_x_ppn = superpage_entries_1_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_u = superpage_entries_1_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_ae_ptw = superpage_entries_1_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_ae_final = superpage_entries_1_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_pf = superpage_entries_1_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_gf = superpage_entries_1_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_sx = superpage_entries_1_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_px = superpage_entries_1_data_0[7]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_3_io_x_c = superpage_entries_1_data_0[1]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_clock = clock;
  assign entries_barrier_4_reset = reset;
  assign entries_barrier_4_io_x_ppn = special_entry_data_0[41:22]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_u = special_entry_data_0[21]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_ae_ptw = special_entry_data_0[19]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_ae_final = special_entry_data_0[18]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_pf = special_entry_data_0[16]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_gf = special_entry_data_0[15]; // @[src/main/scala/rocket/TLB.scala 160:77]
  assign entries_barrier_4_io_x_sx = special_entry_data_0[13]; // @[src/main/scala/rocket/TLB.scala 160:77]
  always @(posedge clock) begin
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_0 <= _GEN_172;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_1 <= _GEN_173;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_2 <= _GEN_174;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_0_data_3 <= _GEN_175;
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_0 <= _GEN_366;
        end else begin
          sectored_entries_0_0_valid_0 <= _GEN_362;
        end
      end else begin
        sectored_entries_0_0_valid_0 <= _GEN_382;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_0 <= _GEN_228;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_1 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_1 <= _GEN_367;
        end else begin
          sectored_entries_0_0_valid_1 <= _GEN_363;
        end
      end else begin
        sectored_entries_0_0_valid_1 <= _GEN_383;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_1 <= _GEN_229;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_2 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_2 <= _GEN_368;
        end else begin
          sectored_entries_0_0_valid_2 <= _GEN_364;
        end
      end else begin
        sectored_entries_0_0_valid_2 <= _GEN_384;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_2 <= _GEN_230;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_0_valid_3 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_3[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_0_valid_3 <= _GEN_369;
        end else begin
          sectored_entries_0_0_valid_3 <= _GEN_365;
        end
      end else begin
        sectored_entries_0_0_valid_3 <= _GEN_385;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_0_valid_3 <= _GEN_231;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_0 <= _GEN_199;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_1 <= _GEN_200;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_2 <= _GEN_201;
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (!(io_ptw_resp_bits_level < 2'h2)) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (waddr_1) begin // @[src/main/scala/rocket/TLB.scala 478:84]
            sectored_entries_0_1_data_3 <= _GEN_202;
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_0 <= _GEN_398;
        end else begin
          sectored_entries_0_1_valid_0 <= _GEN_394;
        end
      end else begin
        sectored_entries_0_1_valid_0 <= _GEN_414;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_0 <= _GEN_239;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_1 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_1 <= _GEN_399;
        end else begin
          sectored_entries_0_1_valid_1 <= _GEN_395;
        end
      end else begin
        sectored_entries_0_1_valid_1 <= _GEN_415;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_1 <= _GEN_240;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_2 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_2 <= _GEN_400;
        end else begin
          sectored_entries_0_1_valid_2 <= _GEN_396;
        end
      end else begin
        sectored_entries_0_1_valid_2 <= _GEN_416;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_2 <= _GEN_241;
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      sectored_entries_0_1_valid_3 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_sector_hits_T_11[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          sectored_entries_0_1_valid_3 <= _GEN_401;
        end else begin
          sectored_entries_0_1_valid_3 <= _GEN_397;
        end
      end else begin
        sectored_entries_0_1_valid_3 <= _GEN_417;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        sectored_entries_0_1_valid_3 <= _GEN_242;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[src/main/scala/rocket/TLB.scala 203:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (~r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_0_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      superpage_entries_0_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_superpage_hits_T[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          superpage_entries_0_valid_0 <= _GEN_423;
        end else begin
          superpage_entries_0_valid_0 <= _GEN_422;
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_427;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        superpage_entries_0_valid_0 <= _GEN_221;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]}; // @[src/main/scala/rocket/TLB.scala 203:16]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
          end
        end
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        if (io_ptw_resp_bits_level < 2'h2) begin // @[src/main/scala/rocket/TLB.scala 468:58]
          if (r_superpage_repl_addr) begin // @[src/main/scala/rocket/TLB.scala 470:91]
            superpage_entries_1_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
          end
        end
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      superpage_entries_1_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_superpage_hits_T_14[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          superpage_entries_1_valid_0 <= _GEN_430;
        end else begin
          superpage_entries_1_valid_0 <= _GEN_429;
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_434;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (!(~io_ptw_resp_bits_homogeneous)) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        superpage_entries_1_valid_0 <= _GEN_226;
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_level <= io_ptw_resp_bits_level; // @[src/main/scala/rocket/TLB.scala 203:16]
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_tag_vpn <= r_refill_tag; // @[src/main/scala/rocket/TLB.scala 201:18]
      end
    end
    if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      if (~io_ptw_resp_bits_homogeneous) begin // @[src/main/scala/rocket/TLB.scala 466:70]
        special_entry_data_0 <= _special_entry_data_0_T; // @[src/main/scala/rocket/TLB.scala 207:15]
      end
    end
    if (multipleHits | reset) begin // @[src/main/scala/rocket/TLB.scala 722:41]
      special_entry_valid_0 <= 1'h0; // @[src/main/scala/rocket/TLB.scala 210:46]
    end else if (io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 708:19]
      if (io_sfence_bits_rs1) begin // @[src/main/scala/rocket/TLB.scala 713:42]
        if (_hitsVec_T_42[26:18] == 9'h0) begin // @[src/main/scala/rocket/TLB.scala 226:72]
          special_entry_valid_0 <= _GEN_437;
        end else begin
          special_entry_valid_0 <= _GEN_436;
        end
      end else begin
        special_entry_valid_0 <= _GEN_441;
      end
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 438:20]
      special_entry_valid_0 <= _GEN_253;
    end
    if (reset) begin // @[src/main/scala/rocket/TLB.scala 341:22]
      state <= 2'h0; // @[src/main/scala/rocket/TLB.scala 341:22]
    end else if (io_ptw_resp_valid) begin // @[src/main/scala/rocket/TLB.scala 703:30]
      state <= 2'h0; // @[src/main/scala/rocket/TLB.scala 704:13]
    end else if (state == 2'h2 & io_sfence_valid) begin // @[src/main/scala/rocket/TLB.scala 699:39]
      state <= 2'h3; // @[src/main/scala/rocket/TLB.scala 700:13]
    end else if (_invalidate_refill_T) begin // @[src/main/scala/rocket/TLB.scala 689:32]
      state <= _GEN_354;
    end else begin
      state <= _GEN_341;
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_refill_tag <= vpn; // @[src/main/scala/rocket/TLB.scala 671:20]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      if (&r_superpage_repl_addr_valids) begin // @[src/main/scala/rocket/TLB.scala 747:8]
        r_superpage_repl_addr <= state_reg_1;
      end else if (_r_superpage_repl_addr_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        r_superpage_repl_addr <= 1'h0;
      end else begin
        r_superpage_repl_addr <= 1'h1;
      end
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      if (&r_sectored_repl_addr_valids) begin // @[src/main/scala/rocket/TLB.scala 747:8]
        r_sectored_repl_addr <= state_vec_0;
      end else if (_r_sectored_repl_addr_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        r_sectored_repl_addr <= 1'h0;
      end else begin
        r_sectored_repl_addr <= 1'h1;
      end
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_sectored_hit_valid <= _T_10; // @[src/main/scala/rocket/TLB.scala 677:28]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_sectored_hit_bits <= state_vec_0_touch_way_sized; // @[src/main/scala/rocket/TLB.scala 678:27]
    end
    if (_T_18 & tlb_miss) begin // @[src/main/scala/rocket/TLB.scala 669:36]
      r_need_gpa <= tlb_hit_if_not_gpa_miss; // @[src/main/scala/rocket/TLB.scala 672:18]
    end
    line_854_valid_reg <= 2'h0 == hitsVec_idx;
    line_855_valid_reg <= 2'h1 == hitsVec_idx;
    line_856_valid_reg <= 2'h2 == hitsVec_idx;
    line_857_valid_reg <= 2'h3 == hitsVec_idx;
    line_858_valid_reg <= 2'h0 == hitsVec_idx;
    line_859_valid_reg <= 2'h1 == hitsVec_idx;
    line_860_valid_reg <= 2'h2 == hitsVec_idx;
    line_861_valid_reg <= 2'h3 == hitsVec_idx;
    line_862_valid_reg <= io_ptw_resp_valid;
    line_863_valid_reg <= _T;
    line_864_valid_reg <= _T;
    line_865_valid_reg <= _T_2;
    line_866_valid_reg <= _T_3;
    line_867_valid_reg <= invalidate_refill;
    line_868_valid_reg <= r_superpage_repl_addr;
    line_869_valid_reg <= invalidate_refill;
    line_870_valid_reg <= _T_2;
    line_871_valid_reg <= _T_5;
    line_872_valid_reg <= _T_6;
    line_873_valid_reg <= 2'h0 == idx;
    line_874_valid_reg <= 2'h1 == idx;
    line_875_valid_reg <= 2'h2 == idx;
    line_876_valid_reg <= 2'h3 == idx;
    line_877_valid_reg <= 2'h0 == idx;
    line_878_valid_reg <= 2'h1 == idx;
    line_879_valid_reg <= 2'h2 == idx;
    line_880_valid_reg <= 2'h3 == idx;
    line_881_valid_reg <= invalidate_refill;
    if (r_sectored_hit_valid) begin // @[src/main/scala/rocket/TLB.scala 477:22]
      line_882_valid_reg <= r_sectored_hit_bits;
    end else begin
      line_882_valid_reg <= r_sectored_repl_addr;
    end
    line_883_valid_reg <= _T_6;
    line_884_valid_reg <= 2'h0 == idx;
    line_885_valid_reg <= 2'h1 == idx;
    line_886_valid_reg <= 2'h2 == idx;
    line_887_valid_reg <= 2'h3 == idx;
    line_888_valid_reg <= 2'h0 == idx;
    line_889_valid_reg <= 2'h1 == idx;
    line_890_valid_reg <= 2'h2 == idx;
    line_891_valid_reg <= 2'h3 == idx;
    line_892_valid_reg <= invalidate_refill;
    line_893_valid_reg <= 2'h0 == hitsVec_idx;
    line_894_valid_reg <= 2'h1 == hitsVec_idx;
    line_895_valid_reg <= 2'h2 == hitsVec_idx;
    line_896_valid_reg <= 2'h3 == hitsVec_idx;
    line_897_valid_reg <= 2'h0 == hitsVec_idx;
    line_898_valid_reg <= 2'h1 == hitsVec_idx;
    line_899_valid_reg <= 2'h2 == hitsVec_idx;
    line_900_valid_reg <= 2'h3 == hitsVec_idx;
    if (reset) begin // @[src/main/scala/util/Replacement.scala 374:17]
      state_vec_0 <= 1'h0; // @[src/main/scala/util/Replacement.scala 374:17]
    end else if (io_req_valid & vm_enabled) begin // @[src/main/scala/rocket/TLB.scala 609:37]
      if (_T_10) begin // @[src/main/scala/rocket/TLB.scala 611:28]
        state_vec_0 <= _state_vec_0_T_1; // @[src/main/scala/util/Replacement.scala 377:20]
      end
    end
    if (reset) begin // @[src/main/scala/util/Replacement.scala 168:72]
      state_reg_1 <= 1'h0; // @[src/main/scala/util/Replacement.scala 168:72]
    end else if (io_req_valid & vm_enabled) begin // @[src/main/scala/rocket/TLB.scala 609:37]
      if (_T_13) begin // @[src/main/scala/rocket/TLB.scala 612:31]
        state_reg_1 <= _state_reg_T_1; // @[src/main/scala/util/Replacement.scala 172:15]
      end
    end
    line_901_valid_reg <= _T_9;
    line_902_valid_reg <= _T_10;
    line_903_valid_reg <= _T_13;
    line_904_valid_reg <= _T_17;
    line_905_valid_reg <= _T_19;
    line_906_valid_reg <= _invalidate_refill_T;
    line_907_valid_reg <= io_sfence_valid;
    line_908_valid_reg <= io_ptw_req_ready;
    line_909_valid_reg <= io_kill;
    line_910_valid_reg <= _T_22;
    line_911_valid_reg <= io_ptw_resp_valid;
    line_912_valid_reg <= io_sfence_valid;
    line_913_valid_reg <= _T_28;
    line_914_valid_reg <= _T_29;
    line_915_valid_reg <= io_sfence_bits_rs1;
    line_916_valid_reg <= _sector_hits_T_5;
    line_917_valid_reg <= _GEN_0;
    line_918_valid_reg <= _GEN_1;
    line_919_valid_reg <= _GEN_2;
    line_920_valid_reg <= _GEN_3;
    line_921_valid_reg <= _T_147;
    line_922_valid_reg <= sectored_entries_0_0_data_0[0];
    line_923_valid_reg <= sectored_entries_0_0_data_1[0];
    line_924_valid_reg <= sectored_entries_0_0_data_2[0];
    line_925_valid_reg <= sectored_entries_0_0_data_3[0];
    line_926_valid_reg <= io_sfence_bits_rs1;
    line_927_valid_reg <= io_sfence_bits_rs2;
    line_928_valid_reg <= _T_343;
    line_929_valid_reg <= _T_346;
    line_930_valid_reg <= _T_349;
    line_931_valid_reg <= _T_352;
    line_932_valid_reg <= io_sfence_bits_rs2;
    line_933_valid_reg <= io_sfence_bits_rs1;
    line_934_valid_reg <= _sector_hits_T_13;
    line_935_valid_reg <= _GEN_0;
    line_936_valid_reg <= _GEN_1;
    line_937_valid_reg <= _GEN_2;
    line_938_valid_reg <= _GEN_3;
    line_939_valid_reg <= _T_568;
    line_940_valid_reg <= sectored_entries_0_1_data_0[0];
    line_941_valid_reg <= sectored_entries_0_1_data_1[0];
    line_942_valid_reg <= sectored_entries_0_1_data_2[0];
    line_943_valid_reg <= sectored_entries_0_1_data_3[0];
    line_944_valid_reg <= io_sfence_bits_rs1;
    line_945_valid_reg <= io_sfence_bits_rs2;
    line_946_valid_reg <= _T_764;
    line_947_valid_reg <= _T_767;
    line_948_valid_reg <= _T_770;
    line_949_valid_reg <= _T_773;
    line_950_valid_reg <= io_sfence_bits_rs2;
    line_951_valid_reg <= io_sfence_bits_rs1;
    line_952_valid_reg <= superpage_hits_0;
    line_953_valid_reg <= _T_891;
    line_954_valid_reg <= superpage_entries_0_data_0[0];
    line_955_valid_reg <= io_sfence_bits_rs1;
    line_956_valid_reg <= io_sfence_bits_rs2;
    line_957_valid_reg <= _T_943;
    line_958_valid_reg <= io_sfence_bits_rs2;
    line_959_valid_reg <= io_sfence_bits_rs1;
    line_960_valid_reg <= superpage_hits_1;
    line_961_valid_reg <= _T_989;
    line_962_valid_reg <= superpage_entries_1_data_0[0];
    line_963_valid_reg <= io_sfence_bits_rs1;
    line_964_valid_reg <= io_sfence_bits_rs2;
    line_965_valid_reg <= _T_1041;
    line_966_valid_reg <= io_sfence_bits_rs2;
    line_967_valid_reg <= io_sfence_bits_rs1;
    line_968_valid_reg <= _hitsVec_T_56;
    line_969_valid_reg <= _T_1087;
    line_970_valid_reg <= special_entry_data_0[0];
    line_971_valid_reg <= io_sfence_bits_rs1;
    line_972_valid_reg <= io_sfence_bits_rs2;
    line_973_valid_reg <= _T_1139;
    line_974_valid_reg <= io_sfence_bits_rs2;
    line_975_valid_reg <= _T_1433;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~reset & ~(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TLB.scala:709 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"
            ); // @[src/main/scala/rocket/TLB.scala 709:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_0_tag_vpn = _RAND_0[26:0];
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_0_data_0 = _RAND_1[41:0];
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_0_data_1 = _RAND_2[41:0];
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_0_data_2 = _RAND_3[41:0];
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_0_data_3 = _RAND_4[41:0];
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_0_valid_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_0_valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_0_valid_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_0_valid_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_0_1_tag_vpn = _RAND_9[26:0];
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_0_1_data_0 = _RAND_10[41:0];
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_0_1_data_1 = _RAND_11[41:0];
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_0_1_data_2 = _RAND_12[41:0];
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_0_1_data_3 = _RAND_13[41:0];
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_0_1_valid_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_0_1_valid_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_0_1_valid_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_0_1_valid_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  superpage_entries_0_tag_vpn = _RAND_19[26:0];
  _RAND_20 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_20[41:0];
  _RAND_21 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  superpage_entries_1_tag_vpn = _RAND_23[26:0];
  _RAND_24 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_24[41:0];
  _RAND_25 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  special_entry_level = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  special_entry_tag_vpn = _RAND_27[26:0];
  _RAND_28 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_28[41:0];
  _RAND_29 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  r_refill_tag = _RAND_31[26:0];
  _RAND_32 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_sectored_hit_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_sectored_hit_bits = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_need_gpa = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_854_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_855_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_856_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_857_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_858_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_859_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_860_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_861_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_862_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_863_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_864_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_865_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_866_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_867_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_868_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_869_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_870_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_871_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_872_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_873_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_874_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_875_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_876_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_877_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_878_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_879_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_880_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_881_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_882_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_883_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_884_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_885_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_886_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_887_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_888_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_889_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_890_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_891_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_892_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_893_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_894_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_895_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_896_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_897_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_898_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_899_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_900_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  state_vec_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  state_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_901_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_902_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_903_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_904_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_905_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_906_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_907_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_908_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_909_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_910_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_911_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_912_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_913_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_914_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_915_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_916_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_917_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_918_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_919_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_920_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_921_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_922_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_923_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_924_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_925_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_926_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  line_927_valid_reg = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  line_928_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  line_929_valid_reg = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  line_930_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  line_931_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_932_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_933_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_934_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_935_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_936_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_937_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_938_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_939_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_940_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_941_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_942_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_943_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_944_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_945_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_946_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_947_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_948_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_949_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_950_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_951_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_952_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_953_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_954_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_955_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_956_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_957_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_958_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_959_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_960_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_961_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_962_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_963_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_964_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_965_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_966_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_967_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_968_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_969_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_970_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_971_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_972_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_973_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_974_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_975_valid_reg = _RAND_160[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (io_sfence_valid & ~reset) begin
      assert(~io_sfence_bits_rs1 | io_sfence_bits_addr[38:12] == vpn); // @[src/main/scala/rocket/TLB.scala 709:13]
    end
  end
endmodule
module Frontend(
  input         clock,
  input         reset,
  input         auto_icache_master_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_icache_master_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_icache_master_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_icache_master_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_icache_master_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_icache_master_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_icache_master_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_icache_master_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         io_cpu_might_request, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_req_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [39:0] io_cpu_req_bits_pc, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_req_bits_speculative, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_sfence_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_sfence_bits_rs1, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_sfence_bits_rs2, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [38:0] io_cpu_sfence_bits_addr, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_resp_ready, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_cpu_resp_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output [39:0] io_cpu_resp_bits_pc, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output [31:0] io_cpu_resp_bits_data, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_cpu_resp_bits_xcpt_pf_inst, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_cpu_resp_bits_xcpt_ae_inst, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_cpu_resp_bits_replay, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_btb_update_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_bht_update_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_flush_icache, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output [39:0] io_cpu_npc, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_cpu_progress, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_req_ready, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_ptw_req_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_ptw_req_bits_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output [26:0] io_ptw_req_bits_bits_addr, // @[src/main/scala/rocket/Frontend.scala 81:14]
  output        io_ptw_req_bits_bits_need_gpa, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_valid, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_ae_ptw, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_ae_final, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pf, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [43:0] io_ptw_resp_bits_pte_ppn, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_d, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_a, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_g, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_u, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_x, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_w, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_r, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_pte_v, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [1:0]  io_ptw_resp_bits_level, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input         io_ptw_resp_bits_homogeneous, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [3:0]  io_ptw_ptbr_mode, // @[src/main/scala/rocket/Frontend.scala 81:14]
  input  [1:0]  io_ptw_status_prv // @[src/main/scala/rocket/Frontend.scala 81:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  icache_clock; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_reset; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_auto_master_out_a_ready; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_auto_master_out_a_valid; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [31:0] icache_auto_master_out_a_bits_address; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_auto_master_out_d_valid; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [2:0] icache_auto_master_out_d_bits_opcode; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [2:0] icache_auto_master_out_d_bits_size; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [63:0] icache_auto_master_out_d_bits_data; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_auto_master_out_d_bits_corrupt; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_req_ready; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_req_valid; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [38:0] icache_io_req_bits_addr; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [31:0] icache_io_s1_paddr; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_s1_kill; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_s2_kill; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_resp_valid; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire [31:0] icache_io_resp_bits_data; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_resp_bits_ae; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  icache_io_invalidate; // @[src/main/scala/rocket/Frontend.scala 66:26]
  wire  fq_clock; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_reset; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_enq_ready; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_enq_valid; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire [39:0] fq_io_enq_bits_pc; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire [31:0] fq_io_enq_bits_data; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_enq_bits_xcpt_pf_inst; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_enq_bits_xcpt_ae_inst; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_enq_bits_replay; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_deq_ready; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_deq_valid; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire [39:0] fq_io_deq_bits_pc; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire [31:0] fq_io_deq_bits_data; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_deq_bits_xcpt_pf_inst; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_deq_bits_xcpt_ae_inst; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  fq_io_deq_bits_replay; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire [4:0] fq_io_mask; // @[src/main/scala/rocket/Frontend.scala 87:64]
  wire  tlb_clock; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_reset; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_req_ready; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_req_valid; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [1:0] tlb_io_req_bits_prv; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_resp_miss; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [31:0] tlb_io_resp_paddr; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_resp_pf_inst; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_resp_ae_inst; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_resp_cacheable; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_sfence_valid; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_sfence_bits_rs1; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_sfence_bits_rs2; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_req_ready; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_req_valid; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_req_bits_valid; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_valid; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pf; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [43:0] tlb_io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  tlb_io_kill; // @[src/main/scala/rocket/Frontend.scala 101:19]
  wire  _T_9 = ~reset; // @[src/main/scala/rocket/Frontend.scala 92:9]
  wire  line_976_clock;
  wire  line_976_reset;
  wire  line_976_valid;
  reg  line_976_valid_reg;
  wire  _T_10 = ~(~(io_cpu_req_valid | io_cpu_sfence_valid | io_cpu_flush_icache | io_cpu_bht_update_valid |
    io_cpu_btb_update_valid) | io_cpu_might_request); // @[src/main/scala/rocket/Frontend.scala 92:9]
  wire  line_977_clock;
  wire  line_977_reset;
  wire  line_977_valid;
  reg  line_977_valid_reg;
  reg  s1_valid; // @[src/main/scala/rocket/Frontend.scala 103:21]
  reg  s2_valid; // @[src/main/scala/rocket/Frontend.scala 104:25]
  wire  _s0_fq_has_space_T_4 = ~s1_valid; // @[src/main/scala/rocket/Frontend.scala 107:45]
  wire  _s0_fq_has_space_T_5 = ~s2_valid; // @[src/main/scala/rocket/Frontend.scala 107:58]
  wire  _s0_fq_has_space_T_7 = ~fq_io_mask[3] & (~s1_valid | ~s2_valid); // @[src/main/scala/rocket/Frontend.scala 107:41]
  wire  _s0_fq_has_space_T_8 = ~fq_io_mask[2] | _s0_fq_has_space_T_7; // @[src/main/scala/rocket/Frontend.scala 106:40]
  wire  _s0_fq_has_space_T_14 = ~fq_io_mask[4] & (_s0_fq_has_space_T_4 & _s0_fq_has_space_T_5); // @[src/main/scala/rocket/Frontend.scala 108:41]
  wire  s0_fq_has_space = _s0_fq_has_space_T_8 | _s0_fq_has_space_T_14; // @[src/main/scala/rocket/Frontend.scala 107:70]
  wire  s0_valid = io_cpu_req_valid | s0_fq_has_space; // @[src/main/scala/rocket/Frontend.scala 109:35]
  reg [39:0] s1_pc; // @[src/main/scala/rocket/Frontend.scala 111:18]
  reg  s1_speculative; // @[src/main/scala/rocket/Frontend.scala 112:27]
  reg [39:0] s2_pc; // @[src/main/scala/rocket/Frontend.scala 113:22]
  reg  s2_tlb_resp_miss; // @[src/main/scala/rocket/Frontend.scala 117:24]
  reg  s2_tlb_resp_pf_inst; // @[src/main/scala/rocket/Frontend.scala 117:24]
  reg  s2_tlb_resp_ae_inst; // @[src/main/scala/rocket/Frontend.scala 117:24]
  reg  s2_tlb_resp_cacheable; // @[src/main/scala/rocket/Frontend.scala 117:24]
  wire  s2_xcpt = s2_tlb_resp_ae_inst | s2_tlb_resp_pf_inst; // @[src/main/scala/rocket/Frontend.scala 118:37]
  reg  s2_speculative; // @[src/main/scala/rocket/Frontend.scala 119:31]
  wire [39:0] _s1_base_pc_T = ~s1_pc; // @[src/main/scala/rocket/Frontend.scala 124:22]
  wire [39:0] _s1_base_pc_T_1 = _s1_base_pc_T | 40'h3; // @[src/main/scala/rocket/Frontend.scala 124:29]
  wire [39:0] s1_base_pc = ~_s1_base_pc_T_1; // @[src/main/scala/rocket/Frontend.scala 124:20]
  wire [39:0] ntpc = s1_base_pc + 40'h4; // @[src/main/scala/rocket/Frontend.scala 125:25]
  wire  _s2_replay_T = fq_io_enq_ready & fq_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  s2_replay_REG; // @[src/main/scala/rocket/Frontend.scala 130:56]
  wire  s2_replay = s2_valid & ~_s2_replay_T | s2_replay_REG; // @[src/main/scala/rocket/Frontend.scala 130:46]
  wire [39:0] npc = s2_replay ? s2_pc : ntpc; // @[src/main/scala/rocket/Frontend.scala 131:16]
  wire  s0_speculative = s1_speculative | s2_valid & ~s2_speculative; // @[src/main/scala/rocket/Frontend.scala 137:41]
  wire  _T_11 = ~s2_replay; // @[src/main/scala/rocket/Frontend.scala 143:9]
  wire  line_978_clock;
  wire  line_978_reset;
  wire  line_978_valid;
  reg  line_978_valid_reg;
  wire  _GEN_11 = ~s2_replay & ~io_cpu_req_valid; // @[src/main/scala/rocket/Frontend.scala 142:12 143:21 144:14]
  reg [1:0] recent_progress_counter; // @[src/main/scala/rocket/Frontend.scala 151:40]
  wire  recent_progress = recent_progress_counter > 2'h0; // @[src/main/scala/rocket/Frontend.scala 152:49]
  wire  _T_12 = io_ptw_req_ready & io_ptw_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_13 = _T_12 & recent_progress; // @[src/main/scala/rocket/Frontend.scala 153:24]
  wire  line_979_clock;
  wire  line_979_reset;
  wire  line_979_valid;
  reg  line_979_valid_reg;
  wire [1:0] _recent_progress_counter_T_1 = recent_progress_counter - 2'h1; // @[src/main/scala/rocket/Frontend.scala 153:97]
  wire  line_980_clock;
  wire  line_980_reset;
  wire  line_980_valid;
  reg  line_980_valid_reg;
  wire  s2_kill_speculative_tlb_refill = s2_speculative & ~recent_progress; // @[src/main/scala/rocket/Frontend.scala 156:55]
  reg  fq_io_enq_valid_REG; // @[src/main/scala/rocket/Frontend.scala 180:29]
  wire  _fq_io_enq_valid_T_1 = s2_kill_speculative_tlb_refill & s2_tlb_resp_miss; // @[src/main/scala/rocket/Frontend.scala 180:112]
  wire [39:0] _io_cpu_npc_T = io_cpu_req_valid ? io_cpu_req_bits_pc : npc; // @[src/main/scala/rocket/Frontend.scala 182:28]
  wire [39:0] _io_cpu_npc_T_1 = ~_io_cpu_npc_T; // @[src/main/scala/rocket/Frontend.scala 377:29]
  wire [39:0] _io_cpu_npc_T_2 = _io_cpu_npc_T_1 | 40'h1; // @[src/main/scala/rocket/Frontend.scala 377:33]
  wire  line_981_clock;
  wire  line_981_reset;
  wire  line_981_valid;
  reg  line_981_valid_reg;
  wire  _T_21 = icache_io_resp_valid & icache_io_resp_bits_ae; // @[src/main/scala/rocket/Frontend.scala 191:30]
  wire  line_982_clock;
  wire  line_982_reset;
  wire  line_982_valid;
  reg  line_982_valid_reg;
  wire  line_983_clock;
  wire  line_983_reset;
  wire  line_983_valid;
  reg  line_983_valid_reg;
  ICache icache ( // @[src/main/scala/rocket/Frontend.scala 66:26]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_master_out_a_ready(icache_auto_master_out_a_ready),
    .auto_master_out_a_valid(icache_auto_master_out_a_valid),
    .auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),
    .auto_master_out_d_valid(icache_auto_master_out_d_valid),
    .auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),
    .auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),
    .auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),
    .auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),
    .io_req_ready(icache_io_req_ready),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_paddr(icache_io_s1_paddr),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_ae(icache_io_resp_bits_ae),
    .io_invalidate(icache_io_invalidate)
  );
  ShiftQueue fq ( // @[src/main/scala/rocket/Frontend.scala 87:64]
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_pc(fq_io_enq_bits_pc),
    .io_enq_bits_data(fq_io_enq_bits_data),
    .io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),
    .io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
    .io_enq_bits_replay(fq_io_enq_bits_replay),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_pc(fq_io_deq_bits_pc),
    .io_deq_bits_data(fq_io_deq_bits_data),
    .io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),
    .io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
    .io_deq_bits_replay(fq_io_deq_bits_replay),
    .io_mask(fq_io_mask)
  );
  TLB_1 tlb ( // @[src/main/scala/rocket/Frontend.scala 101:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_prv(tlb_io_req_bits_prv),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_req_bits_bits_need_gpa(tlb_io_ptw_req_bits_bits_need_gpa),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_ptw(tlb_io_ptw_resp_bits_ae_ptw),
    .io_ptw_resp_bits_ae_final(tlb_io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pf(tlb_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_kill(tlb_io_kill)
  );
  GEN_w1_line #(.COVER_INDEX(976)) line_976 (
    .clock(line_976_clock),
    .reset(line_976_reset),
    .valid(line_976_valid)
  );
  GEN_w1_line #(.COVER_INDEX(977)) line_977 (
    .clock(line_977_clock),
    .reset(line_977_reset),
    .valid(line_977_valid)
  );
  GEN_w1_line #(.COVER_INDEX(978)) line_978 (
    .clock(line_978_clock),
    .reset(line_978_reset),
    .valid(line_978_valid)
  );
  GEN_w1_line #(.COVER_INDEX(979)) line_979 (
    .clock(line_979_clock),
    .reset(line_979_reset),
    .valid(line_979_valid)
  );
  GEN_w1_line #(.COVER_INDEX(980)) line_980 (
    .clock(line_980_clock),
    .reset(line_980_reset),
    .valid(line_980_valid)
  );
  GEN_w1_line #(.COVER_INDEX(981)) line_981 (
    .clock(line_981_clock),
    .reset(line_981_reset),
    .valid(line_981_valid)
  );
  GEN_w1_line #(.COVER_INDEX(982)) line_982 (
    .clock(line_982_clock),
    .reset(line_982_reset),
    .valid(line_982_valid)
  );
  GEN_w1_line #(.COVER_INDEX(983)) line_983 (
    .clock(line_983_clock),
    .reset(line_983_reset),
    .valid(line_983_valid)
  );
  assign line_976_clock = clock;
  assign line_976_reset = reset;
  assign line_976_valid = _T_9 ^ line_976_valid_reg;
  assign line_977_clock = clock;
  assign line_977_reset = reset;
  assign line_977_valid = _T_10 ^ line_977_valid_reg;
  assign line_978_clock = clock;
  assign line_978_reset = reset;
  assign line_978_valid = _T_11 ^ line_978_valid_reg;
  assign line_979_clock = clock;
  assign line_979_reset = reset;
  assign line_979_valid = _T_13 ^ line_979_valid_reg;
  assign line_980_clock = clock;
  assign line_980_reset = reset;
  assign line_980_valid = io_cpu_progress ^ line_980_valid_reg;
  assign line_981_clock = clock;
  assign line_981_reset = reset;
  assign line_981_valid = _T_9 ^ line_981_valid_reg;
  assign line_982_clock = clock;
  assign line_982_reset = reset;
  assign line_982_valid = _T_21 ^ line_982_valid_reg;
  assign line_983_clock = clock;
  assign line_983_reset = reset;
  assign line_983_valid = io_cpu_req_valid ^ line_983_valid_reg;
  assign auto_icache_master_out_a_valid = icache_auto_master_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_icache_master_out_a_bits_address = icache_auto_master_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign io_cpu_resp_valid = fq_io_deq_valid; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_resp_bits_data = fq_io_deq_bits_data; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_resp_bits_xcpt_pf_inst = fq_io_deq_bits_xcpt_pf_inst; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign io_cpu_npc = ~_io_cpu_npc_T_2; // @[src/main/scala/rocket/Frontend.scala 377:27]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign io_ptw_req_bits_valid = tlb_io_ptw_req_bits_valid; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign io_ptw_req_bits_bits_need_gpa = tlb_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign icache_clock = clock; // @[src/main/scala/rocket/Frontend.scala 97:16]
  assign icache_reset = reset;
  assign icache_auto_master_out_a_ready = auto_icache_master_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_auto_master_out_d_valid = auto_icache_master_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_auto_master_out_d_bits_opcode = auto_icache_master_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_auto_master_out_d_bits_size = auto_icache_master_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_auto_master_out_d_bits_data = auto_icache_master_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_auto_master_out_d_bits_corrupt = auto_icache_master_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign icache_io_req_valid = io_cpu_req_valid | s0_fq_has_space; // @[src/main/scala/rocket/Frontend.scala 109:35]
  assign icache_io_req_bits_addr = io_cpu_npc[38:0]; // @[src/main/scala/rocket/Frontend.scala 170:27]
  assign icache_io_s1_paddr = tlb_io_resp_paddr; // @[src/main/scala/rocket/Frontend.scala 172:22]
  assign icache_io_s1_kill = io_cpu_req_valid | tlb_io_resp_miss | s2_replay; // @[src/main/scala/rocket/Frontend.scala 174:56]
  assign icache_io_s2_kill = s2_speculative & ~s2_tlb_resp_cacheable | s2_xcpt; // @[src/main/scala/rocket/Frontend.scala 176:71]
  assign icache_io_invalidate = io_cpu_flush_icache; // @[src/main/scala/rocket/Frontend.scala 171:24]
  assign fq_clock = clock;
  assign fq_reset = reset | io_cpu_req_valid; // @[src/main/scala/rocket/Frontend.scala 87:35]
  assign fq_io_enq_valid = fq_io_enq_valid_REG & s2_valid & (icache_io_resp_valid | s2_kill_speculative_tlb_refill &
    s2_tlb_resp_miss | ~s2_tlb_resp_miss & icache_io_s2_kill); // @[src/main/scala/rocket/Frontend.scala 180:52]
  assign fq_io_enq_bits_pc = s2_pc; // @[src/main/scala/rocket/Frontend.scala 181:21]
  assign fq_io_enq_bits_data = icache_io_resp_bits_data; // @[src/main/scala/rocket/Frontend.scala 184:23]
  assign fq_io_enq_bits_xcpt_pf_inst = s2_tlb_resp_pf_inst; // @[src/main/scala/rocket/Frontend.scala 189:23]
  assign fq_io_enq_bits_xcpt_ae_inst = icache_io_resp_valid & icache_io_resp_bits_ae | s2_tlb_resp_ae_inst; // @[src/main/scala/rocket/Frontend.scala 189:23 191:{57,87}]
  assign fq_io_enq_bits_replay = icache_io_s2_kill & ~icache_io_resp_valid & ~s2_xcpt | _fq_io_enq_valid_T_1; // @[src/main/scala/rocket/Frontend.scala 186:115]
  assign fq_io_deq_ready = io_cpu_resp_ready; // @[src/main/scala/rocket/Frontend.scala 346:15]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid & _T_11; // @[src/main/scala/rocket/Frontend.scala 159:32]
  assign tlb_io_req_bits_vaddr = s1_pc; // @[src/main/scala/rocket/Frontend.scala 161:25]
  assign tlb_io_req_bits_prv = io_ptw_status_prv; // @[src/main/scala/rocket/Frontend.scala 164:23]
  assign tlb_io_sfence_valid = io_cpu_sfence_valid; // @[src/main/scala/rocket/Frontend.scala 166:17]
  assign tlb_io_sfence_bits_rs1 = io_cpu_sfence_bits_rs1; // @[src/main/scala/rocket/Frontend.scala 166:17]
  assign tlb_io_sfence_bits_rs2 = io_cpu_sfence_bits_rs2; // @[src/main/scala/rocket/Frontend.scala 166:17]
  assign tlb_io_sfence_bits_addr = io_cpu_sfence_bits_addr; // @[src/main/scala/rocket/Frontend.scala 166:17]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_ae_ptw = io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_ae_final = io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pf = io_ptw_resp_bits_pf; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[src/main/scala/rocket/Frontend.scala 158:10]
  assign tlb_io_kill = _s0_fq_has_space_T_5 | s2_kill_speculative_tlb_refill; // @[src/main/scala/rocket/Frontend.scala 167:28]
  always @(posedge clock) begin
    line_976_valid_reg <= _T_9;
    line_977_valid_reg <= _T_10;
    s1_valid <= io_cpu_req_valid | s0_fq_has_space; // @[src/main/scala/rocket/Frontend.scala 109:35]
    if (reset) begin // @[src/main/scala/rocket/Frontend.scala 104:25]
      s2_valid <= 1'h0; // @[src/main/scala/rocket/Frontend.scala 104:25]
    end else begin
      s2_valid <= _GEN_11;
    end
    s1_pc <= io_cpu_npc; // @[src/main/scala/rocket/Frontend.scala 133:9]
    if (io_cpu_req_valid) begin // @[src/main/scala/rocket/Frontend.scala 139:24]
      s1_speculative <= io_cpu_req_bits_speculative;
    end else if (s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 139:75]
      s1_speculative <= s2_speculative;
    end else begin
      s1_speculative <= s0_speculative;
    end
    if (reset) begin // @[src/main/scala/rocket/Frontend.scala 113:22]
      s2_pc <= 40'h10000000; // @[src/main/scala/rocket/Frontend.scala 113:22]
    end else if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_pc <= s1_pc; // @[src/main/scala/rocket/Frontend.scala 145:11]
    end
    if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_tlb_resp_miss <= tlb_io_resp_miss; // @[src/main/scala/rocket/Frontend.scala 147:17]
    end
    if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_tlb_resp_pf_inst <= tlb_io_resp_pf_inst; // @[src/main/scala/rocket/Frontend.scala 147:17]
    end
    if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst; // @[src/main/scala/rocket/Frontend.scala 147:17]
    end
    if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_tlb_resp_cacheable <= tlb_io_resp_cacheable; // @[src/main/scala/rocket/Frontend.scala 147:17]
    end
    if (reset) begin // @[src/main/scala/rocket/Frontend.scala 119:31]
      s2_speculative <= 1'h0; // @[src/main/scala/rocket/Frontend.scala 119:31]
    end else if (~s2_replay) begin // @[src/main/scala/rocket/Frontend.scala 143:21]
      s2_speculative <= s1_speculative; // @[src/main/scala/rocket/Frontend.scala 146:20]
    end
    s2_replay_REG <= reset | s2_replay & ~s0_valid; // @[src/main/scala/rocket/Frontend.scala 130:{56,56,56}]
    line_978_valid_reg <= _T_11;
    if (reset) begin // @[src/main/scala/rocket/Frontend.scala 151:40]
      recent_progress_counter <= 2'h3; // @[src/main/scala/rocket/Frontend.scala 151:40]
    end else if (io_cpu_progress) begin // @[src/main/scala/rocket/Frontend.scala 154:25]
      recent_progress_counter <= 2'h3; // @[src/main/scala/rocket/Frontend.scala 154:51]
    end else if (_T_12 & recent_progress) begin // @[src/main/scala/rocket/Frontend.scala 153:44]
      recent_progress_counter <= _recent_progress_counter_T_1; // @[src/main/scala/rocket/Frontend.scala 153:70]
    end
    line_979_valid_reg <= _T_13;
    line_980_valid_reg <= io_cpu_progress;
    fq_io_enq_valid_REG <= s1_valid; // @[src/main/scala/rocket/Frontend.scala 180:29]
    line_981_valid_reg <= _T_9;
    line_982_valid_reg <= _T_21;
    line_983_valid_reg <= io_cpu_req_valid;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_cpu_req_valid | io_cpu_sfence_valid | io_cpu_flush_icache | io_cpu_bht_update_valid |
          io_cpu_btb_update_valid) | io_cpu_might_request)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Frontend.scala:92 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n"
            ); // @[src/main/scala/rocket/Frontend.scala 92:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_976_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_977_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s1_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s2_valid = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  s1_pc = _RAND_4[39:0];
  _RAND_5 = {1{`RANDOM}};
  s1_speculative = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  s2_pc = _RAND_6[39:0];
  _RAND_7 = {1{`RANDOM}};
  s2_tlb_resp_miss = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s2_tlb_resp_pf_inst = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s2_tlb_resp_ae_inst = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  s2_tlb_resp_cacheable = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  s2_speculative = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s2_replay_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_978_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  recent_progress_counter = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  line_979_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_980_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  fq_io_enq_valid_REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_981_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_982_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_983_valid_reg = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_cpu_req_valid | io_cpu_sfence_valid | io_cpu_flush_icache | io_cpu_bht_update_valid |
        io_cpu_btb_update_valid) | io_cpu_might_request); // @[src/main/scala/rocket/Frontend.scala 92:9]
    end
    //
    if (_T_9) begin
      assert(1'h1); // @[src/main/scala/rocket/Frontend.scala 190:9]
    end
  end
endmodule
module TLWidthWidget_8(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLFragmenter_1(
  input   clock,
  input   reset
);
endmodule
module TLWidthWidget_9(
  input   clock,
  input   reset
);
endmodule
module TLBuffer_6(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_size = auto_out_b_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_source = auto_out_b_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_c_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_e_ready = auto_out_e_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_a_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_valid = auto_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_source = auto_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_c_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_d_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_valid = auto_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_e_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLBuffer_7(
  input   clock,
  input   reset
);
endmodule
module HellaCacheArbiter(
  input         clock,
  input         reset,
  output        io_requestor_0_req_ready, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_requestor_0_req_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [39:0] io_requestor_0_req_bits_addr, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_requestor_0_s1_kill, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_0_s2_nack, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_0_resp_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [63:0] io_requestor_0_resp_bits_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_0_s2_xcpt_ae_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_req_ready, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_requestor_1_req_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [39:0] io_requestor_1_req_bits_addr, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [6:0]  io_requestor_1_req_bits_tag, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [4:0]  io_requestor_1_req_bits_cmd, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [1:0]  io_requestor_1_req_bits_size, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_requestor_1_req_bits_signed, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [1:0]  io_requestor_1_req_bits_dprv, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_requestor_1_s1_kill, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [63:0] io_requestor_1_s1_data_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_nack, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_resp_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [6:0]  io_requestor_1_resp_bits_tag, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [63:0] io_requestor_1_resp_bits_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_resp_bits_replay, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_resp_bits_has_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [63:0] io_requestor_1_resp_bits_data_word_bypass, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_replay_next, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_ma_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_ma_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_pf_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_pf_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_ae_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_s2_xcpt_ae_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_ordered, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_perf_release, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_requestor_1_perf_grant, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_req_ready, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_mem_req_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [39:0] io_mem_req_bits_addr, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [6:0]  io_mem_req_bits_tag, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [4:0]  io_mem_req_bits_cmd, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [1:0]  io_mem_req_bits_size, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_mem_req_bits_signed, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [1:0]  io_mem_req_bits_dprv, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_mem_req_bits_phys, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output        io_mem_s1_kill, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  output [63:0] io_mem_s1_data_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_nack, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_resp_valid, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [6:0]  io_mem_resp_bits_tag, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [63:0] io_mem_resp_bits_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_resp_bits_replay, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_resp_bits_has_data, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input  [63:0] io_mem_resp_bits_data_word_bypass, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_replay_next, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_ma_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_ma_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_pf_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_pf_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_ae_ld, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_s2_xcpt_ae_st, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_ordered, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_perf_release, // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
  input         io_mem_perf_grant // @[src/main/scala/rocket/HellaCacheArbiter.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  s1_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 20:20]
  reg  s2_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 21:24]
  wire [7:0] _io_mem_req_bits_tag_T = {io_requestor_1_req_bits_tag,1'h1}; // @[src/main/scala/rocket/HellaCacheArbiter.scala 34:35]
  wire  line_984_clock;
  wire  line_984_reset;
  wire  line_984_valid;
  reg  line_984_valid_reg;
  wire [7:0] _GEN_4 = io_requestor_0_req_valid ? 8'h0 : _io_mem_req_bits_tag_T; // @[src/main/scala/rocket/HellaCacheArbiter.scala 50:26 34:{29,29}]
  wire  _T = ~s1_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 51:21]
  wire  line_985_clock;
  wire  line_985_reset;
  wire  line_985_valid;
  reg  line_985_valid_reg;
  wire  _T_1 = ~s2_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 52:21]
  wire  line_986_clock;
  wire  line_986_reset;
  wire  line_986_valid;
  reg  line_986_valid_reg;
  wire  tag_hit = ~io_mem_resp_bits_tag[0]; // @[src/main/scala/rocket/HellaCacheArbiter.scala 60:57]
  GEN_w1_line #(.COVER_INDEX(984)) line_984 (
    .clock(line_984_clock),
    .reset(line_984_reset),
    .valid(line_984_valid)
  );
  GEN_w1_line #(.COVER_INDEX(985)) line_985 (
    .clock(line_985_clock),
    .reset(line_985_reset),
    .valid(line_985_valid)
  );
  GEN_w1_line #(.COVER_INDEX(986)) line_986 (
    .clock(line_986_clock),
    .reset(line_986_reset),
    .valid(line_986_valid)
  );
  assign line_984_clock = clock;
  assign line_984_reset = reset;
  assign line_984_valid = io_requestor_0_req_valid ^ line_984_valid_reg;
  assign line_985_clock = clock;
  assign line_985_reset = reset;
  assign line_985_valid = _T ^ line_985_valid_reg;
  assign line_986_clock = clock;
  assign line_986_reset = reset;
  assign line_986_valid = _T_1 ^ line_986_valid_reg;
  assign io_requestor_0_req_ready = io_mem_req_ready; // @[src/main/scala/rocket/HellaCacheArbiter.scala 26:31]
  assign io_requestor_0_s2_nack = io_mem_s2_nack & _T_1; // @[src/main/scala/rocket/HellaCacheArbiter.scala 67:49]
  assign io_requestor_0_resp_valid = io_mem_resp_valid & tag_hit; // @[src/main/scala/rocket/HellaCacheArbiter.scala 61:39]
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data; // @[src/main/scala/rocket/HellaCacheArbiter.scala 72:17]
  assign io_requestor_0_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_req_ready = io_requestor_0_req_ready & ~io_requestor_0_req_valid; // @[src/main/scala/rocket/HellaCacheArbiter.scala 28:64]
  assign io_requestor_1_s2_nack = io_mem_s2_nack & s2_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 67:49]
  assign io_requestor_1_resp_valid = io_mem_resp_valid & io_mem_resp_bits_tag[0]; // @[src/main/scala/rocket/HellaCacheArbiter.scala 61:39]
  assign io_requestor_1_resp_bits_tag = {{1'd0}, io_mem_resp_bits_tag[6:1]}; // @[src/main/scala/rocket/HellaCacheArbiter.scala 73:21]
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data; // @[src/main/scala/rocket/HellaCacheArbiter.scala 72:17]
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay; // @[src/main/scala/rocket/HellaCacheArbiter.scala 72:17]
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data; // @[src/main/scala/rocket/HellaCacheArbiter.scala 72:17]
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass; // @[src/main/scala/rocket/HellaCacheArbiter.scala 72:17]
  assign io_requestor_1_replay_next = io_mem_replay_next; // @[src/main/scala/rocket/HellaCacheArbiter.scala 75:35]
  assign io_requestor_1_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st; // @[src/main/scala/rocket/HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_ordered = io_mem_ordered; // @[src/main/scala/rocket/HellaCacheArbiter.scala 65:31]
  assign io_requestor_1_perf_release = io_mem_perf_release; // @[src/main/scala/rocket/HellaCacheArbiter.scala 66:28]
  assign io_requestor_1_perf_grant = io_mem_perf_grant; // @[src/main/scala/rocket/HellaCacheArbiter.scala 66:28]
  assign io_mem_req_valid = io_requestor_0_req_valid | io_requestor_1_req_valid; // @[src/main/scala/rocket/HellaCacheArbiter.scala 25:63]
  assign io_mem_req_bits_addr = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_req_bits_tag = _GEN_4[6:0];
  assign io_mem_req_bits_cmd = io_requestor_0_req_valid ? 5'h0 : io_requestor_1_req_bits_cmd; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_req_bits_size = io_requestor_0_req_valid ? 2'h3 : io_requestor_1_req_bits_size; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_req_bits_signed = io_requestor_0_req_valid ? 1'h0 : io_requestor_1_req_bits_signed; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_req_bits_dprv = io_requestor_0_req_valid ? 2'h1 : io_requestor_1_req_bits_dprv; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_req_bits_phys = io_requestor_0_req_valid; // @[src/main/scala/rocket/HellaCacheArbiter.scala 33:{25,25} 50:26]
  assign io_mem_s1_kill = ~s1_id ? io_requestor_0_s1_kill : io_requestor_1_s1_kill; // @[src/main/scala/rocket/HellaCacheArbiter.scala 38:{24,24} 51:30]
  assign io_mem_s1_data_data = ~s1_id ? 64'h0 : io_requestor_1_s1_data_data; // @[src/main/scala/rocket/HellaCacheArbiter.scala 39:{24,24} 51:30]
  always @(posedge clock) begin
    if (io_requestor_0_req_valid) begin // @[src/main/scala/rocket/HellaCacheArbiter.scala 50:26]
      s1_id <= 1'h0; // @[src/main/scala/rocket/HellaCacheArbiter.scala 35:15]
    end else begin
      s1_id <= 1'h1; // @[src/main/scala/rocket/HellaCacheArbiter.scala 35:15]
    end
    s2_id <= s1_id; // @[src/main/scala/rocket/HellaCacheArbiter.scala 21:24]
    line_984_valid_reg <= io_requestor_0_req_valid;
    line_985_valid_reg <= _T;
    line_986_valid_reg <= _T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_id = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_id = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_984_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_985_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_986_valid_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [26:0] io_in_0_bits_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_0_bits_bits_need_gpa, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_bits_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input  [26:0] io_in_1_bits_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_in_1_bits_bits_need_gpa, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output [26:0] io_out_bits_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_out_bits_bits_need_gpa, // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 134:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  line_987_clock;
  wire  line_987_reset;
  wire  line_987_valid;
  reg  line_987_valid_reg;
  wire  grant_1 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  GEN_w1_line #(.COVER_INDEX(987)) line_987 (
    .clock(line_987_clock),
    .reset(line_987_reset),
    .valid(line_987_valid)
  );
  assign line_987_clock = clock;
  assign line_987_reset = reset;
  assign line_987_valid = io_in_0_valid ^ line_987_valid_reg;
  assign io_in_0_ready = io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 147:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 148:31]
  assign io_out_bits_valid = io_in_0_valid | io_in_1_bits_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_bits_addr = io_in_0_valid ? io_in_0_bits_bits_addr : io_in_1_bits_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_out_bits_bits_need_gpa = io_in_0_valid ? io_in_0_bits_bits_need_gpa : io_in_1_bits_bits_need_gpa; // @[src/main/scala/chisel3/util/Arbiter.scala 137:15 139:26 141:19]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 136:13 139:26 140:17]
  always @(posedge clock) begin
    line_987_valid_reg <= io_in_0_valid;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_987_valid_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OptimizationBarrier_18(
  input        clock,
  input        reset,
  input  [2:0] io_x, // @[src/main/scala/util/package.scala 260:18]
  output [2:0] io_y // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y = io_x; // @[src/main/scala/util/package.scala 264:12]
endmodule
module OptimizationBarrier_19(
  input         clock,
  input         reset,
  input  [43:0] io_x_ppn, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_d, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_a, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_g, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_u, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_x, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_w, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_r, // @[src/main/scala/util/package.scala 260:18]
  input         io_x_v, // @[src/main/scala/util/package.scala 260:18]
  output [43:0] io_y_ppn, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_d, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_a, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_g, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_u, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_x, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_w, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_r, // @[src/main/scala/util/package.scala 260:18]
  output        io_y_v // @[src/main/scala/util/package.scala 260:18]
);
  assign io_y_ppn = io_x_ppn; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_d = io_x_d; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_a = io_x_a; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_g = io_x_g; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_u = io_x_u; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_x = io_x_x; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_w = io_x_w; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_r = io_x_r; // @[src/main/scala/util/package.scala 264:12]
  assign io_y_v = io_x_v; // @[src/main/scala/util/package.scala 264:12]
endmodule
module PTW(
  input         clock,
  input         reset,
  output        io_requestor_0_req_ready, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_requestor_0_req_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [26:0] io_requestor_0_req_bits_bits_addr, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_requestor_0_req_bits_bits_need_gpa, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_ae_ptw, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_ae_final, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pf, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [43:0] io_requestor_0_resp_bits_pte_ppn, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_d, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_a, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_g, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_u, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_x, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_w, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_r, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_pte_v, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [1:0]  io_requestor_0_resp_bits_level, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_resp_bits_homogeneous, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [3:0]  io_requestor_0_ptbr_mode, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_status_mxr, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_0_status_sum, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_req_ready, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_requestor_1_req_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_requestor_1_req_bits_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [26:0] io_requestor_1_req_bits_bits_addr, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_requestor_1_req_bits_bits_need_gpa, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_ae_ptw, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_ae_final, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pf, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [43:0] io_requestor_1_resp_bits_pte_ppn, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_d, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_a, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_g, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_u, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_x, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_w, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_r, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_pte_v, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [1:0]  io_requestor_1_resp_bits_level, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_requestor_1_resp_bits_homogeneous, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [3:0]  io_requestor_1_ptbr_mode, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [1:0]  io_requestor_1_status_prv, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_mem_req_ready, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_mem_req_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  output [39:0] io_mem_req_bits_addr, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_mem_s1_kill, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_mem_s2_nack, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_mem_resp_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [63:0] io_mem_resp_bits_data, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_mem_s2_xcpt_ae_ld, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [3:0]  io_dpath_ptbr_mode, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [43:0] io_dpath_ptbr_ppn, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_dpath_sfence_valid, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_dpath_sfence_bits_rs1, // @[src/main/scala/rocket/PTW.scala 220:14]
  input  [1:0]  io_dpath_status_prv, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_dpath_status_mxr, // @[src/main/scala/rocket/PTW.scala 220:14]
  input         io_dpath_status_sum, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_dpath_perf_l2hit, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_dpath_perf_pte_miss, // @[src/main/scala/rocket/PTW.scala 220:14]
  output        io_dpath_perf_pte_hit // @[src/main/scala/rocket/PTW.scala 220:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
`endif // RANDOMIZE_REG_INIT
  wire  arb_clock; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_reset; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_0_ready; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_0_valid; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire [26:0] arb_io_in_0_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_0_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_1_ready; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_1_valid; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_1_bits_valid; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire [26:0] arb_io_in_1_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_in_1_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_out_ready; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_out_valid; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_out_bits_valid; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire [26:0] arb_io_out_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_out_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  arb_io_chosen; // @[src/main/scala/rocket/PTW.scala 236:19]
  wire  state_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  state_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [2:0] state_barrier_io_x; // @[src/main/scala/util/package.scala 259:25]
  wire [2:0] state_barrier_io_y; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_clock; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_reset; // @[src/main/scala/util/package.scala 259:25]
  wire [43:0] r_pte_barrier_io_x_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_d; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_a; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_g; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_u; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_x; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_w; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_r; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_x_v; // @[src/main/scala/util/package.scala 259:25]
  wire [43:0] r_pte_barrier_io_y_ppn; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_d; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_a; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_g; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_u; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_x; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_w; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_r; // @[src/main/scala/util/package.scala 259:25]
  wire  r_pte_barrier_io_y_v; // @[src/main/scala/util/package.scala 259:25]
  reg [2:0] state; // @[src/main/scala/rocket/PTW.scala 233:22]
  reg  l2_refill; // @[src/main/scala/rocket/PTW.scala 410:26]
  reg  resp_valid_0; // @[src/main/scala/rocket/PTW.scala 242:27]
  reg  resp_valid_1; // @[src/main/scala/rocket/PTW.scala 242:27]
  wire  _clock_en_T = state != 3'h0; // @[src/main/scala/rocket/PTW.scala 244:24]
  reg  invalidated; // @[src/main/scala/rocket/PTW.scala 251:24]
  reg [1:0] count; // @[src/main/scala/rocket/PTW.scala 259:18]
  reg  resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 260:24]
  reg  resp_ae_final; // @[src/main/scala/rocket/PTW.scala 261:26]
  reg  resp_pf; // @[src/main/scala/rocket/PTW.scala 262:20]
  reg [26:0] r_req_addr; // @[src/main/scala/rocket/PTW.scala 270:18]
  reg  r_req_need_gpa; // @[src/main/scala/rocket/PTW.scala 270:18]
  reg  r_req_dest; // @[src/main/scala/rocket/PTW.scala 272:23]
  reg [43:0] r_pte_ppn; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_d; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_a; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_g; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_u; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_x; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_w; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_r; // @[src/main/scala/rocket/PTW.scala 275:18]
  reg  r_pte_v; // @[src/main/scala/rocket/PTW.scala 275:18]
  wire [43:0] vpn = {{17'd0}, r_req_addr}; // @[src/main/scala/rocket/PTW.scala 291:16]
  reg  mem_resp_valid; // @[src/main/scala/rocket/PTW.scala 293:31]
  reg [63:0] mem_resp_data; // @[src/main/scala/rocket/PTW.scala 294:30]
  wire  tmp_v = mem_resp_data[0]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_r = mem_resp_data[1]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_w = mem_resp_data[2]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_x = mem_resp_data[3]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_u = mem_resp_data[4]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_g = mem_resp_data[5]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_a = mem_resp_data[6]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire  tmp_d = mem_resp_data[7]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire [43:0] tmp_ppn = mem_resp_data[53:10]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire [9:0] tmp_reserved_for_future = mem_resp_data[63:54]; // @[src/main/scala/rocket/PTW.scala 305:37]
  wire [26:0] _res_ppn_T_4 = {{7'd0}, tmp_ppn[19:0]}; // @[src/main/scala/rocket/PTW.scala 307:19]
  wire  _T_1 = tmp_r | tmp_w | tmp_x; // @[src/main/scala/rocket/PTW.scala 308:26]
  wire  line_988_clock;
  wire  line_988_reset;
  wire  line_988_valid;
  reg  line_988_valid_reg;
  wire  _T_5 = count <= 2'h0 & tmp_ppn[17:9] != 9'h0; // @[src/main/scala/rocket/PTW.scala 311:28]
  wire  line_989_clock;
  wire  line_989_reset;
  wire  line_989_valid;
  reg  line_989_valid_reg;
  wire  _GEN_66 = count <= 2'h0 & tmp_ppn[17:9] != 9'h0 ? 1'h0 : tmp_v; // @[src/main/scala/rocket/PTW.scala 311:{106,114} 306:26]
  wire  _T_9 = count <= 2'h1 & tmp_ppn[8:0] != 9'h0; // @[src/main/scala/rocket/PTW.scala 311:28]
  wire  line_990_clock;
  wire  line_990_reset;
  wire  line_990_valid;
  reg  line_990_valid_reg;
  wire  _GEN_67 = count <= 2'h1 & tmp_ppn[8:0] != 9'h0 ? 1'h0 : _GEN_66; // @[src/main/scala/rocket/PTW.scala 311:{106,114}]
  wire  pte_v = tmp_r | tmp_w | tmp_x ? _GEN_67 : tmp_v; // @[src/main/scala/rocket/PTW.scala 306:26 308:36]
  wire  invalid_paddr = tmp_ppn[43:20] != 24'h0; // @[src/main/scala/rocket/PTW.scala 313:93]
  wire  _traverse_T_13 = pte_v & ~tmp_r & ~tmp_w & ~tmp_x & ~tmp_d & ~tmp_a & ~tmp_u & tmp_reserved_for_future == 10'h0; // @[src/main/scala/rocket/PTW.scala 139:69]
  wire  _traverse_T_16 = count < 2'h2; // @[src/main/scala/rocket/PTW.scala 316:57]
  wire  traverse = _traverse_T_13 & ~invalid_paddr & count < 2'h2; // @[src/main/scala/rocket/PTW.scala 316:48]
  wire [8:0] pte_addr_vpn_idxs_0 = vpn[26:18]; // @[src/main/scala/rocket/PTW.scala 321:48]
  wire [8:0] pte_addr_vpn_idxs_1 = vpn[17:9]; // @[src/main/scala/rocket/PTW.scala 321:48]
  wire [8:0] pte_addr_vpn_idxs_2 = vpn[8:0]; // @[src/main/scala/rocket/PTW.scala 321:48]
  wire [8:0] _pte_addr_vpn_idx_T_1 = count == 2'h1 ? pte_addr_vpn_idxs_1 : pte_addr_vpn_idxs_0; // @[src/main/scala/util/package.scala 33:76]
  wire  _pte_addr_vpn_idx_T_2 = count == 2'h2; // @[src/main/scala/util/package.scala 33:86]
  wire [8:0] _pte_addr_vpn_idx_T_3 = count == 2'h2 ? pte_addr_vpn_idxs_2 : _pte_addr_vpn_idx_T_1; // @[src/main/scala/util/package.scala 33:76]
  wire [8:0] pte_addr_vpn_idx = count == 2'h3 ? pte_addr_vpn_idxs_2 : _pte_addr_vpn_idx_T_3; // @[src/main/scala/util/package.scala 33:76]
  wire [52:0] _pte_addr_raw_pte_addr_T = {r_pte_ppn, 9'h0}; // @[src/main/scala/rocket/PTW.scala 325:36]
  wire [52:0] _GEN_272 = {{44'd0}, pte_addr_vpn_idx}; // @[src/main/scala/rocket/PTW.scala 325:52]
  wire [52:0] _pte_addr_raw_pte_addr_T_1 = _pte_addr_raw_pte_addr_T | _GEN_272; // @[src/main/scala/rocket/PTW.scala 325:52]
  wire [55:0] pte_addr_raw_pte_addr = {_pte_addr_raw_pte_addr_T_1, 3'h0}; // @[src/main/scala/rocket/PTW.scala 325:63]
  wire [31:0] pte_addr = pte_addr_raw_pte_addr[31:0]; // @[src/main/scala/rocket/PTW.scala 329:23]
  reg  state_reg; // @[src/main/scala/util/Replacement.scala 168:72]
  reg [1:0] valid; // @[src/main/scala/rocket/PTW.scala 364:24]
  reg [31:0] tags__0; // @[src/main/scala/rocket/PTW.scala 365:19]
  reg [31:0] tags__1; // @[src/main/scala/rocket/PTW.scala 365:19]
  reg [19:0] data__0; // @[src/main/scala/rocket/PTW.scala 367:19]
  reg [19:0] data__1; // @[src/main/scala/rocket/PTW.scala 367:19]
  wire [32:0] tag = {1'h0,pte_addr}; // @[src/main/scala/rocket/PTW.scala 376:15]
  wire [32:0] _GEN_273 = {{1'd0}, tags__0}; // @[src/main/scala/rocket/PTW.scala 378:27]
  wire  _hits_T = _GEN_273 == tag; // @[src/main/scala/rocket/PTW.scala 378:27]
  wire [32:0] _GEN_274 = {{1'd0}, tags__1}; // @[src/main/scala/rocket/PTW.scala 378:27]
  wire  _hits_T_1 = _GEN_274 == tag; // @[src/main/scala/rocket/PTW.scala 378:27]
  wire [1:0] _hits_T_2 = {_hits_T_1,_hits_T}; // @[src/main/scala/util/package.scala 37:27]
  wire [1:0] hits = _hits_T_2 & valid; // @[src/main/scala/rocket/PTW.scala 378:43]
  wire  _hit_T = |hits; // @[src/main/scala/rocket/PTW.scala 379:20]
  wire  pte_cache_hit = |hits & _traverse_T_16; // @[src/main/scala/rocket/PTW.scala 379:24]
  wire  _T_22 = mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated; // @[src/main/scala/rocket/PTW.scala 381:65]
  wire  line_991_clock;
  wire  line_991_reset;
  wire  line_991_valid;
  reg  line_991_valid_reg;
  wire [1:0] _r_T_2 = ~valid; // @[src/main/scala/rocket/PTW.scala 382:57]
  wire  _r_T_5 = _r_T_2[0] ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  r = &valid ? state_reg : _r_T_5; // @[src/main/scala/rocket/PTW.scala 382:18]
  wire [1:0] _valid_T = 2'h1 << r; // @[src/main/scala/chisel3/util/OneHot.scala 58:35]
  wire [1:0] _valid_T_1 = valid | _valid_T; // @[src/main/scala/rocket/PTW.scala 383:22]
  wire  _GEN_3 = ~r; // @[src/main/scala/rocket/PTW.scala 384:15]
  wire  line_992_clock;
  wire  line_992_reset;
  wire  line_992_valid;
  reg  line_992_valid_reg;
  wire  line_993_clock;
  wire  line_993_reset;
  wire  line_993_valid;
  reg  line_993_valid_reg;
  wire  line_994_clock;
  wire  line_994_reset;
  wire  line_994_valid;
  reg  line_994_valid_reg;
  wire [43:0] pte_ppn = {{17'd0}, _res_ppn_T_4}; // @[src/main/scala/rocket/PTW.scala 306:26 307:13]
  wire  line_995_clock;
  wire  line_995_reset;
  wire  line_995_valid;
  reg  line_995_valid_reg;
  wire  _T_23 = state == 3'h1; // @[src/main/scala/rocket/PTW.scala 389:24]
  wire  _T_24 = pte_cache_hit & state == 3'h1; // @[src/main/scala/rocket/PTW.scala 389:15]
  wire  line_996_clock;
  wire  line_996_reset;
  wire  line_996_valid;
  reg  line_996_valid_reg;
  wire  state_reg_touch_way_sized_1 = hits[1]; // @[src/main/scala/chisel3/util/CircuitMath.scala 28:8]
  wire  _state_reg_T_3 = ~state_reg_touch_way_sized_1; // @[src/main/scala/util/Replacement.scala 218:7]
  wire  _T_29 = io_dpath_sfence_valid & ~io_dpath_sfence_bits_rs1; // @[src/main/scala/rocket/PTW.scala 390:33]
  wire  line_997_clock;
  wire  line_997_reset;
  wire  line_997_valid;
  reg  line_997_valid_reg;
  wire [19:0] _T_40 = hits[0] ? data__0 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] _T_41 = state_reg_touch_way_sized_1 ? data__1 : 20'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [19:0] pte_cache_data = _T_40 | _T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  line_998_clock;
  wire  line_998_reset;
  wire  line_998_valid;
  reg  line_998_valid_reg;
  reg  pte_hit; // @[src/main/scala/rocket/PTW.scala 404:24]
  wire  _T_74 = ~reset; // @[src/main/scala/rocket/PTW.scala 407:9]
  wire  line_999_clock;
  wire  line_999_reset;
  wire  line_999_valid;
  reg  line_999_valid_reg;
  wire  _T_75 = ~(~(io_dpath_perf_l2hit & (io_dpath_perf_pte_miss | io_dpath_perf_pte_hit))); // @[src/main/scala/rocket/PTW.scala 407:9]
  wire  line_1000_clock;
  wire  line_1000_reset;
  wire  line_1000_valid;
  reg  line_1000_valid_reg;
  wire [55:0] _pmaPgLevelHomogeneous_T = {r_pte_ppn, 12'h0}; // @[src/main/scala/rocket/PTW.scala 555:88]
  wire [55:0] _pmaPgLevelHomogeneous_T_1 = _pmaPgLevelHomogeneous_T ^ 56'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [56:0] _pmaPgLevelHomogeneous_T_2 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_1)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [56:0] _pmaPgLevelHomogeneous_T_4 = $signed(_pmaPgLevelHomogeneous_T_2) & -57'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  pmaPgLevelHomogeneous_0 = $signed(_pmaPgLevelHomogeneous_T_4) == 57'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire [55:0] _pmaPgLevelHomogeneous_T_21 = _pmaPgLevelHomogeneous_T ^ 56'h10000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [56:0] _pmaPgLevelHomogeneous_T_22 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_21)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [56:0] _pmaPgLevelHomogeneous_T_24 = $signed(_pmaPgLevelHomogeneous_T_22) & -57'sh10000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  _pmaPgLevelHomogeneous_T_25 = $signed(_pmaPgLevelHomogeneous_T_24) == 57'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  wire  pmaPgLevelHomogeneous_2 = _pmaPgLevelHomogeneous_T_25 | pmaPgLevelHomogeneous_0; // @[src/main/scala/rocket/TLBPermissions.scala 101:65]
  wire  _pmaHomogeneous_T_1 = count == 2'h1 ? pmaPgLevelHomogeneous_0 : pmaPgLevelHomogeneous_0; // @[src/main/scala/util/package.scala 33:76]
  wire  _pmaHomogeneous_T_3 = count == 2'h2 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_1; // @[src/main/scala/util/package.scala 33:76]
  wire  pmaHomogeneous = count == 2'h3 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_3; // @[src/main/scala/util/package.scala 33:76]
  wire  _T_76 = 3'h0 == state; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  line_1001_clock;
  wire  line_1001_reset;
  wire  line_1001_valid;
  reg  line_1001_valid_reg;
  wire  _T_77 = arb_io_out_ready & arb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1002_clock;
  wire  line_1002_reset;
  wire  line_1002_valid;
  reg  line_1002_valid_reg;
  wire [2:0] _next_state_T = arb_io_out_bits_valid ? 3'h1 : 3'h0; // @[src/main/scala/rocket/PTW.scala 604:26]
  wire  line_1003_clock;
  wire  line_1003_reset;
  wire  line_1003_valid;
  reg  line_1003_valid_reg;
  wire  _T_82 = ~(~arb_io_out_bits_bits_need_gpa); // @[src/main/scala/rocket/PTW.scala 622:15]
  wire  line_1004_clock;
  wire  line_1004_reset;
  wire  line_1004_valid;
  reg  line_1004_valid_reg;
  wire [2:0] _GEN_98 = _T_77 ? _next_state_T : state; // @[src/main/scala/rocket/PTW.scala 596:30 604:20 590:31]
  wire  _GEN_105 = _T_77 ? 1'h0 : resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 596:30 612:21 260:24]
  wire  _GEN_106 = _T_77 ? 1'h0 : resp_ae_final; // @[src/main/scala/rocket/PTW.scala 596:30 613:23 261:26]
  wire  _GEN_107 = _T_77 ? 1'h0 : resp_pf; // @[src/main/scala/rocket/PTW.scala 596:30 614:17 262:20]
  wire  line_1005_clock;
  wire  line_1005_reset;
  wire  line_1005_valid;
  reg  line_1005_valid_reg;
  wire  _T_83 = 3'h1 == state; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  line_1006_clock;
  wire  line_1006_reset;
  wire  line_1006_valid;
  reg  line_1006_valid_reg;
  wire  line_1007_clock;
  wire  line_1007_reset;
  wire  line_1007_valid;
  reg  line_1007_valid_reg;
  wire [1:0] _count_T_2 = count + 2'h1; // @[src/main/scala/rocket/PTW.scala 637:24]
  wire  line_1008_clock;
  wire  line_1008_reset;
  wire  line_1008_valid;
  reg  line_1008_valid_reg;
  wire [2:0] _next_state_T_1 = io_mem_req_ready ? 3'h2 : 3'h1; // @[src/main/scala/rocket/PTW.scala 640:26]
  wire [2:0] _GEN_119 = pte_cache_hit ? state : _next_state_T_1; // @[src/main/scala/rocket/PTW.scala 590:31 636:34 640:20]
  wire  line_1009_clock;
  wire  line_1009_reset;
  wire  line_1009_valid;
  reg  line_1009_valid_reg;
  wire  _T_86 = 3'h2 == state; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  line_1010_clock;
  wire  line_1010_reset;
  wire  line_1010_valid;
  reg  line_1010_valid_reg;
  wire  line_1011_clock;
  wire  line_1011_reset;
  wire  line_1011_valid;
  reg  line_1011_valid_reg;
  wire  _T_87 = 3'h4 == state; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  line_1012_clock;
  wire  line_1012_reset;
  wire  line_1012_valid;
  reg  line_1012_valid_reg;
  wire  line_1013_clock;
  wire  line_1013_reset;
  wire  line_1013_valid;
  reg  line_1013_valid_reg;
  wire  _GEN_27 = ~r_req_dest; // @[src/main/scala/rocket/PTW.scala 653:32]
  wire  line_1014_clock;
  wire  line_1014_reset;
  wire  line_1014_valid;
  reg  line_1014_valid_reg;
  wire  line_1015_clock;
  wire  line_1015_reset;
  wire  line_1015_valid;
  reg  line_1015_valid_reg;
  wire  _GEN_128 = io_mem_s2_xcpt_ae_ld | resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 650:35 651:21 260:24]
  wire [2:0] _GEN_129 = io_mem_s2_xcpt_ae_ld ? 3'h0 : 3'h5; // @[src/main/scala/rocket/PTW.scala 648:18 650:35 652:20]
  wire  _GEN_130 = io_mem_s2_xcpt_ae_ld & _GEN_27; // @[src/main/scala/rocket/PTW.scala 242:27 650:35]
  wire  _GEN_131 = io_mem_s2_xcpt_ae_ld & r_req_dest; // @[src/main/scala/rocket/PTW.scala 242:27 650:35]
  wire  line_1016_clock;
  wire  line_1016_reset;
  wire  line_1016_valid;
  reg  line_1016_valid_reg;
  wire  _T_90 = 3'h7 == state; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  line_1017_clock;
  wire  line_1017_reset;
  wire  line_1017_valid;
  reg  line_1017_valid_reg;
  wire  line_1018_clock;
  wire  line_1018_reset;
  wire  line_1018_valid;
  reg  line_1018_valid_reg;
  wire  line_1019_clock;
  wire  line_1019_reset;
  wire  line_1019_valid;
  reg  line_1019_valid_reg;
  wire  _T_93 = ~pmaHomogeneous; // @[src/main/scala/rocket/PTW.scala 659:13]
  wire  line_1020_clock;
  wire  line_1020_reset;
  wire  line_1020_valid;
  reg  line_1020_valid_reg;
  wire [1:0] _GEN_134 = ~pmaHomogeneous ? 2'h2 : count; // @[src/main/scala/rocket/PTW.scala 659:27 660:15 259:18]
  wire [2:0] _GEN_137 = 3'h7 == state ? 3'h0 : state; // @[src/main/scala/rocket/PTW.scala 594:18 657:18 590:31]
  wire  _GEN_138 = 3'h7 == state & _GEN_27; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire  _GEN_139 = 3'h7 == state & r_req_dest; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire [1:0] _GEN_140 = 3'h7 == state ? _GEN_134 : count; // @[src/main/scala/rocket/PTW.scala 259:18 594:18]
  wire [2:0] _GEN_142 = 3'h4 == state ? _GEN_129 : _GEN_137; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  _GEN_143 = 3'h4 == state & _traverse_T_16; // @[src/main/scala/rocket/PTW.scala 594:18 405:26 649:30]
  wire  _GEN_144 = 3'h4 == state ? _GEN_128 : resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 594:18 260:24]
  wire  _GEN_145 = 3'h4 == state ? _GEN_130 : _GEN_138; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  _GEN_146 = 3'h4 == state ? _GEN_131 : _GEN_139; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire [1:0] _GEN_147 = 3'h4 == state ? count : _GEN_140; // @[src/main/scala/rocket/PTW.scala 259:18 594:18]
  wire [2:0] _GEN_149 = 3'h2 == state ? 3'h4 : _GEN_142; // @[src/main/scala/rocket/PTW.scala 594:18 645:18]
  wire  _GEN_150 = 3'h2 == state ? 1'h0 : _GEN_143; // @[src/main/scala/rocket/PTW.scala 594:18 405:26]
  wire  _GEN_151 = 3'h2 == state ? resp_ae_ptw : _GEN_144; // @[src/main/scala/rocket/PTW.scala 594:18 260:24]
  wire  _GEN_152 = 3'h2 == state ? 1'h0 : _GEN_145; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire  _GEN_153 = 3'h2 == state ? 1'h0 : _GEN_146; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire [2:0] _GEN_162 = 3'h1 == state ? _GEN_119 : _GEN_149; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  _GEN_163 = 3'h1 == state ? 1'h0 : _GEN_150; // @[src/main/scala/rocket/PTW.scala 594:18 405:26]
  wire  _GEN_164 = 3'h1 == state ? resp_ae_ptw : _GEN_151; // @[src/main/scala/rocket/PTW.scala 594:18 260:24]
  wire  _GEN_165 = 3'h1 == state ? 1'h0 : _GEN_152; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire  _GEN_166 = 3'h1 == state ? 1'h0 : _GEN_153; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire [2:0] _GEN_173 = 3'h0 == state ? _GEN_98 : _GEN_162; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  _GEN_180 = 3'h0 == state ? _GEN_105 : _GEN_164; // @[src/main/scala/rocket/PTW.scala 594:18]
  wire  _GEN_181 = 3'h0 == state ? _GEN_106 : resp_ae_final; // @[src/main/scala/rocket/PTW.scala 594:18 261:26]
  wire  _GEN_182 = 3'h0 == state ? _GEN_107 : resp_pf; // @[src/main/scala/rocket/PTW.scala 594:18 262:20]
  wire  _GEN_194 = 3'h0 == state ? 1'h0 : _GEN_165; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire  _GEN_195 = 3'h0 == state ? 1'h0 : _GEN_166; // @[src/main/scala/rocket/PTW.scala 594:18 242:27]
  wire [43:0] _r_pte_T_17 = {r_pte_ppn[43:18],r_req_addr[17:0]}; // @[src/main/scala/rocket/PTW.scala 355:44]
  wire [43:0] _r_pte_T_20 = {r_pte_ppn[43:9],r_req_addr[8:0]}; // @[src/main/scala/rocket/PTW.scala 355:44]
  wire  r_pte_truncIdx = count[0]; // @[src/main/scala/util/package.scala 32:47]
  wire [43:0] r_pte_pte_3_ppn = r_pte_truncIdx ? _r_pte_T_20 : _r_pte_T_17; // @[src/main/scala/util/package.scala 33:76]
  wire [43:0] _r_pte_T_25_ppn = _T_77 ? io_dpath_ptbr_ppn : r_pte_ppn; // @[src/main/scala/rocket/PTW.scala 691:8]
  wire [43:0] _r_pte_T_26_ppn = state == 3'h7 & _T_93 & count != 2'h2 ? r_pte_pte_3_ppn : _r_pte_T_25_ppn; // @[src/main/scala/rocket/PTW.scala 689:8]
  wire [43:0] _r_pte_T_27_ppn = mem_resp_valid ? pte_ppn : _r_pte_T_26_ppn; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_d = mem_resp_valid ? tmp_d : r_pte_d; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_a = mem_resp_valid ? tmp_a : r_pte_a; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_g = mem_resp_valid ? tmp_g : r_pte_g; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_u = mem_resp_valid ? tmp_u : r_pte_u; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_x = mem_resp_valid ? tmp_x : r_pte_x; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_w = mem_resp_valid ? tmp_w : r_pte_w; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_r = mem_resp_valid ? tmp_r : r_pte_r; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  _r_pte_T_27_v = mem_resp_valid ? pte_v : r_pte_v; // @[src/main/scala/rocket/PTW.scala 687:8]
  wire  ae = pte_v & invalid_paddr; // @[src/main/scala/rocket/PTW.scala 708:22]
  wire  pf = pte_v & tmp_reserved_for_future != 10'h0; // @[src/main/scala/rocket/PTW.scala 709:22]
  wire  success = pte_v & ~ae & ~pf; // @[src/main/scala/rocket/PTW.scala 710:34]
  wire [43:0] r_pte_pte_1_ppn = {{24'd0}, pte_cache_data}; // @[src/main/scala/rocket/PTW.scala 780:26 781:13]
  wire  line_1021_clock;
  wire  line_1021_reset;
  wire  line_1021_valid;
  reg  line_1021_valid_reg;
  wire  _T_101 = ~(_T_23 | state == 3'h2); // @[src/main/scala/rocket/PTW.scala 695:11]
  wire  line_1022_clock;
  wire  line_1022_reset;
  wire  line_1022_valid;
  reg  line_1022_valid_reg;
  wire  line_1023_clock;
  wire  line_1023_reset;
  wire  line_1023_valid;
  reg  line_1023_valid_reg;
  wire  _GEN_196 = _GEN_27 | _GEN_194; // @[src/main/scala/rocket/PTW.scala 697:{28,28}]
  wire  line_1024_clock;
  wire  line_1024_reset;
  wire  line_1024_valid;
  reg  line_1024_valid_reg;
  wire  _GEN_197 = r_req_dest | _GEN_195; // @[src/main/scala/rocket/PTW.scala 697:{28,28}]
  wire  line_1025_clock;
  wire  line_1025_reset;
  wire  line_1025_valid;
  reg  line_1025_valid_reg;
  wire  line_1026_clock;
  wire  line_1026_reset;
  wire  line_1026_valid;
  reg  line_1026_valid_reg;
  wire  _T_107 = ~(state == 3'h5); // @[src/main/scala/rocket/PTW.scala 701:11]
  wire  line_1027_clock;
  wire  line_1027_reset;
  wire  line_1027_valid;
  reg  line_1027_valid_reg;
  wire  line_1028_clock;
  wire  line_1028_reset;
  wire  line_1028_valid;
  reg  line_1028_valid_reg;
  wire  line_1029_clock;
  wire  line_1029_reset;
  wire  line_1029_valid;
  reg  line_1029_valid_reg;
  wire  _l2_refill_T_3 = success & _pte_addr_vpn_idx_T_2 & ~r_req_need_gpa; // @[src/main/scala/rocket/PTW.scala 722:58]
  wire  line_1030_clock;
  wire  line_1030_reset;
  wire  line_1030_valid;
  reg  line_1030_valid_reg;
  wire  line_1031_clock;
  wire  line_1031_reset;
  wire  line_1031_valid;
  reg  line_1031_valid_reg;
  wire  _resp_ae_ptw_T_16 = ae & _traverse_T_16 & _traverse_T_13; // @[src/main/scala/rocket/PTW.scala 734:53]
  wire  _GEN_231 = traverse ? 1'h0 : _l2_refill_T_3; // @[src/main/scala/rocket/PTW.scala 703:21 410:26]
  wire [2:0] _GEN_232 = traverse ? 3'h1 : 3'h0; // @[src/main/scala/rocket/PTW.scala 702:16 703:21]
  wire [2:0] _GEN_242 = mem_resp_valid ? _GEN_232 : _GEN_173; // @[src/main/scala/rocket/PTW.scala 700:25]
  wire  line_1032_clock;
  wire  line_1032_reset;
  wire  line_1032_valid;
  reg  line_1032_valid_reg;
  wire  line_1033_clock;
  wire  line_1033_reset;
  wire  line_1033_valid;
  reg  line_1033_valid_reg;
  wire  _T_125 = ~(state == 3'h4); // @[src/main/scala/rocket/PTW.scala 745:11]
  wire  line_1034_clock;
  wire  line_1034_reset;
  wire  line_1034_valid;
  reg  line_1034_valid_reg;
  Arbiter arb ( // @[src/main/scala/rocket/PTW.scala 236:19]
    .clock(arb_clock),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_bits_addr(arb_io_in_0_bits_bits_addr),
    .io_in_0_bits_bits_need_gpa(arb_io_in_0_bits_bits_need_gpa),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_valid(arb_io_in_1_bits_valid),
    .io_in_1_bits_bits_addr(arb_io_in_1_bits_bits_addr),
    .io_in_1_bits_bits_need_gpa(arb_io_in_1_bits_bits_need_gpa),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_valid(arb_io_out_bits_valid),
    .io_out_bits_bits_addr(arb_io_out_bits_bits_addr),
    .io_out_bits_bits_need_gpa(arb_io_out_bits_bits_need_gpa),
    .io_chosen(arb_io_chosen)
  );
  OptimizationBarrier_18 state_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(state_barrier_clock),
    .reset(state_barrier_reset),
    .io_x(state_barrier_io_x),
    .io_y(state_barrier_io_y)
  );
  OptimizationBarrier_19 r_pte_barrier ( // @[src/main/scala/util/package.scala 259:25]
    .clock(r_pte_barrier_clock),
    .reset(r_pte_barrier_reset),
    .io_x_ppn(r_pte_barrier_io_x_ppn),
    .io_x_d(r_pte_barrier_io_x_d),
    .io_x_a(r_pte_barrier_io_x_a),
    .io_x_g(r_pte_barrier_io_x_g),
    .io_x_u(r_pte_barrier_io_x_u),
    .io_x_x(r_pte_barrier_io_x_x),
    .io_x_w(r_pte_barrier_io_x_w),
    .io_x_r(r_pte_barrier_io_x_r),
    .io_x_v(r_pte_barrier_io_x_v),
    .io_y_ppn(r_pte_barrier_io_y_ppn),
    .io_y_d(r_pte_barrier_io_y_d),
    .io_y_a(r_pte_barrier_io_y_a),
    .io_y_g(r_pte_barrier_io_y_g),
    .io_y_u(r_pte_barrier_io_y_u),
    .io_y_x(r_pte_barrier_io_y_x),
    .io_y_w(r_pte_barrier_io_y_w),
    .io_y_r(r_pte_barrier_io_y_r),
    .io_y_v(r_pte_barrier_io_y_v)
  );
  GEN_w1_line #(.COVER_INDEX(988)) line_988 (
    .clock(line_988_clock),
    .reset(line_988_reset),
    .valid(line_988_valid)
  );
  GEN_w1_line #(.COVER_INDEX(989)) line_989 (
    .clock(line_989_clock),
    .reset(line_989_reset),
    .valid(line_989_valid)
  );
  GEN_w1_line #(.COVER_INDEX(990)) line_990 (
    .clock(line_990_clock),
    .reset(line_990_reset),
    .valid(line_990_valid)
  );
  GEN_w1_line #(.COVER_INDEX(991)) line_991 (
    .clock(line_991_clock),
    .reset(line_991_reset),
    .valid(line_991_valid)
  );
  GEN_w1_line #(.COVER_INDEX(992)) line_992 (
    .clock(line_992_clock),
    .reset(line_992_reset),
    .valid(line_992_valid)
  );
  GEN_w1_line #(.COVER_INDEX(993)) line_993 (
    .clock(line_993_clock),
    .reset(line_993_reset),
    .valid(line_993_valid)
  );
  GEN_w1_line #(.COVER_INDEX(994)) line_994 (
    .clock(line_994_clock),
    .reset(line_994_reset),
    .valid(line_994_valid)
  );
  GEN_w1_line #(.COVER_INDEX(995)) line_995 (
    .clock(line_995_clock),
    .reset(line_995_reset),
    .valid(line_995_valid)
  );
  GEN_w1_line #(.COVER_INDEX(996)) line_996 (
    .clock(line_996_clock),
    .reset(line_996_reset),
    .valid(line_996_valid)
  );
  GEN_w1_line #(.COVER_INDEX(997)) line_997 (
    .clock(line_997_clock),
    .reset(line_997_reset),
    .valid(line_997_valid)
  );
  GEN_w1_line #(.COVER_INDEX(998)) line_998 (
    .clock(line_998_clock),
    .reset(line_998_reset),
    .valid(line_998_valid)
  );
  GEN_w1_line #(.COVER_INDEX(999)) line_999 (
    .clock(line_999_clock),
    .reset(line_999_reset),
    .valid(line_999_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1000)) line_1000 (
    .clock(line_1000_clock),
    .reset(line_1000_reset),
    .valid(line_1000_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1001)) line_1001 (
    .clock(line_1001_clock),
    .reset(line_1001_reset),
    .valid(line_1001_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1002)) line_1002 (
    .clock(line_1002_clock),
    .reset(line_1002_reset),
    .valid(line_1002_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1003)) line_1003 (
    .clock(line_1003_clock),
    .reset(line_1003_reset),
    .valid(line_1003_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1004)) line_1004 (
    .clock(line_1004_clock),
    .reset(line_1004_reset),
    .valid(line_1004_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1005)) line_1005 (
    .clock(line_1005_clock),
    .reset(line_1005_reset),
    .valid(line_1005_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1006)) line_1006 (
    .clock(line_1006_clock),
    .reset(line_1006_reset),
    .valid(line_1006_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1007)) line_1007 (
    .clock(line_1007_clock),
    .reset(line_1007_reset),
    .valid(line_1007_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1008)) line_1008 (
    .clock(line_1008_clock),
    .reset(line_1008_reset),
    .valid(line_1008_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1009)) line_1009 (
    .clock(line_1009_clock),
    .reset(line_1009_reset),
    .valid(line_1009_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1010)) line_1010 (
    .clock(line_1010_clock),
    .reset(line_1010_reset),
    .valid(line_1010_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1011)) line_1011 (
    .clock(line_1011_clock),
    .reset(line_1011_reset),
    .valid(line_1011_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1012)) line_1012 (
    .clock(line_1012_clock),
    .reset(line_1012_reset),
    .valid(line_1012_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1013)) line_1013 (
    .clock(line_1013_clock),
    .reset(line_1013_reset),
    .valid(line_1013_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1014)) line_1014 (
    .clock(line_1014_clock),
    .reset(line_1014_reset),
    .valid(line_1014_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1015)) line_1015 (
    .clock(line_1015_clock),
    .reset(line_1015_reset),
    .valid(line_1015_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1016)) line_1016 (
    .clock(line_1016_clock),
    .reset(line_1016_reset),
    .valid(line_1016_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1017)) line_1017 (
    .clock(line_1017_clock),
    .reset(line_1017_reset),
    .valid(line_1017_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1018)) line_1018 (
    .clock(line_1018_clock),
    .reset(line_1018_reset),
    .valid(line_1018_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1019)) line_1019 (
    .clock(line_1019_clock),
    .reset(line_1019_reset),
    .valid(line_1019_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1020)) line_1020 (
    .clock(line_1020_clock),
    .reset(line_1020_reset),
    .valid(line_1020_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1021)) line_1021 (
    .clock(line_1021_clock),
    .reset(line_1021_reset),
    .valid(line_1021_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1022)) line_1022 (
    .clock(line_1022_clock),
    .reset(line_1022_reset),
    .valid(line_1022_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1023)) line_1023 (
    .clock(line_1023_clock),
    .reset(line_1023_reset),
    .valid(line_1023_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1024)) line_1024 (
    .clock(line_1024_clock),
    .reset(line_1024_reset),
    .valid(line_1024_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1025)) line_1025 (
    .clock(line_1025_clock),
    .reset(line_1025_reset),
    .valid(line_1025_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1026)) line_1026 (
    .clock(line_1026_clock),
    .reset(line_1026_reset),
    .valid(line_1026_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1027)) line_1027 (
    .clock(line_1027_clock),
    .reset(line_1027_reset),
    .valid(line_1027_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1028)) line_1028 (
    .clock(line_1028_clock),
    .reset(line_1028_reset),
    .valid(line_1028_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1029)) line_1029 (
    .clock(line_1029_clock),
    .reset(line_1029_reset),
    .valid(line_1029_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1030)) line_1030 (
    .clock(line_1030_clock),
    .reset(line_1030_reset),
    .valid(line_1030_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1031)) line_1031 (
    .clock(line_1031_clock),
    .reset(line_1031_reset),
    .valid(line_1031_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1032)) line_1032 (
    .clock(line_1032_clock),
    .reset(line_1032_reset),
    .valid(line_1032_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1033)) line_1033 (
    .clock(line_1033_clock),
    .reset(line_1033_reset),
    .valid(line_1033_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1034)) line_1034 (
    .clock(line_1034_clock),
    .reset(line_1034_reset),
    .valid(line_1034_valid)
  );
  assign line_988_clock = clock;
  assign line_988_reset = reset;
  assign line_988_valid = _T_1 ^ line_988_valid_reg;
  assign line_989_clock = clock;
  assign line_989_reset = reset;
  assign line_989_valid = _T_5 ^ line_989_valid_reg;
  assign line_990_clock = clock;
  assign line_990_reset = reset;
  assign line_990_valid = _T_9 ^ line_990_valid_reg;
  assign line_991_clock = clock;
  assign line_991_reset = reset;
  assign line_991_valid = _T_22 ^ line_991_valid_reg;
  assign line_992_clock = clock;
  assign line_992_reset = reset;
  assign line_992_valid = ~r ^ line_992_valid_reg;
  assign line_993_clock = clock;
  assign line_993_reset = reset;
  assign line_993_valid = r ^ line_993_valid_reg;
  assign line_994_clock = clock;
  assign line_994_reset = reset;
  assign line_994_valid = ~r ^ line_994_valid_reg;
  assign line_995_clock = clock;
  assign line_995_reset = reset;
  assign line_995_valid = r ^ line_995_valid_reg;
  assign line_996_clock = clock;
  assign line_996_reset = reset;
  assign line_996_valid = _T_24 ^ line_996_valid_reg;
  assign line_997_clock = clock;
  assign line_997_reset = reset;
  assign line_997_valid = _T_29 ^ line_997_valid_reg;
  assign line_998_clock = clock;
  assign line_998_reset = reset;
  assign line_998_valid = _T_29 ^ line_998_valid_reg;
  assign line_999_clock = clock;
  assign line_999_reset = reset;
  assign line_999_valid = _T_74 ^ line_999_valid_reg;
  assign line_1000_clock = clock;
  assign line_1000_reset = reset;
  assign line_1000_valid = _T_75 ^ line_1000_valid_reg;
  assign line_1001_clock = clock;
  assign line_1001_reset = reset;
  assign line_1001_valid = _T_76 ^ line_1001_valid_reg;
  assign line_1002_clock = clock;
  assign line_1002_reset = reset;
  assign line_1002_valid = _T_77 ^ line_1002_valid_reg;
  assign line_1003_clock = clock;
  assign line_1003_reset = reset;
  assign line_1003_valid = _T_74 ^ line_1003_valid_reg;
  assign line_1004_clock = clock;
  assign line_1004_reset = reset;
  assign line_1004_valid = _T_82 ^ line_1004_valid_reg;
  assign line_1005_clock = clock;
  assign line_1005_reset = reset;
  assign line_1005_valid = _T_76 ^ line_1005_valid_reg;
  assign line_1006_clock = clock;
  assign line_1006_reset = reset;
  assign line_1006_valid = _T_83 ^ line_1006_valid_reg;
  assign line_1007_clock = clock;
  assign line_1007_reset = reset;
  assign line_1007_valid = pte_cache_hit ^ line_1007_valid_reg;
  assign line_1008_clock = clock;
  assign line_1008_reset = reset;
  assign line_1008_valid = pte_cache_hit ^ line_1008_valid_reg;
  assign line_1009_clock = clock;
  assign line_1009_reset = reset;
  assign line_1009_valid = _T_83 ^ line_1009_valid_reg;
  assign line_1010_clock = clock;
  assign line_1010_reset = reset;
  assign line_1010_valid = _T_86 ^ line_1010_valid_reg;
  assign line_1011_clock = clock;
  assign line_1011_reset = reset;
  assign line_1011_valid = _T_86 ^ line_1011_valid_reg;
  assign line_1012_clock = clock;
  assign line_1012_reset = reset;
  assign line_1012_valid = _T_87 ^ line_1012_valid_reg;
  assign line_1013_clock = clock;
  assign line_1013_reset = reset;
  assign line_1013_valid = io_mem_s2_xcpt_ae_ld ^ line_1013_valid_reg;
  assign line_1014_clock = clock;
  assign line_1014_reset = reset;
  assign line_1014_valid = ~r_req_dest ^ line_1014_valid_reg;
  assign line_1015_clock = clock;
  assign line_1015_reset = reset;
  assign line_1015_valid = r_req_dest ^ line_1015_valid_reg;
  assign line_1016_clock = clock;
  assign line_1016_reset = reset;
  assign line_1016_valid = _T_87 ^ line_1016_valid_reg;
  assign line_1017_clock = clock;
  assign line_1017_reset = reset;
  assign line_1017_valid = _T_90 ^ line_1017_valid_reg;
  assign line_1018_clock = clock;
  assign line_1018_reset = reset;
  assign line_1018_valid = ~r_req_dest ^ line_1018_valid_reg;
  assign line_1019_clock = clock;
  assign line_1019_reset = reset;
  assign line_1019_valid = r_req_dest ^ line_1019_valid_reg;
  assign line_1020_clock = clock;
  assign line_1020_reset = reset;
  assign line_1020_valid = _T_93 ^ line_1020_valid_reg;
  assign line_1021_clock = clock;
  assign line_1021_reset = reset;
  assign line_1021_valid = _T_74 ^ line_1021_valid_reg;
  assign line_1022_clock = clock;
  assign line_1022_reset = reset;
  assign line_1022_valid = _T_101 ^ line_1022_valid_reg;
  assign line_1023_clock = clock;
  assign line_1023_reset = reset;
  assign line_1023_valid = ~r_req_dest ^ line_1023_valid_reg;
  assign line_1024_clock = clock;
  assign line_1024_reset = reset;
  assign line_1024_valid = r_req_dest ^ line_1024_valid_reg;
  assign line_1025_clock = clock;
  assign line_1025_reset = reset;
  assign line_1025_valid = mem_resp_valid ^ line_1025_valid_reg;
  assign line_1026_clock = clock;
  assign line_1026_reset = reset;
  assign line_1026_valid = _T_74 ^ line_1026_valid_reg;
  assign line_1027_clock = clock;
  assign line_1027_reset = reset;
  assign line_1027_valid = _T_107 ^ line_1027_valid_reg;
  assign line_1028_clock = clock;
  assign line_1028_reset = reset;
  assign line_1028_valid = traverse ^ line_1028_valid_reg;
  assign line_1029_clock = clock;
  assign line_1029_reset = reset;
  assign line_1029_valid = traverse ^ line_1029_valid_reg;
  assign line_1030_clock = clock;
  assign line_1030_reset = reset;
  assign line_1030_valid = ~r_req_dest ^ line_1030_valid_reg;
  assign line_1031_clock = clock;
  assign line_1031_reset = reset;
  assign line_1031_valid = r_req_dest ^ line_1031_valid_reg;
  assign line_1032_clock = clock;
  assign line_1032_reset = reset;
  assign line_1032_valid = io_mem_s2_nack ^ line_1032_valid_reg;
  assign line_1033_clock = clock;
  assign line_1033_reset = reset;
  assign line_1033_valid = _T_74 ^ line_1033_valid_reg;
  assign line_1034_clock = clock;
  assign line_1034_reset = reset;
  assign line_1034_valid = _T_125 ^ line_1034_valid_reg;
  assign io_requestor_0_req_ready = arb_io_in_0_ready; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign io_requestor_0_resp_valid = resp_valid_0; // @[src/main/scala/rocket/PTW.scala 563:32]
  assign io_requestor_0_resp_bits_ae_ptw = resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 564:38]
  assign io_requestor_0_resp_bits_ae_final = resp_ae_final; // @[src/main/scala/rocket/PTW.scala 565:40]
  assign io_requestor_0_resp_bits_pf = resp_pf; // @[src/main/scala/rocket/PTW.scala 566:34]
  assign io_requestor_0_resp_bits_pte_ppn = r_pte_ppn; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_d = r_pte_d; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_a = r_pte_a; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_g = r_pte_g; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_u = r_pte_u; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_x = r_pte_x; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_w = r_pte_w; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_r = r_pte_r; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_pte_v = r_pte_v; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_0_resp_bits_level = count; // @[src/main/scala/rocket/PTW.scala 290:25]
  assign io_requestor_0_resp_bits_homogeneous = count == 2'h3 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_3; // @[src/main/scala/util/package.scala 33:76]
  assign io_requestor_0_ptbr_mode = io_dpath_ptbr_mode; // @[src/main/scala/rocket/PTW.scala 579:26]
  assign io_requestor_0_status_mxr = io_dpath_status_mxr; // @[src/main/scala/rocket/PTW.scala 583:28]
  assign io_requestor_0_status_sum = io_dpath_status_sum; // @[src/main/scala/rocket/PTW.scala 583:28]
  assign io_requestor_1_req_ready = arb_io_in_1_ready; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign io_requestor_1_resp_valid = resp_valid_1; // @[src/main/scala/rocket/PTW.scala 563:32]
  assign io_requestor_1_resp_bits_ae_ptw = resp_ae_ptw; // @[src/main/scala/rocket/PTW.scala 564:38]
  assign io_requestor_1_resp_bits_ae_final = resp_ae_final; // @[src/main/scala/rocket/PTW.scala 565:40]
  assign io_requestor_1_resp_bits_pf = resp_pf; // @[src/main/scala/rocket/PTW.scala 566:34]
  assign io_requestor_1_resp_bits_pte_ppn = r_pte_ppn; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_d = r_pte_d; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_a = r_pte_a; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_g = r_pte_g; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_u = r_pte_u; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_x = r_pte_x; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_w = r_pte_w; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_r = r_pte_r; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_pte_v = r_pte_v; // @[src/main/scala/rocket/PTW.scala 571:35]
  assign io_requestor_1_resp_bits_level = count; // @[src/main/scala/rocket/PTW.scala 290:25]
  assign io_requestor_1_resp_bits_homogeneous = count == 2'h3 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_3; // @[src/main/scala/util/package.scala 33:76]
  assign io_requestor_1_ptbr_mode = io_dpath_ptbr_mode; // @[src/main/scala/rocket/PTW.scala 579:26]
  assign io_requestor_1_status_prv = io_dpath_status_prv; // @[src/main/scala/rocket/PTW.scala 583:28]
  assign io_mem_req_valid = _T_23 | state == 3'h3; // @[src/main/scala/rocket/PTW.scala 527:39]
  assign io_mem_req_bits_addr = {{8'd0}, pte_addr}; // @[src/main/scala/rocket/PTW.scala 532:24]
  assign io_mem_s1_kill = state != 3'h2; // @[src/main/scala/rocket/PTW.scala 542:37]
  assign io_dpath_perf_l2hit = 1'h0; // @[src/main/scala/rocket/PTW.scala 413:23]
  assign io_dpath_perf_pte_miss = 3'h0 == state ? 1'h0 : _GEN_163; // @[src/main/scala/rocket/PTW.scala 594:18 405:26]
  assign io_dpath_perf_pte_hit = pte_hit & _T_23 & ~io_dpath_perf_l2hit; // @[src/main/scala/rocket/PTW.scala 406:57]
  assign arb_clock = clock;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_requestor_0_req_valid; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_0_bits_bits_addr = io_requestor_0_req_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_0_bits_bits_need_gpa = io_requestor_0_req_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_1_valid = io_requestor_1_req_valid; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_1_bits_valid = io_requestor_1_req_bits_valid; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_1_bits_bits_addr = io_requestor_1_req_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_in_1_bits_bits_need_gpa = io_requestor_1_req_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 238:13]
  assign arb_io_out_ready = state == 3'h0 & ~l2_refill; // @[src/main/scala/rocket/PTW.scala 240:43]
  assign state_barrier_clock = clock;
  assign state_barrier_reset = reset;
  assign state_barrier_io_x = io_mem_s2_nack ? 3'h1 : _GEN_242; // @[src/main/scala/rocket/PTW.scala 744:25 746:16]
  assign r_pte_barrier_clock = clock;
  assign r_pte_barrier_reset = reset;
  assign r_pte_barrier_io_x_ppn = _T_23 & pte_cache_hit ? r_pte_pte_1_ppn : _r_pte_T_27_ppn; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_d = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_d; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_a = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_a; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_g = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_g; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_u = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_u; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_x = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_x; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_w = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_w; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_r = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_r; // @[src/main/scala/rocket/PTW.scala 683:8]
  assign r_pte_barrier_io_x_v = _T_23 & pte_cache_hit ? 1'h0 : _r_pte_T_27_v; // @[src/main/scala/rocket/PTW.scala 683:8]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rocket/PTW.scala 233:22]
      state <= 3'h0; // @[src/main/scala/rocket/PTW.scala 233:22]
    end else begin
      state <= state_barrier_io_y; // @[src/main/scala/rocket/PTW.scala 591:9]
    end
    l2_refill <= mem_resp_valid & _GEN_231; // @[src/main/scala/rocket/PTW.scala 700:25 410:26]
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        resp_valid_0 <= _GEN_194;
      end else begin
        resp_valid_0 <= _GEN_196;
      end
    end else begin
      resp_valid_0 <= _GEN_194;
    end
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        resp_valid_1 <= _GEN_195;
      end else begin
        resp_valid_1 <= _GEN_197;
      end
    end else begin
      resp_valid_1 <= _GEN_195;
    end
    invalidated <= io_dpath_sfence_valid | invalidated & _clock_en_T; // @[src/main/scala/rocket/PTW.scala 523:40]
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        count <= _count_T_2; // @[src/main/scala/rocket/PTW.scala 705:13]
      end
    end else if (3'h0 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      if (_T_77) begin // @[src/main/scala/rocket/PTW.scala 596:30]
        count <= 2'h0; // @[src/main/scala/rocket/PTW.scala 607:21]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      if (pte_cache_hit) begin // @[src/main/scala/rocket/PTW.scala 636:34]
        count <= _count_T_2; // @[src/main/scala/rocket/PTW.scala 637:15]
      end
    end else if (!(3'h2 == state)) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      count <= _GEN_147;
    end
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        resp_ae_ptw <= _GEN_180;
      end else begin
        resp_ae_ptw <= _resp_ae_ptw_T_16;
      end
    end else begin
      resp_ae_ptw <= _GEN_180;
    end
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        resp_ae_final <= _GEN_181;
      end else begin
        resp_ae_final <= ae;
      end
    end else begin
      resp_ae_final <= _GEN_181;
    end
    if (mem_resp_valid) begin // @[src/main/scala/rocket/PTW.scala 700:25]
      if (traverse) begin // @[src/main/scala/rocket/PTW.scala 703:21]
        resp_pf <= _GEN_182;
      end else begin
        resp_pf <= pf;
      end
    end else begin
      resp_pf <= _GEN_182;
    end
    if (3'h0 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      if (_T_77) begin // @[src/main/scala/rocket/PTW.scala 596:30]
        r_req_addr <= arb_io_out_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 602:15]
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      if (_T_77) begin // @[src/main/scala/rocket/PTW.scala 596:30]
        r_req_need_gpa <= arb_io_out_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 602:15]
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      if (_T_77) begin // @[src/main/scala/rocket/PTW.scala 596:30]
        r_req_dest <= arb_io_chosen; // @[src/main/scala/rocket/PTW.scala 603:20]
      end
    end
    r_pte_ppn <= r_pte_barrier_io_y_ppn; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_d <= r_pte_barrier_io_y_d; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_a <= r_pte_barrier_io_y_a; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_g <= r_pte_barrier_io_y_g; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_u <= r_pte_barrier_io_y_u; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_x <= r_pte_barrier_io_y_x; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_w <= r_pte_barrier_io_y_w; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_r <= r_pte_barrier_io_y_r; // @[src/main/scala/rocket/PTW.scala 677:9]
    r_pte_v <= r_pte_barrier_io_y_v; // @[src/main/scala/rocket/PTW.scala 677:9]
    mem_resp_valid <= io_mem_resp_valid; // @[src/main/scala/rocket/PTW.scala 293:31]
    mem_resp_data <= io_mem_resp_bits_data; // @[src/main/scala/rocket/PTW.scala 294:30]
    line_988_valid_reg <= _T_1;
    line_989_valid_reg <= _T_5;
    line_990_valid_reg <= _T_9;
    if (reset) begin // @[src/main/scala/util/Replacement.scala 168:72]
      state_reg <= 1'h0; // @[src/main/scala/util/Replacement.scala 168:72]
    end else if (pte_cache_hit & state == 3'h1) begin // @[src/main/scala/rocket/PTW.scala 389:35]
      state_reg <= _state_reg_T_3; // @[src/main/scala/util/Replacement.scala 172:15]
    end else if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      state_reg <= _GEN_3; // @[src/main/scala/util/Replacement.scala 172:15]
    end
    if (reset) begin // @[src/main/scala/rocket/PTW.scala 364:24]
      valid <= 2'h0; // @[src/main/scala/rocket/PTW.scala 364:24]
    end else if (io_dpath_sfence_valid & ~io_dpath_sfence_bits_rs1) begin // @[src/main/scala/rocket/PTW.scala 390:113]
      valid <= 2'h0; // @[src/main/scala/rocket/PTW.scala 390:121]
    end else if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      valid <= _valid_T_1; // @[src/main/scala/rocket/PTW.scala 383:13]
    end
    if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      if (~r) begin // @[src/main/scala/rocket/PTW.scala 384:15]
        tags__0 <= tag[31:0]; // @[src/main/scala/rocket/PTW.scala 384:15]
      end
    end
    if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      if (r) begin // @[src/main/scala/rocket/PTW.scala 384:15]
        tags__1 <= tag[31:0]; // @[src/main/scala/rocket/PTW.scala 384:15]
      end
    end
    if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      if (~r) begin // @[src/main/scala/rocket/PTW.scala 385:15]
        data__0 <= pte_ppn[19:0]; // @[src/main/scala/rocket/PTW.scala 385:15]
      end
    end
    if (mem_resp_valid & traverse & _traverse_T_16 & ~_hit_T & ~invalidated) begin // @[src/main/scala/rocket/PTW.scala 381:82]
      if (r) begin // @[src/main/scala/rocket/PTW.scala 385:15]
        data__1 <= pte_ppn[19:0]; // @[src/main/scala/rocket/PTW.scala 385:15]
      end
    end
    line_991_valid_reg <= _T_22;
    line_992_valid_reg <= ~r;
    if (&valid) begin // @[src/main/scala/rocket/PTW.scala 382:18]
      line_993_valid_reg <= state_reg;
    end else if (_r_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
      line_993_valid_reg <= 1'h0;
    end else begin
      line_993_valid_reg <= 1'h1;
    end
    line_994_valid_reg <= ~r;
    if (&valid) begin // @[src/main/scala/rocket/PTW.scala 382:18]
      line_995_valid_reg <= state_reg;
    end else if (_r_T_2[0]) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
      line_995_valid_reg <= 1'h0;
    end else begin
      line_995_valid_reg <= 1'h1;
    end
    line_996_valid_reg <= _T_24;
    line_997_valid_reg <= _T_29;
    line_998_valid_reg <= _T_29;
    if (3'h0 == state) begin // @[src/main/scala/rocket/PTW.scala 594:18]
      pte_hit <= 1'h0; // @[src/main/scala/rocket/PTW.scala 404:24]
    end else begin
      pte_hit <= 3'h1 == state & pte_cache_hit;
    end
    line_999_valid_reg <= _T_74;
    line_1000_valid_reg <= _T_75;
    line_1001_valid_reg <= _T_76;
    line_1002_valid_reg <= _T_77;
    line_1003_valid_reg <= _T_74;
    line_1004_valid_reg <= _T_82;
    line_1005_valid_reg <= _T_76;
    line_1006_valid_reg <= _T_83;
    line_1007_valid_reg <= pte_cache_hit;
    line_1008_valid_reg <= pte_cache_hit;
    line_1009_valid_reg <= _T_83;
    line_1010_valid_reg <= _T_86;
    line_1011_valid_reg <= _T_86;
    line_1012_valid_reg <= _T_87;
    line_1013_valid_reg <= io_mem_s2_xcpt_ae_ld;
    line_1014_valid_reg <= ~r_req_dest;
    line_1015_valid_reg <= r_req_dest;
    line_1016_valid_reg <= _T_87;
    line_1017_valid_reg <= _T_90;
    line_1018_valid_reg <= ~r_req_dest;
    line_1019_valid_reg <= r_req_dest;
    line_1020_valid_reg <= _T_93;
    line_1021_valid_reg <= _T_74;
    line_1022_valid_reg <= _T_101;
    line_1023_valid_reg <= ~r_req_dest;
    line_1024_valid_reg <= r_req_dest;
    line_1025_valid_reg <= mem_resp_valid;
    line_1026_valid_reg <= _T_74;
    line_1027_valid_reg <= _T_107;
    line_1028_valid_reg <= traverse;
    line_1029_valid_reg <= traverse;
    line_1030_valid_reg <= ~r_req_dest;
    line_1031_valid_reg <= r_req_dest;
    line_1032_valid_reg <= io_mem_s2_nack;
    line_1033_valid_reg <= _T_74;
    line_1034_valid_reg <= _T_125;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(io_dpath_perf_l2hit & (io_dpath_perf_pte_miss | io_dpath_perf_pte_hit)))) begin
          $fwrite(32'h80000002,
            "Assertion failed: PTE Cache Hit/Miss Performance Monitor Events are lower priority than L2TLB Hit event\n    at PTW.scala:407 assert(!(io.dpath.perf.l2hit && (io.dpath.perf.pte_miss || io.dpath.perf.pte_hit)),\n"
            ); // @[src/main/scala/rocket/PTW.scala 407:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_76 & _T_77 & _T_74 & ~(~arb_io_out_bits_bits_need_gpa)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at PTW.scala:622 assert(!arb.io.out.bits.bits.need_gpa || arb.io.out.bits.bits.stage2)\n"
            ); // @[src/main/scala/rocket/PTW.scala 622:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (mem_resp_valid & _T_74 & ~(state == 3'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:701 assert(state === s_wait3)\n"); // @[src/main/scala/rocket/PTW.scala 701:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_s2_nack & _T_74 & ~(state == 3'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:745 assert(state === s_wait2)\n"); // @[src/main/scala/rocket/PTW.scala 745:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  l2_refill = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  resp_valid_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  resp_valid_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  invalidated = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  count = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  resp_ae_ptw = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  resp_ae_final = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  resp_pf = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_req_addr = _RAND_9[26:0];
  _RAND_10 = {1{`RANDOM}};
  r_req_need_gpa = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_req_dest = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  r_pte_ppn = _RAND_12[43:0];
  _RAND_13 = {1{`RANDOM}};
  r_pte_d = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_pte_a = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_pte_g = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_pte_u = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_pte_x = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_pte_w = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_pte_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_pte_v = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mem_resp_valid = _RAND_21[0:0];
  _RAND_22 = {2{`RANDOM}};
  mem_resp_data = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  line_988_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  line_989_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  line_990_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  state_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  tags__0 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  tags__1 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  data__0 = _RAND_30[19:0];
  _RAND_31 = {1{`RANDOM}};
  data__1 = _RAND_31[19:0];
  _RAND_32 = {1{`RANDOM}};
  line_991_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  line_992_valid_reg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  line_993_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  line_994_valid_reg = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  line_995_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_996_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_997_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_998_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  pte_hit = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_999_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_1000_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_1001_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_1002_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_1003_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_1004_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_1005_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_1006_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_1007_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_1008_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_1009_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_1010_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_1011_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_1012_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_1013_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_1014_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_1015_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_1016_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_1017_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_1018_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_1019_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_1020_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_1021_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_1022_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_1023_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_1024_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_1025_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_1026_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_1027_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_1028_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_1029_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_1030_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_1031_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  line_1032_valid_reg = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_1033_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_1034_valid_reg = _RAND_76[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(io_dpath_perf_l2hit & (io_dpath_perf_pte_miss | io_dpath_perf_pte_hit))); // @[src/main/scala/rocket/PTW.scala 407:9]
    end
    //
    if (_T_76 & _T_77 & _T_74) begin
      assert(~arb_io_out_bits_bits_need_gpa); // @[src/main/scala/rocket/PTW.scala 622:15]
    end
    //
    if (mem_resp_valid & _T_74) begin
      assert(state == 3'h5); // @[src/main/scala/rocket/PTW.scala 701:11]
    end
    //
    if (io_mem_s2_nack & _T_74) begin
      assert(state == 3'h4); // @[src/main/scala/rocket/PTW.scala 745:11]
    end
  end
endmodule
module RVCExpander(
  input         clock,
  input         reset,
  input  [31:0] io_in, // @[src/main/scala/rocket/RVC.scala 159:14]
  output [31:0] io_out_bits, // @[src/main/scala/rocket/RVC.scala 159:14]
  output [4:0]  io_out_rd, // @[src/main/scala/rocket/RVC.scala 159:14]
  output [4:0]  io_out_rs1, // @[src/main/scala/rocket/RVC.scala 159:14]
  output [4:0]  io_out_rs2, // @[src/main/scala/rocket/RVC.scala 159:14]
  output        io_rvc // @[src/main/scala/rocket/RVC.scala 159:14]
);
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f; // @[src/main/scala/rocket/RVC.scala 53:20]
  wire [4:0] _io_out_s_T_6 = {2'h1,io_in[4:2]}; // @[src/main/scala/rocket/RVC.scala 31:17]
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc}; // @[src/main/scala/rocket/RVC.scala 54:15]
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0}; // @[src/main/scala/rocket/RVC.scala 36:18]
  wire [4:0] _io_out_s_T_17 = {2'h1,io_in[9:7]}; // @[src/main/scala/rocket/RVC.scala 30:17]
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[src/main/scala/rocket/RVC.scala 58:23]
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[src/main/scala/rocket/RVC.scala 35:18]
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/rocket/RVC.scala 57:22]
  wire [27:0] _io_out_s_T_51 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/rocket/RVC.scala 56:22]
  wire [26:0] _io_out_s_T_73 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f}; // @[src/main/scala/rocket/RVC.scala 63:25]
  wire [27:0] _io_out_s_T_93 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27}; // @[src/main/scala/rocket/RVC.scala 66:23]
  wire [26:0] _io_out_s_T_115 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23}; // @[src/main/scala/rocket/RVC.scala 65:22]
  wire [27:0] _io_out_s_T_135 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h23}; // @[src/main/scala/rocket/RVC.scala 64:22]
  wire [6:0] _io_out_s_T_144 = io_in[12] ? 7'h7f : 7'h0; // @[src/main/scala/rocket/RVC.scala 43:25]
  wire [11:0] _io_out_s_T_146 = {_io_out_s_T_144,io_in[6:2]}; // @[src/main/scala/rocket/RVC.scala 43:20]
  wire [31:0] io_out_s_8_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/rocket/RVC.scala 75:24]
  wire  _io_out_s_opc_T_3 = |io_in[11:7]; // @[src/main/scala/rocket/RVC.scala 77:24]
  wire [6:0] io_out_s_opc_1 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[src/main/scala/rocket/RVC.scala 77:20]
  wire [31:0] io_out_s_9_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],io_out_s_opc_1}; // @[src/main/scala/rocket/RVC.scala 78:15]
  wire [31:0] io_out_s_10_bits = {_io_out_s_T_144,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[src/main/scala/rocket/RVC.scala 84:22]
  wire  _io_out_s_opc_T_8 = |_io_out_s_T_146; // @[src/main/scala/rocket/RVC.scala 90:29]
  wire [6:0] io_out_s_opc_2 = |_io_out_s_T_146 ? 7'h37 : 7'h3f; // @[src/main/scala/rocket/RVC.scala 90:20]
  wire [14:0] _io_out_s_me_T_1 = io_in[12] ? 15'h7fff : 15'h0; // @[src/main/scala/rocket/RVC.scala 41:24]
  wire [31:0] _io_out_s_me_T_3 = {_io_out_s_me_T_1,io_in[6:2],12'h0}; // @[src/main/scala/rocket/RVC.scala 41:19]
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_3[31:12],io_in[11:7],io_out_s_opc_2}; // @[src/main/scala/rocket/RVC.scala 91:24]
  wire [6:0] io_out_s_opc_3 = _io_out_s_opc_T_8 ? 7'h13 : 7'h1f; // @[src/main/scala/rocket/RVC.scala 86:20]
  wire [2:0] _io_out_s_T_183 = io_in[12] ? 3'h7 : 3'h0; // @[src/main/scala/rocket/RVC.scala 42:29]
  wire [31:0] io_out_s_res_bits = {_io_out_s_T_183,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:
    7],io_out_s_opc_3}; // @[src/main/scala/rocket/RVC.scala 87:15]
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_bits : io_out_s_me_bits; // @[src/main/scala/rocket/RVC.scala 92:10]
  wire [4:0] io_out_s_11_rd = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_in[11:7] : io_in[11:7]; // @[src/main/scala/rocket/RVC.scala 92:10]
  wire [4:0] io_out_s_11_rs2 = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? _io_out_s_T_6 : _io_out_s_T_6; // @[src/main/scala/rocket/RVC.scala 92:10]
  wire [25:0] _io_out_s_T_204 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/rocket/RVC.scala 98:21]
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_204}; // @[src/main/scala/rocket/RVC.scala 99:23]
  wire [30:0] _io_out_s_T_213 = _GEN_0 | 31'h40000000; // @[src/main/scala/rocket/RVC.scala 99:23]
  wire [31:0] _io_out_s_T_222 = {_io_out_s_T_144,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/rocket/RVC.scala 100:21]
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]}; // @[src/main/scala/rocket/RVC.scala 102:68]
  wire [2:0] _io_out_s_funct_T_4 = _io_out_s_funct_T_2 == 3'h1 ? 3'h4 : 3'h0; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] _io_out_s_funct_T_6 = _io_out_s_funct_T_2 == 3'h2 ? 3'h6 : _io_out_s_funct_T_4; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] _io_out_s_funct_T_8 = _io_out_s_funct_T_2 == 3'h3 ? 3'h7 : _io_out_s_funct_T_6; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] _io_out_s_funct_T_10 = _io_out_s_funct_T_2 == 3'h4 ? 3'h0 : _io_out_s_funct_T_8; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] _io_out_s_funct_T_12 = _io_out_s_funct_T_2 == 3'h5 ? 3'h0 : _io_out_s_funct_T_10; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] _io_out_s_funct_T_14 = _io_out_s_funct_T_2 == 3'h6 ? 3'h2 : _io_out_s_funct_T_12; // @[src/main/scala/util/package.scala 33:76]
  wire [2:0] io_out_s_funct = _io_out_s_funct_T_2 == 3'h7 ? 3'h3 : _io_out_s_funct_T_14; // @[src/main/scala/util/package.scala 33:76]
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[src/main/scala/rocket/RVC.scala 103:22]
  wire [6:0] io_out_s_opc_4 = io_in[12] ? 7'h3b : 7'h33; // @[src/main/scala/rocket/RVC.scala 104:22]
  wire [24:0] _io_out_s_T_229 = {2'h1,io_in[4:2],2'h1,io_in[9:7],io_out_s_funct,2'h1,io_in[9:7],io_out_s_opc_4}; // @[src/main/scala/rocket/RVC.scala 105:12]
  wire [30:0] _GEN_1 = {{6'd0}, _io_out_s_T_229}; // @[src/main/scala/rocket/RVC.scala 105:43]
  wire [30:0] _io_out_s_T_230 = _GEN_1 | io_out_s_sub; // @[src/main/scala/rocket/RVC.scala 105:43]
  wire [30:0] _io_out_s_T_233 = io_in[11:10] == 2'h1 ? _io_out_s_T_213 : {{5'd0}, _io_out_s_T_204}; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_s_T_235 = io_in[11:10] == 2'h2 ? _io_out_s_T_222 : {{1'd0}, _io_out_s_T_233}; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_12_bits = io_in[11:10] == 2'h3 ? {{1'd0}, _io_out_s_T_230} : _io_out_s_T_235; // @[src/main/scala/util/package.scala 33:76]
  wire [9:0] _io_out_s_T_246 = io_in[12] ? 10'h3ff : 10'h0; // @[src/main/scala/rocket/RVC.scala 44:22]
  wire [20:0] _io_out_s_T_254 = {_io_out_s_T_246,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    }; // @[src/main/scala/rocket/RVC.scala 44:17]
  wire [31:0] io_out_s_13_bits = {_io_out_s_T_254[20],_io_out_s_T_254[10:1],_io_out_s_T_254[11],_io_out_s_T_254[19:12],5'h0
    ,7'h6f}; // @[src/main/scala/rocket/RVC.scala 94:21]
  wire [4:0] _io_out_s_T_296 = io_in[12] ? 5'h1f : 5'h0; // @[src/main/scala/rocket/RVC.scala 45:22]
  wire [12:0] _io_out_s_T_301 = {_io_out_s_T_296,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[src/main/scala/rocket/RVC.scala 45:17]
  wire [31:0] io_out_s_14_bits = {_io_out_s_T_301[12],_io_out_s_T_301[10:5],5'h0,2'h1,io_in[9:7],3'h0,_io_out_s_T_301[4:
    1],_io_out_s_T_301[11],7'h63}; // @[src/main/scala/rocket/RVC.scala 95:24]
  wire [31:0] io_out_s_15_bits = {_io_out_s_T_301[12],_io_out_s_T_301[10:5],5'h0,2'h1,io_in[9:7],3'h1,_io_out_s_T_301[4:
    1],_io_out_s_T_301[11],7'h63}; // @[src/main/scala/rocket/RVC.scala 96:24]
  wire [6:0] io_out_s_load_opc = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[src/main/scala/rocket/RVC.scala 113:23]
  wire [25:0] _io_out_s_T_378 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[src/main/scala/rocket/RVC.scala 114:24]
  wire [28:0] _io_out_s_T_388 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[src/main/scala/rocket/RVC.scala 117:25]
  wire [27:0] _io_out_s_T_397 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/rocket/RVC.scala 116:24]
  wire [28:0] _io_out_s_T_406 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/rocket/RVC.scala 115:24]
  wire [24:0] _io_out_s_mv_T_2 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[src/main/scala/rocket/RVC.scala 132:22]
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[src/main/scala/rocket/RVC.scala 134:25]
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[src/main/scala/rocket/RVC.scala 135:19]
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f}; // @[src/main/scala/rocket/RVC.scala 136:25]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[src/main/scala/rocket/RVC.scala 137:33]
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2]; // @[src/main/scala/rocket/RVC.scala 138:27]
  wire [31:0] io_out_s_mv_bits = {{7'd0}, _io_out_s_mv_T_2}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[src/main/scala/rocket/RVC.scala 138:22]
  wire [4:0] io_out_s_jr_mv_rd = |io_in[6:2] ? io_in[11:7] : 5'h0; // @[src/main/scala/rocket/RVC.scala 138:22]
  wire [4:0] io_out_s_jr_mv_rs1 = |io_in[6:2] ? 5'h0 : io_in[11:7]; // @[src/main/scala/rocket/RVC.scala 138:22]
  wire [4:0] io_out_s_jr_mv_rs2 = |io_in[6:2] ? io_in[6:2] : io_in[6:2]; // @[src/main/scala/rocket/RVC.scala 138:22]
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[src/main/scala/rocket/RVC.scala 139:21]
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73}; // @[src/main/scala/rocket/RVC.scala 140:23]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000; // @[src/main/scala/rocket/RVC.scala 140:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[src/main/scala/rocket/RVC.scala 141:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[src/main/scala/rocket/RVC.scala 142:25]
  wire [4:0] io_out_s_jalr_add_rd = _io_out_s_jr_mv_T_1 ? io_in[11:7] : 5'h1; // @[src/main/scala/rocket/RVC.scala 142:25]
  wire [4:0] io_out_s_jalr_add_rs1 = _io_out_s_jr_mv_T_1 ? io_in[11:7] : io_in[11:7]; // @[src/main/scala/rocket/RVC.scala 142:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[src/main/scala/rocket/RVC.scala 143:10]
  wire [4:0] io_out_s_20_rd = io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd; // @[src/main/scala/rocket/RVC.scala 143:10]
  wire [4:0] io_out_s_20_rs1 = io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1; // @[src/main/scala/rocket/RVC.scala 143:10]
  wire [4:0] io_out_s_20_rs2 = io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2; // @[src/main/scala/rocket/RVC.scala 143:10]
  wire [8:0] _io_out_s_T_413 = {io_in[9:7],io_in[12:10],3'h0}; // @[src/main/scala/rocket/RVC.scala 40:20]
  wire [28:0] _io_out_s_T_420 = {_io_out_s_T_413[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_413[4:0],7'h27}; // @[src/main/scala/rocket/RVC.scala 124:25]
  wire [7:0] _io_out_s_T_426 = {io_in[8:7],io_in[12:9],2'h0}; // @[src/main/scala/rocket/RVC.scala 39:20]
  wire [27:0] _io_out_s_T_433 = {_io_out_s_T_426[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_426[4:0],7'h23}; // @[src/main/scala/rocket/RVC.scala 123:24]
  wire [28:0] _io_out_s_T_446 = {_io_out_s_T_413[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_413[4:0],7'h23}; // @[src/main/scala/rocket/RVC.scala 122:24]
  wire [4:0] io_out_s_24_rs1 = io_in[19:15]; // @[src/main/scala/rocket/RVC.scala 20:57]
  wire [4:0] io_out_s_24_rs2 = io_in[24:20]; // @[src/main/scala/rocket/RVC.scala 20:79]
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]}; // @[src/main/scala/rocket/RVC.scala 154:10]
  wire [31:0] io_out_s_1_bits = {{4'd0}, _io_out_s_T_20}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_0_bits = {{2'd0}, _io_out_s_T_7}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_4_bits = _io_out_T_2 == 5'h1 ? io_out_s_1_bits : io_out_s_0_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_4_rd = _io_out_T_2 == 5'h1 ? _io_out_s_T_6 : _io_out_s_T_6; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_4_rs1 = _io_out_T_2 == 5'h1 ? _io_out_s_T_17 : 5'h2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_2_bits = {{5'd0}, _io_out_s_T_36}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_6_bits = _io_out_T_2 == 5'h2 ? io_out_s_2_bits : _io_out_T_4_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_6_rd = _io_out_T_2 == 5'h2 ? _io_out_s_T_6 : _io_out_T_4_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_6_rs1 = _io_out_T_2 == 5'h2 ? _io_out_s_T_17 : _io_out_T_4_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_3_bits = {{4'd0}, _io_out_s_T_51}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_8_bits = _io_out_T_2 == 5'h3 ? io_out_s_3_bits : _io_out_T_6_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_8_rd = _io_out_T_2 == 5'h3 ? _io_out_s_T_6 : _io_out_T_6_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_8_rs1 = _io_out_T_2 == 5'h3 ? _io_out_s_T_17 : _io_out_T_6_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_4_bits = {{5'd0}, _io_out_s_T_73}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_10_bits = _io_out_T_2 == 5'h4 ? io_out_s_4_bits : _io_out_T_8_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_10_rd = _io_out_T_2 == 5'h4 ? _io_out_s_T_6 : _io_out_T_8_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_10_rs1 = _io_out_T_2 == 5'h4 ? _io_out_s_T_17 : _io_out_T_8_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_5_bits = {{4'd0}, _io_out_s_T_93}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_12_bits = _io_out_T_2 == 5'h5 ? io_out_s_5_bits : _io_out_T_10_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_12_rd = _io_out_T_2 == 5'h5 ? _io_out_s_T_6 : _io_out_T_10_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_12_rs1 = _io_out_T_2 == 5'h5 ? _io_out_s_T_17 : _io_out_T_10_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_6_bits = {{5'd0}, _io_out_s_T_115}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_14_bits = _io_out_T_2 == 5'h6 ? io_out_s_6_bits : _io_out_T_12_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_14_rd = _io_out_T_2 == 5'h6 ? _io_out_s_T_6 : _io_out_T_12_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_14_rs1 = _io_out_T_2 == 5'h6 ? _io_out_s_T_17 : _io_out_T_12_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_7_bits = {{4'd0}, _io_out_s_T_135}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_16_bits = _io_out_T_2 == 5'h7 ? io_out_s_7_bits : _io_out_T_14_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_16_rd = _io_out_T_2 == 5'h7 ? _io_out_s_T_6 : _io_out_T_14_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_16_rs1 = _io_out_T_2 == 5'h7 ? _io_out_s_T_17 : _io_out_T_14_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_18_bits = _io_out_T_2 == 5'h8 ? io_out_s_8_bits : _io_out_T_16_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_18_rd = _io_out_T_2 == 5'h8 ? io_in[11:7] : _io_out_T_16_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_18_rs1 = _io_out_T_2 == 5'h8 ? io_in[11:7] : _io_out_T_16_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_18_rs2 = _io_out_T_2 == 5'h8 ? _io_out_s_T_6 : _io_out_T_16_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_20_bits = _io_out_T_2 == 5'h9 ? io_out_s_9_bits : _io_out_T_18_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_20_rd = _io_out_T_2 == 5'h9 ? io_in[11:7] : _io_out_T_18_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_20_rs1 = _io_out_T_2 == 5'h9 ? io_in[11:7] : _io_out_T_18_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_20_rs2 = _io_out_T_2 == 5'h9 ? _io_out_s_T_6 : _io_out_T_18_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_22_bits = _io_out_T_2 == 5'ha ? io_out_s_10_bits : _io_out_T_20_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_22_rd = _io_out_T_2 == 5'ha ? io_in[11:7] : _io_out_T_20_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_22_rs1 = _io_out_T_2 == 5'ha ? 5'h0 : _io_out_T_20_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_22_rs2 = _io_out_T_2 == 5'ha ? _io_out_s_T_6 : _io_out_T_20_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_24_bits = _io_out_T_2 == 5'hb ? io_out_s_11_bits : _io_out_T_22_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_24_rd = _io_out_T_2 == 5'hb ? io_out_s_11_rd : _io_out_T_22_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_24_rs1 = _io_out_T_2 == 5'hb ? io_out_s_11_rd : _io_out_T_22_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_24_rs2 = _io_out_T_2 == 5'hb ? io_out_s_11_rs2 : _io_out_T_22_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_26_bits = _io_out_T_2 == 5'hc ? io_out_s_12_bits : _io_out_T_24_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_26_rd = _io_out_T_2 == 5'hc ? _io_out_s_T_17 : _io_out_T_24_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_26_rs1 = _io_out_T_2 == 5'hc ? _io_out_s_T_17 : _io_out_T_24_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_26_rs2 = _io_out_T_2 == 5'hc ? _io_out_s_T_6 : _io_out_T_24_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_28_bits = _io_out_T_2 == 5'hd ? io_out_s_13_bits : _io_out_T_26_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_28_rd = _io_out_T_2 == 5'hd ? 5'h0 : _io_out_T_26_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_28_rs1 = _io_out_T_2 == 5'hd ? _io_out_s_T_17 : _io_out_T_26_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_28_rs2 = _io_out_T_2 == 5'hd ? _io_out_s_T_6 : _io_out_T_26_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_30_bits = _io_out_T_2 == 5'he ? io_out_s_14_bits : _io_out_T_28_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_30_rd = _io_out_T_2 == 5'he ? _io_out_s_T_17 : _io_out_T_28_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_30_rs1 = _io_out_T_2 == 5'he ? _io_out_s_T_17 : _io_out_T_28_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_30_rs2 = _io_out_T_2 == 5'he ? 5'h0 : _io_out_T_28_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_32_bits = _io_out_T_2 == 5'hf ? io_out_s_15_bits : _io_out_T_30_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_32_rd = _io_out_T_2 == 5'hf ? 5'h0 : _io_out_T_30_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_32_rs1 = _io_out_T_2 == 5'hf ? _io_out_s_T_17 : _io_out_T_30_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_32_rs2 = _io_out_T_2 == 5'hf ? 5'h0 : _io_out_T_30_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_16_bits = {{6'd0}, _io_out_s_T_378}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_34_bits = _io_out_T_2 == 5'h10 ? io_out_s_16_bits : _io_out_T_32_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_34_rd = _io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_34_rs1 = _io_out_T_2 == 5'h10 ? io_in[11:7] : _io_out_T_32_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_34_rs2 = _io_out_T_2 == 5'h10 ? io_in[6:2] : _io_out_T_32_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_17_bits = {{3'd0}, _io_out_s_T_388}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_36_bits = _io_out_T_2 == 5'h11 ? io_out_s_17_bits : _io_out_T_34_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_36_rd = _io_out_T_2 == 5'h11 ? io_in[11:7] : _io_out_T_34_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_36_rs1 = _io_out_T_2 == 5'h11 ? 5'h2 : _io_out_T_34_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_36_rs2 = _io_out_T_2 == 5'h11 ? io_in[6:2] : _io_out_T_34_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_18_bits = {{4'd0}, _io_out_s_T_397}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_38_bits = _io_out_T_2 == 5'h12 ? io_out_s_18_bits : _io_out_T_36_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_38_rd = _io_out_T_2 == 5'h12 ? io_in[11:7] : _io_out_T_36_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_38_rs1 = _io_out_T_2 == 5'h12 ? 5'h2 : _io_out_T_36_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_38_rs2 = _io_out_T_2 == 5'h12 ? io_in[6:2] : _io_out_T_36_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_19_bits = {{3'd0}, _io_out_s_T_406}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_40_bits = _io_out_T_2 == 5'h13 ? io_out_s_19_bits : _io_out_T_38_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_40_rd = _io_out_T_2 == 5'h13 ? io_in[11:7] : _io_out_T_38_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_40_rs1 = _io_out_T_2 == 5'h13 ? 5'h2 : _io_out_T_38_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_40_rs2 = _io_out_T_2 == 5'h13 ? io_in[6:2] : _io_out_T_38_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_42_bits = _io_out_T_2 == 5'h14 ? io_out_s_20_bits : _io_out_T_40_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_42_rd = _io_out_T_2 == 5'h14 ? io_out_s_20_rd : _io_out_T_40_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_42_rs1 = _io_out_T_2 == 5'h14 ? io_out_s_20_rs1 : _io_out_T_40_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_42_rs2 = _io_out_T_2 == 5'h14 ? io_out_s_20_rs2 : _io_out_T_40_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_21_bits = {{3'd0}, _io_out_s_T_420}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_44_bits = _io_out_T_2 == 5'h15 ? io_out_s_21_bits : _io_out_T_42_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_44_rd = _io_out_T_2 == 5'h15 ? io_in[11:7] : _io_out_T_42_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_44_rs1 = _io_out_T_2 == 5'h15 ? 5'h2 : _io_out_T_42_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_44_rs2 = _io_out_T_2 == 5'h15 ? io_in[6:2] : _io_out_T_42_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_22_bits = {{4'd0}, _io_out_s_T_433}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_46_bits = _io_out_T_2 == 5'h16 ? io_out_s_22_bits : _io_out_T_44_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_46_rd = _io_out_T_2 == 5'h16 ? io_in[11:7] : _io_out_T_44_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_46_rs1 = _io_out_T_2 == 5'h16 ? 5'h2 : _io_out_T_44_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_46_rs2 = _io_out_T_2 == 5'h16 ? io_in[6:2] : _io_out_T_44_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] io_out_s_23_bits = {{3'd0}, _io_out_s_T_446}; // @[src/main/scala/rocket/RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_48_bits = _io_out_T_2 == 5'h17 ? io_out_s_23_bits : _io_out_T_46_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_48_rd = _io_out_T_2 == 5'h17 ? io_in[11:7] : _io_out_T_46_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_48_rs1 = _io_out_T_2 == 5'h17 ? 5'h2 : _io_out_T_46_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_48_rs2 = _io_out_T_2 == 5'h17 ? io_in[6:2] : _io_out_T_46_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_50_bits = _io_out_T_2 == 5'h18 ? io_in : _io_out_T_48_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_50_rd = _io_out_T_2 == 5'h18 ? io_in[11:7] : _io_out_T_48_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_50_rs1 = _io_out_T_2 == 5'h18 ? io_out_s_24_rs1 : _io_out_T_48_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_50_rs2 = _io_out_T_2 == 5'h18 ? io_out_s_24_rs2 : _io_out_T_48_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_52_bits = _io_out_T_2 == 5'h19 ? io_in : _io_out_T_50_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_52_rd = _io_out_T_2 == 5'h19 ? io_in[11:7] : _io_out_T_50_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_52_rs1 = _io_out_T_2 == 5'h19 ? io_out_s_24_rs1 : _io_out_T_50_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_52_rs2 = _io_out_T_2 == 5'h19 ? io_out_s_24_rs2 : _io_out_T_50_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_54_bits = _io_out_T_2 == 5'h1a ? io_in : _io_out_T_52_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_54_rd = _io_out_T_2 == 5'h1a ? io_in[11:7] : _io_out_T_52_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_54_rs1 = _io_out_T_2 == 5'h1a ? io_out_s_24_rs1 : _io_out_T_52_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_54_rs2 = _io_out_T_2 == 5'h1a ? io_out_s_24_rs2 : _io_out_T_52_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_56_bits = _io_out_T_2 == 5'h1b ? io_in : _io_out_T_54_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_56_rd = _io_out_T_2 == 5'h1b ? io_in[11:7] : _io_out_T_54_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_56_rs1 = _io_out_T_2 == 5'h1b ? io_out_s_24_rs1 : _io_out_T_54_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_56_rs2 = _io_out_T_2 == 5'h1b ? io_out_s_24_rs2 : _io_out_T_54_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_58_bits = _io_out_T_2 == 5'h1c ? io_in : _io_out_T_56_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_58_rd = _io_out_T_2 == 5'h1c ? io_in[11:7] : _io_out_T_56_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_58_rs1 = _io_out_T_2 == 5'h1c ? io_out_s_24_rs1 : _io_out_T_56_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_58_rs2 = _io_out_T_2 == 5'h1c ? io_out_s_24_rs2 : _io_out_T_56_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_60_bits = _io_out_T_2 == 5'h1d ? io_in : _io_out_T_58_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_60_rd = _io_out_T_2 == 5'h1d ? io_in[11:7] : _io_out_T_58_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_60_rs1 = _io_out_T_2 == 5'h1d ? io_out_s_24_rs1 : _io_out_T_58_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_60_rs2 = _io_out_T_2 == 5'h1d ? io_out_s_24_rs2 : _io_out_T_58_rs2; // @[src/main/scala/util/package.scala 33:76]
  wire [31:0] _io_out_T_62_bits = _io_out_T_2 == 5'h1e ? io_in : _io_out_T_60_bits; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_62_rd = _io_out_T_2 == 5'h1e ? io_in[11:7] : _io_out_T_60_rd; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_62_rs1 = _io_out_T_2 == 5'h1e ? io_out_s_24_rs1 : _io_out_T_60_rs1; // @[src/main/scala/util/package.scala 33:76]
  wire [4:0] _io_out_T_62_rs2 = _io_out_T_2 == 5'h1e ? io_out_s_24_rs2 : _io_out_T_60_rs2; // @[src/main/scala/util/package.scala 33:76]
  assign io_out_bits = _io_out_T_2 == 5'h1f ? io_in : _io_out_T_62_bits; // @[src/main/scala/util/package.scala 33:76]
  assign io_out_rd = _io_out_T_2 == 5'h1f ? io_in[11:7] : _io_out_T_62_rd; // @[src/main/scala/util/package.scala 33:76]
  assign io_out_rs1 = _io_out_T_2 == 5'h1f ? io_out_s_24_rs1 : _io_out_T_62_rs1; // @[src/main/scala/util/package.scala 33:76]
  assign io_out_rs2 = _io_out_T_2 == 5'h1f ? io_out_s_24_rs2 : _io_out_T_62_rs2; // @[src/main/scala/util/package.scala 33:76]
  assign io_rvc = io_in[1:0] != 2'h3; // @[src/main/scala/rocket/RVC.scala 166:26]
endmodule
module IBuf(
  input         clock,
  input         reset,
  output        io_imem_ready, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_imem_valid, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input  [39:0] io_imem_bits_pc, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input  [31:0] io_imem_bits_data, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_imem_bits_xcpt_pf_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_imem_bits_xcpt_ae_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_imem_bits_replay, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_kill, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [39:0] io_pc, // @[src/main/scala/rocket/IBuf.scala 22:14]
  input         io_inst_0_ready, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_valid, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_xcpt0_pf_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_xcpt0_ae_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_xcpt1_pf_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_xcpt1_gf_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_xcpt1_ae_inst, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_replay, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output        io_inst_0_bits_rvc, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [31:0] io_inst_0_bits_inst_bits, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [4:0]  io_inst_0_bits_inst_rd, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [4:0]  io_inst_0_bits_inst_rs1, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [4:0]  io_inst_0_bits_inst_rs2, // @[src/main/scala/rocket/IBuf.scala 22:14]
  output [31:0] io_inst_0_bits_raw // @[src/main/scala/rocket/IBuf.scala 22:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  exp_clock; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire  exp_reset; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire [31:0] exp_io_in; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire [31:0] exp_io_out_bits; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire [4:0] exp_io_out_rd; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire [4:0] exp_io_out_rs1; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire [4:0] exp_io_out_rs2; // @[src/main/scala/rocket/IBuf.scala 86:21]
  wire  exp_io_rvc; // @[src/main/scala/rocket/IBuf.scala 86:21]
  reg  nBufValid; // @[src/main/scala/rocket/IBuf.scala 34:47]
  reg [39:0] buf__pc; // @[src/main/scala/rocket/IBuf.scala 35:16]
  reg [31:0] buf__data; // @[src/main/scala/rocket/IBuf.scala 35:16]
  reg  buf__xcpt_pf_inst; // @[src/main/scala/rocket/IBuf.scala 35:16]
  reg  buf__xcpt_ae_inst; // @[src/main/scala/rocket/IBuf.scala 35:16]
  reg  buf__replay; // @[src/main/scala/rocket/IBuf.scala 35:16]
  wire  pcWordBits = io_imem_bits_pc[1]; // @[src/main/scala/util/package.scala 155:13]
  wire [1:0] _GEN_65 = {{1'd0}, pcWordBits}; // @[src/main/scala/rocket/IBuf.scala 41:86]
  wire [1:0] nIC = 2'h2 - _GEN_65; // @[src/main/scala/rocket/IBuf.scala 41:86]
  wire [1:0] _nValid_T = io_imem_valid ? nIC : 2'h0; // @[src/main/scala/rocket/IBuf.scala 43:19]
  wire [1:0] _GEN_66 = {{1'd0}, nBufValid}; // @[src/main/scala/rocket/IBuf.scala 43:45]
  wire [1:0] nValid = _nValid_T + _GEN_66; // @[src/main/scala/rocket/IBuf.scala 43:45]
  wire [3:0] _valid_T = 4'h1 << nValid; // @[src/main/scala/chisel3/util/OneHot.scala 58:35]
  wire [3:0] _valid_T_2 = _valid_T - 4'h1; // @[src/main/scala/rocket/IBuf.scala 74:33]
  wire [1:0] valid = _valid_T_2[1:0]; // @[src/main/scala/rocket/IBuf.scala 74:39]
  wire [1:0] _full_insn_T_2 = {{1'd0}, valid[1]}; // @[src/main/scala/rocket/IBuf.scala 93:42]
  wire [1:0] _bufMask_T = 2'h1 << nBufValid; // @[src/main/scala/chisel3/util/OneHot.scala 58:35]
  wire [1:0] bufMask = _bufMask_T - 2'h1; // @[src/main/scala/rocket/IBuf.scala 75:37]
  wire [1:0] buf_replay = buf__replay ? bufMask : 2'h0; // @[src/main/scala/rocket/IBuf.scala 77:23]
  wire  full_insn = exp_io_rvc | _full_insn_T_2[0] | buf_replay[0]; // @[src/main/scala/rocket/IBuf.scala 93:50]
  wire [1:0] _nReady_T_4 = exp_io_rvc ? 2'h1 : 2'h2; // @[src/main/scala/rocket/IBuf.scala 102:75]
  wire [1:0] nReady = full_insn ? _nReady_T_4 : 2'h0; // @[src/main/scala/rocket/IBuf.scala 102:{60,69} 40:27]
  wire [1:0] nICReady = nReady - _GEN_66; // @[src/main/scala/rocket/IBuf.scala 42:25]
  wire  _io_imem_ready_T = nReady >= _GEN_66; // @[src/main/scala/rocket/IBuf.scala 44:47]
  wire [1:0] _io_imem_ready_T_4 = nIC - nICReady; // @[src/main/scala/rocket/IBuf.scala 44:94]
  wire  _io_imem_ready_T_5 = 2'h1 >= _io_imem_ready_T_4; // @[src/main/scala/rocket/IBuf.scala 44:87]
  wire  line_1035_clock;
  wire  line_1035_reset;
  wire  line_1035_valid;
  reg  line_1035_valid_reg;
  wire  _nBufValid_T_2 = _io_imem_ready_T | ~nBufValid; // @[src/main/scala/util/package.scala 210:38]
  wire [1:0] _nBufValid_T_4 = _GEN_66 - nReady; // @[src/main/scala/rocket/IBuf.scala 48:61]
  wire [1:0] _nBufValid_T_5 = _nBufValid_T_2 ? 2'h0 : _nBufValid_T_4; // @[src/main/scala/rocket/IBuf.scala 48:23]
  wire  _T_7 = io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5; // @[src/main/scala/rocket/IBuf.scala 54:68]
  wire  line_1036_clock;
  wire  line_1036_reset;
  wire  line_1036_valid;
  reg  line_1036_valid_reg;
  wire [1:0] shamt = _GEN_65 + nICReady; // @[src/main/scala/rocket/IBuf.scala 55:32]
  wire [63:0] buf_data_data = {io_imem_bits_data[31:16],io_imem_bits_data[31:16],io_imem_bits_data}; // @[src/main/scala/rocket/IBuf.scala 127:19]
  wire [5:0] _buf_data_T = {shamt, 4'h0}; // @[src/main/scala/rocket/IBuf.scala 128:19]
  wire [63:0] _buf_data_T_1 = buf_data_data >> _buf_data_T; // @[src/main/scala/rocket/IBuf.scala 128:10]
  wire [39:0] _buf_pc_T_1 = io_imem_bits_pc & 40'hfffffffffc; // @[src/main/scala/rocket/IBuf.scala 59:35]
  wire [2:0] _buf_pc_T_2 = {nICReady, 1'h0}; // @[src/main/scala/rocket/IBuf.scala 59:80]
  wire [39:0] _GEN_74 = {{37'd0}, _buf_pc_T_2}; // @[src/main/scala/rocket/IBuf.scala 59:68]
  wire [39:0] _buf_pc_T_4 = io_imem_bits_pc + _GEN_74; // @[src/main/scala/rocket/IBuf.scala 59:68]
  wire [39:0] _buf_pc_T_5 = _buf_pc_T_4 & 40'h3; // @[src/main/scala/rocket/IBuf.scala 59:109]
  wire [39:0] _buf_pc_T_6 = _buf_pc_T_1 | _buf_pc_T_5; // @[src/main/scala/rocket/IBuf.scala 59:49]
  wire [1:0] _GEN_7 = io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5 ? _io_imem_ready_T_4 :
    _nBufValid_T_5; // @[src/main/scala/rocket/IBuf.scala 48:17 54:94 56:19]
  wire [1:0] _GEN_31 = io_inst_0_ready ? _GEN_7 : {{1'd0}, nBufValid}; // @[src/main/scala/rocket/IBuf.scala 47:29 34:47]
  wire  line_1037_clock;
  wire  line_1037_reset;
  wire  line_1037_valid;
  reg  line_1037_valid_reg;
  wire [1:0] _GEN_55 = io_kill ? 2'h0 : _GEN_31; // @[src/main/scala/rocket/IBuf.scala 63:20 64:17]
  wire [1:0] _icShiftAmt_T_1 = 2'h2 + _GEN_66; // @[src/main/scala/rocket/IBuf.scala 68:34]
  wire [1:0] icShiftAmt = _icShiftAmt_T_1 - _GEN_65; // @[src/main/scala/rocket/IBuf.scala 68:46]
  wire [63:0] _icData_T_2 = {io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[src/main/scala/rocket/IBuf.scala 69:33]
  wire [127:0] icData_data = {_icData_T_2[63:48],_icData_T_2[63:48],_icData_T_2[63:48],_icData_T_2[63:48],
    io_imem_bits_data,io_imem_bits_data[15:0],io_imem_bits_data[15:0]}; // @[src/main/scala/rocket/IBuf.scala 120:19]
  wire [5:0] _icData_T_3 = {icShiftAmt, 4'h0}; // @[src/main/scala/rocket/IBuf.scala 121:19]
  wire [190:0] _GEN_8 = {{63'd0}, icData_data}; // @[src/main/scala/rocket/IBuf.scala 121:10]
  wire [190:0] _icData_T_4 = _GEN_8 << _icData_T_3; // @[src/main/scala/rocket/IBuf.scala 121:10]
  wire [31:0] icData = _icData_T_4[95:64]; // @[src/main/scala/util/package.scala 155:13]
  wire [4:0] _icMask_T_1 = {nBufValid, 4'h0}; // @[src/main/scala/rocket/IBuf.scala 71:65]
  wire [62:0] _icMask_T_2 = 63'hffffffff << _icMask_T_1; // @[src/main/scala/rocket/IBuf.scala 71:51]
  wire [31:0] icMask = _icMask_T_2[31:0]; // @[src/main/scala/rocket/IBuf.scala 71:92]
  wire [31:0] _inst_T = icData & icMask; // @[src/main/scala/rocket/IBuf.scala 72:21]
  wire [31:0] _inst_T_1 = ~icMask; // @[src/main/scala/rocket/IBuf.scala 72:43]
  wire [31:0] _inst_T_2 = buf__data & _inst_T_1; // @[src/main/scala/rocket/IBuf.scala 72:41]
  wire  xcpt_1_pf_inst = bufMask[1] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[src/main/scala/rocket/IBuf.scala 76:53]
  wire  xcpt_1_ae_inst = bufMask[1] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[src/main/scala/rocket/IBuf.scala 76:53]
  wire [1:0] _ic_replay_T = ~bufMask; // @[src/main/scala/rocket/IBuf.scala 78:65]
  wire [1:0] _ic_replay_T_1 = valid & _ic_replay_T; // @[src/main/scala/rocket/IBuf.scala 78:63]
  wire [1:0] _ic_replay_T_2 = io_imem_bits_replay ? _ic_replay_T_1 : 2'h0; // @[src/main/scala/rocket/IBuf.scala 78:35]
  wire [1:0] ic_replay = buf_replay | _ic_replay_T_2; // @[src/main/scala/rocket/IBuf.scala 78:30]
  wire  _T_14 = ~reset; // @[src/main/scala/rocket/IBuf.scala 79:9]
  wire  line_1038_clock;
  wire  line_1038_reset;
  wire  line_1038_valid;
  reg  line_1038_valid_reg;
  wire [1:0] _replay_T_5 = {{1'd0}, ic_replay[1]}; // @[src/main/scala/rocket/IBuf.scala 92:61]
  wire [2:0] _io_inst_0_bits_xcpt1_T_4 = {xcpt_1_pf_inst,1'h0,xcpt_1_ae_inst}; // @[src/main/scala/rocket/IBuf.scala 96:65]
  wire [2:0] _io_inst_0_bits_xcpt1_T_5 = exp_io_rvc ? 3'h0 : _io_inst_0_bits_xcpt1_T_4; // @[src/main/scala/rocket/IBuf.scala 96:35]
  wire [1:0] _T_21 = {{1'd0}, bufMask[1]}; // @[src/main/scala/rocket/IBuf.scala 100:50]
  wire  _T_23 = bufMask[0] & exp_io_rvc | _T_21[0]; // @[src/main/scala/rocket/IBuf.scala 100:40]
  wire  line_1039_clock;
  wire  line_1039_reset;
  wire  line_1039_valid;
  reg  line_1039_valid_reg;
  wire  line_1040_clock;
  wire  line_1040_reset;
  wire  line_1040_valid;
  reg  line_1040_valid_reg;
  wire [1:0] _GEN_79 = reset ? 2'h0 : _GEN_55; // @[src/main/scala/rocket/IBuf.scala 34:{47,47}]
  RVCExpander exp ( // @[src/main/scala/rocket/IBuf.scala 86:21]
    .clock(exp_clock),
    .reset(exp_reset),
    .io_in(exp_io_in),
    .io_out_bits(exp_io_out_bits),
    .io_out_rd(exp_io_out_rd),
    .io_out_rs1(exp_io_out_rs1),
    .io_out_rs2(exp_io_out_rs2),
    .io_rvc(exp_io_rvc)
  );
  GEN_w1_line #(.COVER_INDEX(1035)) line_1035 (
    .clock(line_1035_clock),
    .reset(line_1035_reset),
    .valid(line_1035_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1036)) line_1036 (
    .clock(line_1036_clock),
    .reset(line_1036_reset),
    .valid(line_1036_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1037)) line_1037 (
    .clock(line_1037_clock),
    .reset(line_1037_reset),
    .valid(line_1037_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1038)) line_1038 (
    .clock(line_1038_clock),
    .reset(line_1038_reset),
    .valid(line_1038_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1039)) line_1039 (
    .clock(line_1039_clock),
    .reset(line_1039_reset),
    .valid(line_1039_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1040)) line_1040 (
    .clock(line_1040_clock),
    .reset(line_1040_reset),
    .valid(line_1040_valid)
  );
  assign line_1035_clock = clock;
  assign line_1035_reset = reset;
  assign line_1035_valid = io_inst_0_ready ^ line_1035_valid_reg;
  assign line_1036_clock = clock;
  assign line_1036_reset = reset;
  assign line_1036_valid = _T_7 ^ line_1036_valid_reg;
  assign line_1037_clock = clock;
  assign line_1037_reset = reset;
  assign line_1037_valid = io_kill ^ line_1037_valid_reg;
  assign line_1038_clock = clock;
  assign line_1038_reset = reset;
  assign line_1038_valid = _T_14 ^ line_1038_valid_reg;
  assign line_1039_clock = clock;
  assign line_1039_reset = reset;
  assign line_1039_valid = _T_23 ^ line_1039_valid_reg;
  assign line_1040_clock = clock;
  assign line_1040_reset = reset;
  assign line_1040_valid = full_insn ^ line_1040_valid_reg;
  assign io_imem_ready = io_inst_0_ready & nReady >= _GEN_66 & (nICReady >= nIC | 2'h1 >= _io_imem_ready_T_4); // @[src/main/scala/rocket/IBuf.scala 44:60]
  assign io_pc = nBufValid > 1'h0 ? buf__pc : io_imem_bits_pc; // @[src/main/scala/rocket/IBuf.scala 82:15]
  assign io_inst_0_valid = valid[0] & full_insn; // @[src/main/scala/rocket/IBuf.scala 94:36]
  assign io_inst_0_bits_xcpt0_pf_inst = bufMask[0] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[src/main/scala/rocket/IBuf.scala 76:53]
  assign io_inst_0_bits_xcpt0_ae_inst = bufMask[0] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[src/main/scala/rocket/IBuf.scala 76:53]
  assign io_inst_0_bits_xcpt1_pf_inst = _io_inst_0_bits_xcpt1_T_5[2]; // @[src/main/scala/rocket/IBuf.scala 96:81]
  assign io_inst_0_bits_xcpt1_gf_inst = _io_inst_0_bits_xcpt1_T_5[1]; // @[src/main/scala/rocket/IBuf.scala 96:81]
  assign io_inst_0_bits_xcpt1_ae_inst = _io_inst_0_bits_xcpt1_T_5[0]; // @[src/main/scala/rocket/IBuf.scala 96:81]
  assign io_inst_0_bits_replay = ic_replay[0] | ~exp_io_rvc & _replay_T_5[0]; // @[src/main/scala/rocket/IBuf.scala 92:33]
  assign io_inst_0_bits_rvc = exp_io_rvc; // @[src/main/scala/rocket/IBuf.scala 98:27]
  assign io_inst_0_bits_inst_bits = exp_io_out_bits; // @[src/main/scala/rocket/IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rd = exp_io_out_rd; // @[src/main/scala/rocket/IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs1 = exp_io_out_rs1; // @[src/main/scala/rocket/IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs2 = exp_io_out_rs2; // @[src/main/scala/rocket/IBuf.scala 88:26]
  assign io_inst_0_bits_raw = _inst_T | _inst_T_2; // @[src/main/scala/rocket/IBuf.scala 72:30]
  assign exp_clock = clock;
  assign exp_reset = reset;
  assign exp_io_in = _inst_T | _inst_T_2; // @[src/main/scala/rocket/IBuf.scala 72:30]
  always @(posedge clock) begin
    nBufValid <= _GEN_79[0]; // @[src/main/scala/rocket/IBuf.scala 34:{47,47}]
    if (io_inst_0_ready) begin // @[src/main/scala/rocket/IBuf.scala 47:29]
      if (io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5) begin // @[src/main/scala/rocket/IBuf.scala 54:94]
        buf__pc <= _buf_pc_T_6; // @[src/main/scala/rocket/IBuf.scala 59:16]
      end
    end
    if (io_inst_0_ready) begin // @[src/main/scala/rocket/IBuf.scala 47:29]
      if (io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5) begin // @[src/main/scala/rocket/IBuf.scala 54:94]
        buf__data <= {{16'd0}, _buf_data_T_1[15:0]}; // @[src/main/scala/rocket/IBuf.scala 58:18]
      end
    end
    if (io_inst_0_ready) begin // @[src/main/scala/rocket/IBuf.scala 47:29]
      if (io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5) begin // @[src/main/scala/rocket/IBuf.scala 54:94]
        buf__xcpt_pf_inst <= io_imem_bits_xcpt_pf_inst; // @[src/main/scala/rocket/IBuf.scala 57:13]
      end
    end
    if (io_inst_0_ready) begin // @[src/main/scala/rocket/IBuf.scala 47:29]
      if (io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5) begin // @[src/main/scala/rocket/IBuf.scala 54:94]
        buf__xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst; // @[src/main/scala/rocket/IBuf.scala 57:13]
      end
    end
    if (io_inst_0_ready) begin // @[src/main/scala/rocket/IBuf.scala 47:29]
      if (io_imem_valid & _io_imem_ready_T & nICReady < nIC & _io_imem_ready_T_5) begin // @[src/main/scala/rocket/IBuf.scala 54:94]
        buf__replay <= io_imem_bits_replay; // @[src/main/scala/rocket/IBuf.scala 57:13]
      end
    end
    line_1035_valid_reg <= io_inst_0_ready;
    line_1036_valid_reg <= _T_7;
    line_1037_valid_reg <= io_kill;
    line_1038_valid_reg <= _T_14;
    line_1039_valid_reg <= _T_23;
    line_1040_valid_reg <= full_insn;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  nBufValid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  buf__pc = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  buf__data = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buf__xcpt_pf_inst = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buf__xcpt_ae_inst = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  buf__replay = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1035_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1036_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1037_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1038_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1039_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1040_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/rocket/IBuf.scala 79:9]
    end
  end
endmodule
module DelayReg_2(
  input         clock,
  input         reset,
  input         i_valid, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [31:0] i_interrupt, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [31:0] i_exception, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [63:0] i_exceptionPC, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [31:0] i_exceptionInst, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  output        o_valid, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [31:0] o_interrupt, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [31:0] o_exception, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [63:0] o_exceptionPC, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [31:0] o_exceptionInst // @[difftest/src/main/scala/util/Delayer.scala 24:13]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [31:0] REG_interrupt; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [31:0] REG_exception; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_exceptionPC; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [31:0] REG_exceptionInst; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  assign o_valid = REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_interrupt = REG_interrupt; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_exception = REG_exception; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_exceptionPC = REG_exceptionPC; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_exceptionInst = REG_exceptionInst; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_valid <= i_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_interrupt <= 32'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_interrupt <= i_interrupt; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_exception <= 32'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_exception <= i_exception; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_exceptionPC <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_exceptionPC <= i_exceptionPC; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_exceptionInst <= 32'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_exceptionInst <= i_exceptionInst; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_interrupt = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  REG_exception = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  REG_exceptionPC = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  REG_exceptionInst = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_2(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_interrupt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exception, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_exceptionPC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exceptionInst // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_interrupt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exception; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_interrupt(dpic_io_interrupt),
    .io_exception(dpic_io_exception),
    .io_exceptionPC(dpic_io_exceptionPC),
    .io_exceptionInst(dpic_io_exceptionInst),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_interrupt = io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exception = io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionPC = io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionInst = io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_3(
  input         clock,
  input         reset,
  input         io_bits_hasTrap, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_cycleCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_instrCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasTrap; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_instrCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasWFI; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_code; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestTrapEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_hasTrap(dpic_io_hasTrap),
    .io_cycleCnt(dpic_io_cycleCnt),
    .io_instrCnt(dpic_io_instrCnt),
    .io_hasWFI(dpic_io_hasWFI),
    .io_code(dpic_io_code),
    .io_pc(dpic_io_pc),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_hasTrap = io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_cycleCnt = io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instrCnt = io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_hasWFI = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_code = 32'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_ungated_clock, // @[src/main/scala/rocket/CSR.scala 390:14]
  input         io_hartid, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [11:0] io_rw_addr, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [2:0]  io_rw_cmd, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_rw_rdata, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [63:0] io_rw_wdata, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [31:0] io_decode_0_inst, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_fp_illegal, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_fp_csr, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_rocc_illegal, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_read_illegal, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_write_illegal, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_write_flush, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_decode_0_system_illegal, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_csr_stall, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_rw_stall, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_eret, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_singleStep, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_debug, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_cease, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_wfi, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [31:0] io_status_isa, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_dprv, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_dv, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_prv, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_v, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_sd, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [22:0] io_status_zero2, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mpv, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_gva, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mbe, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_sbe, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_sxl, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_uxl, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_sd_rv32, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [7:0]  io_status_zero1, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_tsr, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_tw, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_tvm, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mxr, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_sum, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mprv, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_xs, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_fs, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_mpp, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [1:0]  io_status_vs, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_spp, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mpie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_ube, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_spie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_upie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_mie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_hie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_sie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_status_uie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [3:0]  io_ptbr_mode, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [43:0] io_ptbr_ppn, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [39:0] io_evec, // @[src/main/scala/rocket/CSR.scala 390:14]
  input         io_exception, // @[src/main/scala/rocket/CSR.scala 390:14]
  input         io_retire, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [63:0] io_cause, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [39:0] io_pc, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [39:0] io_tval, // @[src/main/scala/rocket/CSR.scala 390:14]
  input         io_gva, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_time, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_interrupt, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_interrupt_cause, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_csrr_counter, // @[src/main/scala/rocket/CSR.scala 390:14]
  input  [31:0] io_inst_0, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_trace_0_valid, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [39:0] io_trace_0_iaddr, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [31:0] io_trace_0_insn, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_trace_0_exception, // @[src/main/scala/rocket/CSR.scala 390:14]
  output        io_trace_0_interrupt, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_privilegeMode, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mstatus, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_sstatus, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mepc, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_sepc, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mtval, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_stval, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mtvec, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_stvec, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mcause, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_scause, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_satp, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mip, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mie, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mscratch, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_sscratch, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_mideleg, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_difftest_medeleg, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_snapshot_minstret, // @[src/main/scala/rocket/CSR.scala 390:14]
  output [63:0] io_snapshot_mcycle // @[src/main/scala/rocket/CSR.scala 390:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [63:0] _RAND_112;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_delayer_clock; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_reset; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_i_interrupt; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_i_exception; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_i_exceptionPC; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_i_exceptionInst; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_o_interrupt; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_o_exception; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_o_exceptionPC; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_o_exceptionInst; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [1:0] reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_gva; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_tsr; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_tw; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_tvm; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_mxr; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_sum; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_mprv; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg [1:0] reg_mstatus_fs; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg [1:0] reg_mstatus_mpp; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_spp; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_mpie; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 401:28]
  reg  reg_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 401:28]
  wire  system_insn = io_rw_cmd == 3'h4; // @[src/main/scala/rocket/CSR.scala 877:31]
  wire [31:0] _insn_T = {io_rw_addr, 20'h0}; // @[src/main/scala/rocket/CSR.scala 893:44]
  wire [31:0] insn = 32'h73 | _insn_T; // @[src/main/scala/rocket/CSR.scala 893:30]
  wire [31:0] decoded_invInputs = ~insn; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[20]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_1 = decoded_invInputs[21]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_2 = decoded_invInputs[22]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_3 = decoded_invInputs[23]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_4 = decoded_invInputs[24]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_5 = decoded_invInputs[25]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_6 = decoded_invInputs[26]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_7 = decoded_invInputs[27]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_8 = decoded_invInputs[28]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_9 = decoded_invInputs[29]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_10 = decoded_invInputs[30]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_11 = decoded_invInputs[31]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [5:0] decoded_lo = {decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_8,
    decoded_andMatrixInput_9,decoded_andMatrixInput_10,decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_T = {decoded_andMatrixInput_0,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_lo}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_1 = &_decoded_T; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_1; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  decoded_andMatrixInput_0_1 = insn[20]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [11:0] _decoded_T_2 = {decoded_andMatrixInput_0_1,decoded_andMatrixInput_1,decoded_andMatrixInput_2,
    decoded_andMatrixInput_3,decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_lo}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_3 = &_decoded_T_2; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_T_3; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  decoded_andMatrixInput_0_2 = insn[0]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_7_2 = insn[28]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _decoded_T_4 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_2,decoded_andMatrixInput_3,
    decoded_andMatrixInput_4,decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,
    decoded_andMatrixInput_7_2,decoded_andMatrixInput_10,decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_5 = &_decoded_T_4; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_6 = insn[30]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [1:0] _decoded_T_12 = {decoded_andMatrixInput_0_6,decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_13 = &_decoded_T_12; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [1:0] _decoded_orMatrixOutputs_T_3 = {_decoded_T_5,_decoded_T_13}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _decoded_orMatrixOutputs_T_4 = |_decoded_orMatrixOutputs_T_3; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  decoded_andMatrixInput_0_5 = insn[22]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_7_5 = insn[29]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _decoded_T_10 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_3,decoded_andMatrixInput_4,
    decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,
    decoded_andMatrixInput_7_5,decoded_andMatrixInput_10,decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_11 = &_decoded_T_10; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T_2 = |_decoded_T_11; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [9:0] _decoded_T_6 = {decoded_andMatrixInput_0_5,decoded_andMatrixInput_3,decoded_andMatrixInput_4,
    decoded_andMatrixInput_5,decoded_andMatrixInput_6,decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,
    decoded_andMatrixInput_9,decoded_andMatrixInput_10,decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_7 = &_decoded_T_6; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_T_7; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  decoded_andMatrixInput_1_4 = insn[1]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_2_4 = decoded_invInputs[2]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_3_4 = decoded_invInputs[3]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_4_4 = insn[4]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_5_4 = insn[5]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_6_4 = insn[6]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_7_4 = decoded_invInputs[7]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_8_4 = decoded_invInputs[8]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_9_4 = decoded_invInputs[9]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_10_2 = insn[25]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] decoded_lo_4 = {decoded_andMatrixInput_9_4,decoded_andMatrixInput_10_2,decoded_andMatrixInput_6,
    decoded_andMatrixInput_7,decoded_andMatrixInput_7_2,decoded_andMatrixInput_9,decoded_andMatrixInput_10,
    decoded_andMatrixInput_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [16:0] _decoded_T_8 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_1_4,decoded_andMatrixInput_2_4,
    decoded_andMatrixInput_3_4,decoded_andMatrixInput_4_4,decoded_andMatrixInput_5_4,decoded_andMatrixInput_6_4,
    decoded_andMatrixInput_7_4,decoded_andMatrixInput_8_4,decoded_lo_4}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_9 = &_decoded_T_8; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T = |_decoded_T_9; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [8:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,
    _decoded_orMatrixOutputs_T_4,_decoded_orMatrixOutputs_T_2,_decoded_orMatrixOutputs_T_1,_decoded_orMatrixOutputs_T,1'h0
    ,2'h0}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [8:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[8],decoded_orMatrixOutputs[7],decoded_orMatrixOutputs[6
    ],decoded_orMatrixOutputs[5],decoded_orMatrixOutputs[4],decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],
    decoded_orMatrixOutputs[1],decoded_orMatrixOutputs[0]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire  insn_ret = system_insn & decoded_invMatrixOutputs[6]; // @[src/main/scala/rocket/CSR.scala 894:83]
  wire  _T_368 = ~io_rw_addr[9]; // @[src/main/scala/rocket/CSR.scala 1114:32]
  wire  _T_374 = io_rw_addr[10] & io_rw_addr[7]; // @[src/main/scala/rocket/CSR.scala 1131:48]
  reg [1:0] reg_dcsr_prv; // @[src/main/scala/rocket/CSR.scala 409:25]
  wire [1:0] _GEN_276 = io_rw_addr[10] & io_rw_addr[7] ? reg_dcsr_prv : reg_mstatus_mpp; // @[src/main/scala/rocket/CSR.scala 1131:66 1132:15]
  wire [1:0] ret_prv = ~io_rw_addr[9] ? {{1'd0}, reg_mstatus_spp} : _GEN_276; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire  insn_call = system_insn & decoded_invMatrixOutputs[8]; // @[src/main/scala/rocket/CSR.scala 894:83]
  wire  insn_break = system_insn & decoded_invMatrixOutputs[7]; // @[src/main/scala/rocket/CSR.scala 894:83]
  wire  _exception_T = insn_call | insn_break; // @[src/main/scala/rocket/CSR.scala 1019:29]
  wire  exception = insn_call | insn_break | io_exception; // @[src/main/scala/rocket/CSR.scala 1019:43]
  reg  reg_singleStepped; // @[src/main/scala/rocket/CSR.scala 492:30]
  wire [3:0] _GEN_461 = {{2'd0}, reg_mstatus_prv}; // @[src/main/scala/rocket/CSR.scala 959:40]
  wire [3:0] _cause_T_4 = 4'h8 + _GEN_461; // @[src/main/scala/rocket/CSR.scala 959:40]
  wire [63:0] _cause_T_5 = insn_break ? 64'h3 : io_cause; // @[src/main/scala/rocket/CSR.scala 960:14]
  wire [63:0] cause = insn_call ? {{60'd0}, _cause_T_4} : _cause_T_5; // @[src/main/scala/rocket/CSR.scala 959:8]
  wire [7:0] cause_lsbs = cause[7:0]; // @[src/main/scala/rocket/CSR.scala 961:25]
  wire  _causeIsDebugInt_T_1 = cause_lsbs == 8'he; // @[src/main/scala/rocket/CSR.scala 962:53]
  wire  causeIsDebugInt = cause[63] & cause_lsbs == 8'he; // @[src/main/scala/rocket/CSR.scala 962:39]
  wire  _causeIsDebugTrigger_T_1 = ~cause[63]; // @[src/main/scala/rocket/CSR.scala 963:29]
  wire  causeIsDebugTrigger = ~cause[63] & _causeIsDebugInt_T_1; // @[src/main/scala/rocket/CSR.scala 963:44]
  reg  reg_dcsr_ebreakm; // @[src/main/scala/rocket/CSR.scala 409:25]
  reg  reg_dcsr_ebreaks; // @[src/main/scala/rocket/CSR.scala 409:25]
  reg  reg_dcsr_ebreaku; // @[src/main/scala/rocket/CSR.scala 409:25]
  wire [3:0] _causeIsDebugBreak_T_3 = {reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku}; // @[src/main/scala/rocket/CSR.scala 964:62]
  wire [3:0] _causeIsDebugBreak_T_4 = _causeIsDebugBreak_T_3 >> reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 964:134]
  wire  causeIsDebugBreak = _causeIsDebugTrigger_T_1 & insn_break & _causeIsDebugBreak_T_4[0]; // @[src/main/scala/rocket/CSR.scala 964:56]
  reg  reg_debug; // @[src/main/scala/rocket/CSR.scala 488:26]
  wire  trapToDebug = reg_singleStepped | causeIsDebugInt | causeIsDebugTrigger | causeIsDebugBreak | reg_debug; // @[src/main/scala/rocket/CSR.scala 965:119]
  wire  _T_244 = ~reg_debug; // @[src/main/scala/rocket/CSR.scala 1036:13]
  wire [1:0] _GEN_96 = ~reg_debug ? 2'h3 : reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 1036:25 1043:17 403:28]
  wire  _delegate_T = reg_mstatus_prv <= 2'h1; // @[src/main/scala/rocket/CSR.scala 969:55]
  reg [63:0] reg_mideleg; // @[src/main/scala/rocket/CSR.scala 503:18]
  wire [63:0] read_mideleg = reg_mideleg & 64'h222; // @[src/main/scala/rocket/CSR.scala 504:38]
  wire [63:0] _delegate_T_3 = read_mideleg >> cause_lsbs; // @[src/main/scala/rocket/CSR.scala 969:100]
  reg [63:0] reg_medeleg; // @[src/main/scala/rocket/CSR.scala 507:18]
  wire [63:0] read_medeleg = reg_medeleg & 64'hb15d; // @[src/main/scala/rocket/CSR.scala 508:38]
  wire [63:0] _delegate_T_5 = read_medeleg >> cause_lsbs; // @[src/main/scala/rocket/CSR.scala 969:126]
  wire  _delegate_T_7 = cause[63] ? _delegate_T_3[0] : _delegate_T_5[0]; // @[src/main/scala/rocket/CSR.scala 969:72]
  wire  delegate = reg_mstatus_prv <= 2'h1 & _delegate_T_7; // @[src/main/scala/rocket/CSR.scala 969:66]
  wire [1:0] _GEN_115 = delegate ? 2'h1 : 2'h3; // @[src/main/scala/rocket/CSR.scala 1064:35 1076:15 1088:15]
  wire [1:0] _GEN_190 = trapToDebug ? _GEN_96 : _GEN_115; // @[src/main/scala/rocket/CSR.scala 1035:24]
  wire [1:0] _GEN_227 = exception ? _GEN_190 : reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 1034:20 403:28]
  wire [1:0] new_prv = insn_ret ? ret_prv : _GEN_227; // @[src/main/scala/rocket/CSR.scala 1112:19 1151:13]
  reg [2:0] reg_dcsr_cause; // @[src/main/scala/rocket/CSR.scala 409:25]
  reg  reg_dcsr_step; // @[src/main/scala/rocket/CSR.scala 409:25]
  reg [39:0] reg_dpc; // @[src/main/scala/rocket/CSR.scala 489:20]
  reg [63:0] reg_dscratch0; // @[src/main/scala/rocket/CSR.scala 490:26]
  reg [63:0] reg_mie; // @[src/main/scala/rocket/CSR.scala 501:20]
  reg  reg_mip_seip; // @[src/main/scala/rocket/CSR.scala 510:20]
  reg  reg_mip_stip; // @[src/main/scala/rocket/CSR.scala 510:20]
  reg  reg_mip_ssip; // @[src/main/scala/rocket/CSR.scala 510:20]
  reg [39:0] reg_mepc; // @[src/main/scala/rocket/CSR.scala 511:21]
  reg [63:0] reg_mcause; // @[src/main/scala/rocket/CSR.scala 512:27]
  reg [39:0] reg_mtval; // @[src/main/scala/rocket/CSR.scala 513:22]
  reg [63:0] reg_mscratch; // @[src/main/scala/rocket/CSR.scala 515:25]
  reg [31:0] reg_mtvec; // @[src/main/scala/rocket/CSR.scala 518:31]
  reg [31:0] reg_mcounteren; // @[src/main/scala/rocket/CSR.scala 537:22]
  wire [31:0] read_mcounteren = reg_mcounteren & 32'h7; // @[src/main/scala/rocket/CSR.scala 538:32]
  reg [31:0] reg_scounteren; // @[src/main/scala/rocket/CSR.scala 541:22]
  wire [31:0] read_scounteren = reg_scounteren & 32'h7; // @[src/main/scala/rocket/CSR.scala 542:38]
  wire [15:0] _read_hvip_T = {4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0}; // @[src/main/scala/rocket/CSR.scala 561:27]
  reg [39:0] reg_sepc; // @[src/main/scala/rocket/CSR.scala 575:21]
  reg [63:0] reg_scause; // @[src/main/scala/rocket/CSR.scala 576:23]
  reg [39:0] reg_stval; // @[src/main/scala/rocket/CSR.scala 577:22]
  reg [63:0] reg_sscratch; // @[src/main/scala/rocket/CSR.scala 578:25]
  reg [38:0] reg_stvec; // @[src/main/scala/rocket/CSR.scala 579:22]
  reg [3:0] reg_satp_mode; // @[src/main/scala/rocket/CSR.scala 580:21]
  reg [43:0] reg_satp_ppn; // @[src/main/scala/rocket/CSR.scala 580:21]
  reg  reg_wfi; // @[src/main/scala/rocket/CSR.scala 581:54]
  reg [5:0] small_; // @[src/main/scala/util/Counters.scala 45:41]
  wire [5:0] _GEN_462 = {{5'd0}, io_retire}; // @[src/main/scala/util/Counters.scala 46:33]
  wire [6:0] nextSmall = small_ + _GEN_462; // @[src/main/scala/util/Counters.scala 46:33]
  reg [57:0] large_; // @[src/main/scala/util/Counters.scala 50:31]
  wire  line_1041_clock;
  wire  line_1041_reset;
  wire  line_1041_valid;
  reg  line_1041_valid_reg;
  wire [57:0] _large_r_T_1 = large_ + 58'h1; // @[src/main/scala/util/Counters.scala 51:55]
  wire [57:0] _GEN_80 = nextSmall[6] ? _large_r_T_1 : large_; // @[src/main/scala/util/Counters.scala 50:31 51:{46,50}]
  wire [63:0] value = {large_,small_}; // @[src/main/scala/util/Counters.scala 55:30]
  wire  x10 = ~io_csr_stall; // @[src/main/scala/rocket/CSR.scala 594:56]
  reg [5:0] small_1; // @[src/main/scala/util/Counters.scala 45:41]
  wire [5:0] _GEN_463 = {{5'd0}, x10}; // @[src/main/scala/util/Counters.scala 46:33]
  wire [6:0] nextSmall_1 = small_1 + _GEN_463; // @[src/main/scala/util/Counters.scala 46:33]
  reg [57:0] large_1; // @[src/main/scala/util/Counters.scala 50:31]
  wire  line_1042_clock;
  wire  line_1042_reset;
  wire  line_1042_valid;
  reg  line_1042_valid_reg;
  wire [57:0] _large_r_T_3 = large_1 + 58'h1; // @[src/main/scala/util/Counters.scala 51:55]
  wire [57:0] _GEN_82 = nextSmall_1[6] ? _large_r_T_3 : large_1; // @[src/main/scala/util/Counters.scala 50:31 51:{46,50}]
  wire [63:0] value_1 = {large_1,small_1}; // @[src/main/scala/util/Counters.scala 55:30]
  wire [15:0] read_mip = _read_hvip_T & 16'haaa; // @[src/main/scala/rocket/CSR.scala 610:29]
  wire [63:0] _GEN_464 = {{48'd0}, read_mip}; // @[src/main/scala/rocket/CSR.scala 614:56]
  wire [63:0] pending_interrupts = _GEN_464 & reg_mie; // @[src/main/scala/rocket/CSR.scala 614:56]
  wire [63:0] _m_interrupts_T_3 = ~pending_interrupts; // @[src/main/scala/rocket/CSR.scala 620:85]
  wire [63:0] _m_interrupts_T_4 = _m_interrupts_T_3 | read_mideleg; // @[src/main/scala/rocket/CSR.scala 620:105]
  wire [63:0] _m_interrupts_T_5 = ~_m_interrupts_T_4; // @[src/main/scala/rocket/CSR.scala 620:83]
  wire [63:0] m_interrupts = _delegate_T | reg_mstatus_mie ? _m_interrupts_T_5 : 64'h0; // @[src/main/scala/rocket/CSR.scala 620:25]
  wire [63:0] _s_interrupts_T_6 = pending_interrupts & read_mideleg; // @[src/main/scala/rocket/CSR.scala 621:151]
  wire [63:0] s_interrupts = reg_mstatus_prv < 2'h1 | reg_mstatus_prv == 2'h1 & reg_mstatus_sie ? _s_interrupts_T_6 : 64'h0
    ; // @[src/main/scala/rocket/CSR.scala 621:25]
  wire  _any_T_93 = m_interrupts[15] | m_interrupts[14] | m_interrupts[13] | m_interrupts[12] | m_interrupts[11] |
    m_interrupts[3] | m_interrupts[7] | m_interrupts[9] | m_interrupts[1] | m_interrupts[5] | m_interrupts[10] |
    m_interrupts[2] | m_interrupts[6] | m_interrupts[8] | m_interrupts[0] | m_interrupts[4]; // @[src/main/scala/rocket/CSR.scala 1689:90]
  wire  _any_T_108 = _any_T_93 | s_interrupts[15] | s_interrupts[14] | s_interrupts[13] | s_interrupts[12] |
    s_interrupts[11] | s_interrupts[3] | s_interrupts[7] | s_interrupts[9] | s_interrupts[1] | s_interrupts[5] |
    s_interrupts[10] | s_interrupts[2] | s_interrupts[6] | s_interrupts[8] | s_interrupts[0]; // @[src/main/scala/rocket/CSR.scala 1689:90]
  wire  anyInterrupt = _any_T_108 | s_interrupts[4]; // @[src/main/scala/rocket/CSR.scala 1689:90]
  wire [3:0] _which_T_79 = s_interrupts[0] ? 4'h0 : 4'h4; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_80 = s_interrupts[8] ? 4'h8 : _which_T_79; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_81 = s_interrupts[6] ? 4'h6 : _which_T_80; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_82 = s_interrupts[2] ? 4'h2 : _which_T_81; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_83 = s_interrupts[10] ? 4'ha : _which_T_82; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_84 = s_interrupts[5] ? 4'h5 : _which_T_83; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_85 = s_interrupts[1] ? 4'h1 : _which_T_84; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_86 = s_interrupts[9] ? 4'h9 : _which_T_85; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_87 = s_interrupts[7] ? 4'h7 : _which_T_86; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_88 = s_interrupts[3] ? 4'h3 : _which_T_87; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_89 = s_interrupts[11] ? 4'hb : _which_T_88; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_90 = s_interrupts[12] ? 4'hc : _which_T_89; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_91 = s_interrupts[13] ? 4'hd : _which_T_90; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_92 = s_interrupts[14] ? 4'he : _which_T_91; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_93 = s_interrupts[15] ? 4'hf : _which_T_92; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_94 = m_interrupts[4] ? 4'h4 : _which_T_93; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_95 = m_interrupts[0] ? 4'h0 : _which_T_94; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_96 = m_interrupts[8] ? 4'h8 : _which_T_95; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_97 = m_interrupts[6] ? 4'h6 : _which_T_96; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_98 = m_interrupts[2] ? 4'h2 : _which_T_97; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_99 = m_interrupts[10] ? 4'ha : _which_T_98; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_100 = m_interrupts[5] ? 4'h5 : _which_T_99; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_101 = m_interrupts[1] ? 4'h1 : _which_T_100; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_102 = m_interrupts[9] ? 4'h9 : _which_T_101; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_103 = m_interrupts[7] ? 4'h7 : _which_T_102; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_104 = m_interrupts[3] ? 4'h3 : _which_T_103; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_105 = m_interrupts[11] ? 4'hb : _which_T_104; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_106 = m_interrupts[12] ? 4'hc : _which_T_105; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_107 = m_interrupts[13] ? 4'hd : _which_T_106; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _which_T_108 = m_interrupts[14] ? 4'he : _which_T_107; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] whichInterrupt = m_interrupts[15] ? 4'hf : _which_T_108; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [63:0] _GEN_465 = {{60'd0}, whichInterrupt}; // @[src/main/scala/rocket/CSR.scala 625:63]
  wire  _io_interrupt_T = ~io_singleStep; // @[src/main/scala/rocket/CSR.scala 626:36]
  reg [63:0] reg_misa; // @[src/main/scala/rocket/CSR.scala 650:25]
  wire [8:0] read_mstatus_lo_lo = {io_status_spp,io_status_mpie,io_status_ube,io_status_spie,io_status_upie,
    io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[src/main/scala/rocket/CSR.scala 651:32]
  wire [21:0] read_mstatus_lo = {io_status_tw,io_status_tvm,io_status_mxr,io_status_sum,io_status_mprv,io_status_xs,
    io_status_fs,io_status_mpp,io_status_vs,read_mstatus_lo_lo}; // @[src/main/scala/rocket/CSR.scala 651:32]
  wire [64:0] read_mstatus_hi_hi = {io_status_debug,io_status_cease,io_status_wfi,io_status_isa,io_status_dprv,
    io_status_dv,io_status_prv,io_status_v,io_status_sd,io_status_zero2}; // @[src/main/scala/rocket/CSR.scala 651:32]
  wire [82:0] read_mstatus_hi = {read_mstatus_hi_hi,io_status_mpv,io_status_gva,io_status_mbe,io_status_sbe,
    io_status_sxl,io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr}; // @[src/main/scala/rocket/CSR.scala 651:32]
  wire [104:0] _read_mstatus_T = {read_mstatus_hi,read_mstatus_lo}; // @[src/main/scala/rocket/CSR.scala 651:32]
  wire [63:0] read_mstatus = _read_mstatus_T[63:0]; // @[src/main/scala/util/package.scala 155:13]
  wire [7:0] _read_mtvec_T_1 = reg_mtvec[0] ? 8'hfe : 8'h2; // @[src/main/scala/rocket/CSR.scala 1718:39]
  wire [31:0] _read_mtvec_T_3 = {{24'd0}, _read_mtvec_T_1}; // @[src/main/scala/util/package.scala 166:41]
  wire [31:0] _read_mtvec_T_4 = ~_read_mtvec_T_3; // @[src/main/scala/util/package.scala 166:37]
  wire [31:0] _read_mtvec_T_5 = reg_mtvec & _read_mtvec_T_4; // @[src/main/scala/util/package.scala 166:35]
  wire [63:0] read_mtvec = {32'h0,_read_mtvec_T_5}; // @[src/main/scala/util/package.scala 130:15]
  wire [7:0] _read_stvec_T_1 = reg_stvec[0] ? 8'hfe : 8'h2; // @[src/main/scala/rocket/CSR.scala 1718:39]
  wire [38:0] _read_stvec_T_3 = {{31'd0}, _read_stvec_T_1}; // @[src/main/scala/util/package.scala 166:41]
  wire [38:0] _read_stvec_T_4 = ~_read_stvec_T_3; // @[src/main/scala/util/package.scala 166:37]
  wire [38:0] _read_stvec_T_5 = reg_stvec & _read_stvec_T_4; // @[src/main/scala/util/package.scala 166:35]
  wire [24:0] _read_stvec_T_7 = _read_stvec_T_5[38] ? 25'h1ffffff : 25'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] read_stvec = {_read_stvec_T_7,_read_stvec_T_5}; // @[src/main/scala/util/package.scala 124:15]
  wire [39:0] _T_19 = ~reg_mepc; // @[src/main/scala/rocket/CSR.scala 1717:28]
  wire [1:0] _T_21 = reg_misa[2] ? 2'h1 : 2'h3; // @[src/main/scala/rocket/CSR.scala 1717:36]
  wire [39:0] _GEN_466 = {{38'd0}, _T_21}; // @[src/main/scala/rocket/CSR.scala 1717:31]
  wire [39:0] _T_22 = _T_19 | _GEN_466; // @[src/main/scala/rocket/CSR.scala 1717:31]
  wire [39:0] _T_23 = ~_T_22; // @[src/main/scala/rocket/CSR.scala 1717:26]
  wire [23:0] _T_25 = _T_23[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] _T_26 = {_T_25,_T_23}; // @[src/main/scala/util/package.scala 124:15]
  wire [23:0] _T_28 = reg_mtval[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] _T_29 = {_T_28,reg_mtval}; // @[src/main/scala/util/package.scala 124:15]
  wire [10:0] lo_4 = {2'h0,reg_dcsr_cause,1'h0,2'h0,reg_dcsr_step,reg_dcsr_prv}; // @[src/main/scala/rocket/CSR.scala 668:27]
  wire [31:0] _T_30 = {4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,1'h0,lo_4}; // @[src/main/scala/rocket/CSR.scala 668:27]
  wire [39:0] _T_31 = ~reg_dpc; // @[src/main/scala/rocket/CSR.scala 1717:28]
  wire [39:0] _T_34 = _T_31 | _GEN_466; // @[src/main/scala/rocket/CSR.scala 1717:31]
  wire [39:0] _T_35 = ~_T_34; // @[src/main/scala/rocket/CSR.scala 1717:26]
  wire [23:0] _T_37 = _T_35[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] _T_38 = {_T_37,_T_35}; // @[src/main/scala/util/package.scala 124:15]
  wire [63:0] sie_mask = read_mideleg & 64'hefff; // @[src/main/scala/rocket/CSR.scala 756:18]
  wire [63:0] read_sie = reg_mie & sie_mask; // @[src/main/scala/rocket/CSR.scala 760:28]
  wire [63:0] read_sip = _GEN_464 & sie_mask; // @[src/main/scala/rocket/CSR.scala 761:29]
  wire [8:0] sstatus_lo_lo = {io_status_spp,1'h0,1'h0,io_status_spie,1'h0,2'h0,io_status_sie,1'h0}; // @[src/main/scala/rocket/CSR.scala 774:37]
  wire [21:0] sstatus_lo = {2'h0,io_status_mxr,io_status_sum,1'h0,io_status_xs,io_status_fs,2'h0,io_status_vs,
    sstatus_lo_lo}; // @[src/main/scala/rocket/CSR.scala 774:37]
  wire [104:0] _sstatus_T = {37'h0,4'h0,io_status_sd,23'h0,6'h0,io_status_uxl,io_status_sd_rv32,9'h0,sstatus_lo}; // @[src/main/scala/rocket/CSR.scala 774:37]
  wire [23:0] _T_43 = reg_stval[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] _T_44 = {_T_43,reg_stval}; // @[src/main/scala/util/package.scala 124:15]
  wire [19:0] hi_7 = {reg_satp_mode,16'h0}; // @[src/main/scala/rocket/CSR.scala 782:43]
  wire [63:0] _T_45 = {reg_satp_mode,16'h0,reg_satp_ppn}; // @[src/main/scala/rocket/CSR.scala 782:43]
  wire [39:0] _T_46 = ~reg_sepc; // @[src/main/scala/rocket/CSR.scala 1717:28]
  wire [39:0] _T_49 = _T_46 | _GEN_466; // @[src/main/scala/rocket/CSR.scala 1717:31]
  wire [39:0] _T_50 = ~_T_49; // @[src/main/scala/rocket/CSR.scala 1717:26]
  wire [23:0] _T_52 = _T_50[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire [63:0] _T_53 = {_T_52,_T_50}; // @[src/main/scala/util/package.scala 124:15]
  wire [12:0] addr = {io_status_v,io_rw_addr}; // @[src/main/scala/rocket/CSR.scala 859:19]
  wire [11:0] decoded_decoded_plaInput = addr[11:0]; // @[src/main/scala/chisel3/util/experimental/decode/decoder.scala 39:16 src/main/scala/chisel3/util/pla.scala 77:22]
  wire [11:0] decoded_decoded_invInputs = ~decoded_decoded_plaInput; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  decoded_decoded_andMatrixInput_0 = decoded_decoded_invInputs[2]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_1 = decoded_decoded_invInputs[3]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_2 = decoded_decoded_invInputs[4]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_3 = decoded_decoded_invInputs[5]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_4 = decoded_decoded_invInputs[6]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_5 = decoded_decoded_invInputs[7]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_6 = decoded_decoded_plaInput[8]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_decoded_andMatrixInput_7 = decoded_decoded_invInputs[9]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_8 = decoded_decoded_invInputs[10]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_9 = decoded_decoded_invInputs[11]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [4:0] decoded_decoded_lo = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [9:0] _decoded_decoded_T = {decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,
    decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_1 = &_decoded_decoded_T; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_0_1 = decoded_decoded_invInputs[0]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_1_1 = decoded_decoded_invInputs[1]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_decoded_andMatrixInput_2_1 = decoded_decoded_plaInput[2]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] decoded_decoded_lo_1 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_2 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_3 = &_decoded_decoded_T_2; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_0_2 = decoded_decoded_plaInput[0]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [11:0] _decoded_decoded_T_4 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_5 = &_decoded_decoded_T_4; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_0_3 = decoded_decoded_plaInput[1]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [10:0] _decoded_decoded_T_6 = {decoded_decoded_andMatrixInput_0_3,decoded_decoded_andMatrixInput_2_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_7 = &_decoded_decoded_T_6; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_0_4 = decoded_decoded_plaInput[3]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [8:0] _decoded_decoded_T_8 = {decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_9 = &_decoded_decoded_T_8; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_6_5 = decoded_decoded_plaInput[6]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] decoded_decoded_lo_5 = {decoded_decoded_andMatrixInput_6_5,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_10 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_11 = &_decoded_decoded_T_10; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_12 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_13 = &_decoded_decoded_T_12; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_14 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_15 = &_decoded_decoded_T_14; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_16 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_17 = &_decoded_decoded_T_16; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [9:0] _decoded_decoded_T_18 = {decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_6_5,
    decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_7,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_19 = &_decoded_decoded_T_18; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_0_10 = decoded_decoded_plaInput[7]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [4:0] _decoded_decoded_T_20 = {decoded_decoded_andMatrixInput_0_10,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_21 = &_decoded_decoded_T_20; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_9_9 = decoded_decoded_plaInput[9]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] decoded_decoded_lo_11 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_22 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_23 = &_decoded_decoded_T_22; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_24 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_25 = &_decoded_decoded_T_24; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_26 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_27 = &_decoded_decoded_T_26; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_28 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_29 = &_decoded_decoded_T_28; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_30 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_31 = &_decoded_decoded_T_30; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_32 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_33 = &_decoded_decoded_T_32; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [4:0] decoded_decoded_lo_17 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _decoded_decoded_T_34 = {decoded_decoded_andMatrixInput_0_3,decoded_decoded_andMatrixInput_2_1,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_17}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_35 = &_decoded_decoded_T_34; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _decoded_decoded_T_36 = {decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_37 = &_decoded_decoded_T_36; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_4_19 = decoded_decoded_plaInput[5]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [10:0] _decoded_decoded_T_38 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_19,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_17}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_39 = &_decoded_decoded_T_38; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [10:0] _decoded_decoded_T_40 = {decoded_decoded_andMatrixInput_0_3,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_4_19,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_17}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_41 = &_decoded_decoded_T_40; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_42 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_43 = &_decoded_decoded_T_42; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_44 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_45 = &_decoded_decoded_T_44; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_46 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_47 = &_decoded_decoded_T_46; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_48 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_49 = &_decoded_decoded_T_48; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_50 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_51 = &_decoded_decoded_T_50; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_52 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_53 = &_decoded_decoded_T_52; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_54 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_55 = &_decoded_decoded_T_54; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_56 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_57 = &_decoded_decoded_T_56; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_58 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_59 = &_decoded_decoded_T_58; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_60 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_61 = &_decoded_decoded_T_60; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_62 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_63 = &_decoded_decoded_T_62; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_64 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_65 = &_decoded_decoded_T_64; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_4_33 = decoded_decoded_plaInput[4]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [11:0] _decoded_decoded_T_66 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_67 = &_decoded_decoded_T_66; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_68 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_69 = &_decoded_decoded_T_68; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_70 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_71 = &_decoded_decoded_T_70; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_72 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_73 = &_decoded_decoded_T_72; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_74 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_75 = &_decoded_decoded_T_74; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_76 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_77 = &_decoded_decoded_T_76; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_78 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_79 = &_decoded_decoded_T_78; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_80 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_81 = &_decoded_decoded_T_80; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_82 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_83 = &_decoded_decoded_T_82; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_84 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_85 = &_decoded_decoded_T_84; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_86 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_87 = &_decoded_decoded_T_86; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_88 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_89 = &_decoded_decoded_T_88; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_90 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_91 = &_decoded_decoded_T_90; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_92 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_93 = &_decoded_decoded_T_92; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_94 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_95 = &_decoded_decoded_T_94; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_96 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_97 = &_decoded_decoded_T_96; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] decoded_decoded_lo_49 = {decoded_decoded_andMatrixInput_6_5,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_98 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_49}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_99 = &_decoded_decoded_T_98; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_100 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_49}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_101 = &_decoded_decoded_T_100; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_102 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_49}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_103 = &_decoded_decoded_T_102; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_104 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_49}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_105 = &_decoded_decoded_T_104; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [9:0] _decoded_decoded_T_106 = {decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,
    decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,decoded_decoded_andMatrixInput_6_5,
    decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,
    decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_107 = &_decoded_decoded_T_106; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_10_48 = decoded_decoded_plaInput[10]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] decoded_decoded_lo_54 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_0_10,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_10_48,
    decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_108 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_54}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_109 = &_decoded_decoded_T_108; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_110 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_4_19,decoded_decoded_lo_54}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_111 = &_decoded_decoded_T_110; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [4:0] decoded_decoded_lo_56 = {decoded_decoded_andMatrixInput_0_10,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_10_48,decoded_decoded_andMatrixInput_9}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _decoded_decoded_T_112 = {decoded_decoded_andMatrixInput_0_3,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,decoded_decoded_andMatrixInput_4_19,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_56}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_113 = &_decoded_decoded_T_112; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_10_51 = decoded_decoded_plaInput[11]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [4:0] decoded_decoded_lo_57 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _decoded_decoded_T_114 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_57}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_115 = &_decoded_decoded_T_114; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] decoded_decoded_lo_58 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_8,
    decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_116 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_117 = &_decoded_decoded_T_116; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_118 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_119 = &_decoded_decoded_T_118; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_120 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_121 = &_decoded_decoded_T_120; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_122 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_123 = &_decoded_decoded_T_122; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_124 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_125 = &_decoded_decoded_T_124; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_126 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_127 = &_decoded_decoded_T_126; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_128 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_129 = &_decoded_decoded_T_128; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_130 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_131 = &_decoded_decoded_T_130; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_132 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_133 = &_decoded_decoded_T_132; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_134 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_135 = &_decoded_decoded_T_134; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_136 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_137 = &_decoded_decoded_T_136; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_138 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_139 = &_decoded_decoded_T_138; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_140 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_141 = &_decoded_decoded_T_140; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_142 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_143 = &_decoded_decoded_T_142; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_144 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_145 = &_decoded_decoded_T_144; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_146 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_147 = &_decoded_decoded_T_146; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_148 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_149 = &_decoded_decoded_T_148; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_150 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_151 = &_decoded_decoded_T_150; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_152 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_153 = &_decoded_decoded_T_152; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_154 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_155 = &_decoded_decoded_T_154; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_156 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_157 = &_decoded_decoded_T_156; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_158 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_159 = &_decoded_decoded_T_158; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_160 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_161 = &_decoded_decoded_T_160; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_162 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_163 = &_decoded_decoded_T_162; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_164 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_165 = &_decoded_decoded_T_164; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_166 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_167 = &_decoded_decoded_T_166; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_168 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_169 = &_decoded_decoded_T_168; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_170 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_171 = &_decoded_decoded_T_170; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_172 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_173 = &_decoded_decoded_T_172; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_174 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_58}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_175 = &_decoded_decoded_T_174; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_decoded_andMatrixInput_7_87 = decoded_decoded_invInputs[8]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [4:0] decoded_decoded_lo_88 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_7_87,
    decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_10_48,decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _decoded_decoded_T_176 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_88}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_177 = &_decoded_decoded_T_176; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] decoded_decoded_lo_89 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_7_87,decoded_decoded_andMatrixInput_7,decoded_decoded_andMatrixInput_10_48,
    decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_178 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_179 = &_decoded_decoded_T_178; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_180 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_181 = &_decoded_decoded_T_180; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_182 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_183 = &_decoded_decoded_T_182; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_184 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_185 = &_decoded_decoded_T_184; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_186 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_187 = &_decoded_decoded_T_186; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_188 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_189 = &_decoded_decoded_T_188; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_190 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_191 = &_decoded_decoded_T_190; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_192 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_193 = &_decoded_decoded_T_192; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_194 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_195 = &_decoded_decoded_T_194; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_196 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_197 = &_decoded_decoded_T_196; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_198 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_199 = &_decoded_decoded_T_198; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_200 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_201 = &_decoded_decoded_T_200; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_202 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_203 = &_decoded_decoded_T_202; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_204 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_2,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_205 = &_decoded_decoded_T_204; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_206 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_207 = &_decoded_decoded_T_206; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_208 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_209 = &_decoded_decoded_T_208; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_210 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_211 = &_decoded_decoded_T_210; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_212 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_213 = &_decoded_decoded_T_212; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_214 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_215 = &_decoded_decoded_T_214; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_216 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_217 = &_decoded_decoded_T_216; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_218 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_219 = &_decoded_decoded_T_218; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_220 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_221 = &_decoded_decoded_T_220; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_222 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_223 = &_decoded_decoded_T_222; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_224 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_225 = &_decoded_decoded_T_224; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_226 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_227 = &_decoded_decoded_T_226; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_228 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_229 = &_decoded_decoded_T_228; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_230 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_231 = &_decoded_decoded_T_230; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_232 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_233 = &_decoded_decoded_T_232; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_234 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_235 = &_decoded_decoded_T_234; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_236 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_0_4,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_237 = &_decoded_decoded_T_236; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [4:0] decoded_decoded_lo_119 = {decoded_decoded_andMatrixInput_5,decoded_decoded_andMatrixInput_6,
    decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_10_48,decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _decoded_decoded_T_238 = {decoded_decoded_andMatrixInput_1_1,decoded_decoded_andMatrixInput_0,
    decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,decoded_decoded_andMatrixInput_3,
    decoded_decoded_andMatrixInput_4,decoded_decoded_lo_119}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_239 = &_decoded_decoded_T_238; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] decoded_decoded_lo_120 = {decoded_decoded_andMatrixInput_4,decoded_decoded_andMatrixInput_5,
    decoded_decoded_andMatrixInput_6,decoded_decoded_andMatrixInput_9_9,decoded_decoded_andMatrixInput_10_48,
    decoded_decoded_andMatrixInput_10_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_decoded_T_240 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_120}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_241 = &_decoded_decoded_T_240; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_242 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_0_3,
    decoded_decoded_andMatrixInput_0,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_120}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_243 = &_decoded_decoded_T_242; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_244 = {decoded_decoded_andMatrixInput_0_1,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_120}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_245 = &_decoded_decoded_T_244; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [11:0] _decoded_decoded_T_246 = {decoded_decoded_andMatrixInput_0_2,decoded_decoded_andMatrixInput_1_1,
    decoded_decoded_andMatrixInput_2_1,decoded_decoded_andMatrixInput_1,decoded_decoded_andMatrixInput_4_33,
    decoded_decoded_andMatrixInput_3,decoded_decoded_lo_120}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_decoded_T_247 = &_decoded_decoded_T_246; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_decoded_orMatrixOutputs_T = |_decoded_decoded_T_247; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_1 = |_decoded_decoded_T_243; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_2 = |_decoded_decoded_T_239; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_3 = |_decoded_decoded_T_241; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_4 = |_decoded_decoded_T_9; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_5 = |_decoded_decoded_T_27; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_6 = |_decoded_decoded_T_29; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_7 = |_decoded_decoded_T_7; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_8 = |_decoded_decoded_T_5; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_9 = |_decoded_decoded_T_13; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_10 = |_decoded_decoded_T_21; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_11 = |_decoded_decoded_T_17; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_12 = |_decoded_decoded_T_15; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_13 = |_decoded_decoded_T_11; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_14 = |_decoded_decoded_T_3; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_15 = |_decoded_decoded_T_19; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_16 = |_decoded_decoded_T_1; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_17 = |_decoded_decoded_T_37; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_18 = |_decoded_decoded_T_179; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_19 = |_decoded_decoded_T_177; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_20 = |_decoded_decoded_T_35; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_21 = |_decoded_decoded_T_237; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_22 = |_decoded_decoded_T_175; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_23 = |_decoded_decoded_T_97; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_24 = |_decoded_decoded_T_235; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_25 = |_decoded_decoded_T_173; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_26 = |_decoded_decoded_T_95; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_27 = |_decoded_decoded_T_233; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_28 = |_decoded_decoded_T_171; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_29 = |_decoded_decoded_T_93; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_30 = |_decoded_decoded_T_231; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_31 = |_decoded_decoded_T_169; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_32 = |_decoded_decoded_T_91; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_33 = |_decoded_decoded_T_229; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_34 = |_decoded_decoded_T_167; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_35 = |_decoded_decoded_T_89; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_36 = |_decoded_decoded_T_227; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_37 = |_decoded_decoded_T_165; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_38 = |_decoded_decoded_T_87; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_39 = |_decoded_decoded_T_225; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_40 = |_decoded_decoded_T_163; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_41 = |_decoded_decoded_T_85; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_42 = |_decoded_decoded_T_223; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_43 = |_decoded_decoded_T_161; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_44 = |_decoded_decoded_T_83; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_45 = |_decoded_decoded_T_221; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_46 = |_decoded_decoded_T_159; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_47 = |_decoded_decoded_T_81; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_48 = |_decoded_decoded_T_219; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_49 = |_decoded_decoded_T_157; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_50 = |_decoded_decoded_T_79; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_51 = |_decoded_decoded_T_217; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_52 = |_decoded_decoded_T_155; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_53 = |_decoded_decoded_T_77; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_54 = |_decoded_decoded_T_215; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_55 = |_decoded_decoded_T_153; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_56 = |_decoded_decoded_T_75; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_57 = |_decoded_decoded_T_213; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_58 = |_decoded_decoded_T_151; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_59 = |_decoded_decoded_T_73; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_60 = |_decoded_decoded_T_211; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_61 = |_decoded_decoded_T_149; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_62 = |_decoded_decoded_T_71; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_63 = |_decoded_decoded_T_209; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_64 = |_decoded_decoded_T_147; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_65 = |_decoded_decoded_T_69; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_66 = |_decoded_decoded_T_207; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_67 = |_decoded_decoded_T_145; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_68 = |_decoded_decoded_T_67; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_69 = |_decoded_decoded_T_205; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_70 = |_decoded_decoded_T_143; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_71 = |_decoded_decoded_T_65; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_72 = |_decoded_decoded_T_203; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_73 = |_decoded_decoded_T_141; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_74 = |_decoded_decoded_T_63; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_75 = |_decoded_decoded_T_201; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_76 = |_decoded_decoded_T_139; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_77 = |_decoded_decoded_T_61; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_78 = |_decoded_decoded_T_199; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_79 = |_decoded_decoded_T_137; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_80 = |_decoded_decoded_T_59; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_81 = |_decoded_decoded_T_197; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_82 = |_decoded_decoded_T_135; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_83 = |_decoded_decoded_T_57; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_84 = |_decoded_decoded_T_195; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_85 = |_decoded_decoded_T_133; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_86 = |_decoded_decoded_T_55; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_87 = |_decoded_decoded_T_193; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_88 = |_decoded_decoded_T_131; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_89 = |_decoded_decoded_T_53; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_90 = |_decoded_decoded_T_191; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_91 = |_decoded_decoded_T_129; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_92 = |_decoded_decoded_T_51; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_93 = |_decoded_decoded_T_189; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_94 = |_decoded_decoded_T_127; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_95 = |_decoded_decoded_T_49; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_96 = |_decoded_decoded_T_187; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_97 = |_decoded_decoded_T_125; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_98 = |_decoded_decoded_T_47; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_99 = |_decoded_decoded_T_185; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_100 = |_decoded_decoded_T_123; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_101 = |_decoded_decoded_T_45; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_102 = |_decoded_decoded_T_183; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_103 = |_decoded_decoded_T_121; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_104 = |_decoded_decoded_T_43; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_105 = |_decoded_decoded_T_181; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_106 = |_decoded_decoded_T_119; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_107 = |_decoded_decoded_T_41; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_108 = |_decoded_decoded_T_117; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_109 = |_decoded_decoded_T_115; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_110 = |_decoded_decoded_T_39; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_111 = |_decoded_decoded_T_113; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_112 = |_decoded_decoded_T_111; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_113 = |_decoded_decoded_T_109; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_114 = |_decoded_decoded_T_245; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_115 = |_decoded_decoded_T_103; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_116 = |_decoded_decoded_T_105; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_117 = |_decoded_decoded_T_101; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_118 = |_decoded_decoded_T_99; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_119 = |_decoded_decoded_T_31; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_120 = |_decoded_decoded_T_107; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_121 = |_decoded_decoded_T_33; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_122 = |_decoded_decoded_T_23; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_decoded_orMatrixOutputs_T_123 = |_decoded_decoded_T_25; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_6,
    _decoded_decoded_orMatrixOutputs_T_5,_decoded_decoded_orMatrixOutputs_T_4,_decoded_decoded_orMatrixOutputs_T_3,
    _decoded_decoded_orMatrixOutputs_T_2,_decoded_decoded_orMatrixOutputs_T_1,_decoded_decoded_orMatrixOutputs_T}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [14:0] decoded_decoded_orMatrixOutputs_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_14,
    _decoded_decoded_orMatrixOutputs_T_13,_decoded_decoded_orMatrixOutputs_T_12,_decoded_decoded_orMatrixOutputs_T_11,
    _decoded_decoded_orMatrixOutputs_T_10,_decoded_decoded_orMatrixOutputs_T_9,_decoded_decoded_orMatrixOutputs_T_8,
    _decoded_decoded_orMatrixOutputs_T_7,decoded_decoded_orMatrixOutputs_lo_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [7:0] decoded_decoded_orMatrixOutputs_lo_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_22,
    _decoded_decoded_orMatrixOutputs_T_21,_decoded_decoded_orMatrixOutputs_T_20,_decoded_decoded_orMatrixOutputs_T_19,
    _decoded_decoded_orMatrixOutputs_T_18,_decoded_decoded_orMatrixOutputs_T_17,_decoded_decoded_orMatrixOutputs_T_16,
    _decoded_decoded_orMatrixOutputs_T_15}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [30:0] decoded_decoded_orMatrixOutputs_lo_lo = {_decoded_decoded_orMatrixOutputs_T_30,
    _decoded_decoded_orMatrixOutputs_T_29,_decoded_decoded_orMatrixOutputs_T_28,_decoded_decoded_orMatrixOutputs_T_27,
    _decoded_decoded_orMatrixOutputs_T_26,_decoded_decoded_orMatrixOutputs_T_25,_decoded_decoded_orMatrixOutputs_T_24,
    _decoded_decoded_orMatrixOutputs_T_23,decoded_decoded_orMatrixOutputs_lo_lo_hi_lo,
    decoded_decoded_orMatrixOutputs_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [6:0] decoded_decoded_orMatrixOutputs_lo_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_37,
    _decoded_decoded_orMatrixOutputs_T_36,_decoded_decoded_orMatrixOutputs_T_35,_decoded_decoded_orMatrixOutputs_T_34,
    _decoded_decoded_orMatrixOutputs_T_33,_decoded_decoded_orMatrixOutputs_T_32,_decoded_decoded_orMatrixOutputs_T_31}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [14:0] decoded_decoded_orMatrixOutputs_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_45,
    _decoded_decoded_orMatrixOutputs_T_44,_decoded_decoded_orMatrixOutputs_T_43,_decoded_decoded_orMatrixOutputs_T_42,
    _decoded_decoded_orMatrixOutputs_T_41,_decoded_decoded_orMatrixOutputs_T_40,_decoded_decoded_orMatrixOutputs_T_39,
    _decoded_decoded_orMatrixOutputs_T_38,decoded_decoded_orMatrixOutputs_lo_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [7:0] decoded_decoded_orMatrixOutputs_lo_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_53,
    _decoded_decoded_orMatrixOutputs_T_52,_decoded_decoded_orMatrixOutputs_T_51,_decoded_decoded_orMatrixOutputs_T_50,
    _decoded_decoded_orMatrixOutputs_T_49,_decoded_decoded_orMatrixOutputs_T_48,_decoded_decoded_orMatrixOutputs_T_47,
    _decoded_decoded_orMatrixOutputs_T_46}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [30:0] decoded_decoded_orMatrixOutputs_lo_hi = {_decoded_decoded_orMatrixOutputs_T_61,
    _decoded_decoded_orMatrixOutputs_T_60,_decoded_decoded_orMatrixOutputs_T_59,_decoded_decoded_orMatrixOutputs_T_58,
    _decoded_decoded_orMatrixOutputs_T_57,_decoded_decoded_orMatrixOutputs_T_56,_decoded_decoded_orMatrixOutputs_T_55,
    _decoded_decoded_orMatrixOutputs_T_54,decoded_decoded_orMatrixOutputs_lo_hi_hi_lo,
    decoded_decoded_orMatrixOutputs_lo_hi_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [6:0] decoded_decoded_orMatrixOutputs_hi_lo_lo_lo = {_decoded_decoded_orMatrixOutputs_T_68,
    _decoded_decoded_orMatrixOutputs_T_67,_decoded_decoded_orMatrixOutputs_T_66,_decoded_decoded_orMatrixOutputs_T_65,
    _decoded_decoded_orMatrixOutputs_T_64,_decoded_decoded_orMatrixOutputs_T_63,_decoded_decoded_orMatrixOutputs_T_62}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [14:0] decoded_decoded_orMatrixOutputs_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_76,
    _decoded_decoded_orMatrixOutputs_T_75,_decoded_decoded_orMatrixOutputs_T_74,_decoded_decoded_orMatrixOutputs_T_73,
    _decoded_decoded_orMatrixOutputs_T_72,_decoded_decoded_orMatrixOutputs_T_71,_decoded_decoded_orMatrixOutputs_T_70,
    _decoded_decoded_orMatrixOutputs_T_69,decoded_decoded_orMatrixOutputs_hi_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [7:0] decoded_decoded_orMatrixOutputs_hi_lo_hi_lo = {_decoded_decoded_orMatrixOutputs_T_84,
    _decoded_decoded_orMatrixOutputs_T_83,_decoded_decoded_orMatrixOutputs_T_82,_decoded_decoded_orMatrixOutputs_T_81,
    _decoded_decoded_orMatrixOutputs_T_80,_decoded_decoded_orMatrixOutputs_T_79,_decoded_decoded_orMatrixOutputs_T_78,
    _decoded_decoded_orMatrixOutputs_T_77}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [30:0] decoded_decoded_orMatrixOutputs_hi_lo = {_decoded_decoded_orMatrixOutputs_T_92,
    _decoded_decoded_orMatrixOutputs_T_91,_decoded_decoded_orMatrixOutputs_T_90,_decoded_decoded_orMatrixOutputs_T_89,
    _decoded_decoded_orMatrixOutputs_T_88,_decoded_decoded_orMatrixOutputs_T_87,_decoded_decoded_orMatrixOutputs_T_86,
    _decoded_decoded_orMatrixOutputs_T_85,decoded_decoded_orMatrixOutputs_hi_lo_hi_lo,
    decoded_decoded_orMatrixOutputs_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [6:0] decoded_decoded_orMatrixOutputs_hi_hi_lo_lo = {_decoded_decoded_orMatrixOutputs_T_99,
    _decoded_decoded_orMatrixOutputs_T_98,_decoded_decoded_orMatrixOutputs_T_97,_decoded_decoded_orMatrixOutputs_T_96,
    _decoded_decoded_orMatrixOutputs_T_95,_decoded_decoded_orMatrixOutputs_T_94,_decoded_decoded_orMatrixOutputs_T_93}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [14:0] decoded_decoded_orMatrixOutputs_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_107,
    _decoded_decoded_orMatrixOutputs_T_106,_decoded_decoded_orMatrixOutputs_T_105,_decoded_decoded_orMatrixOutputs_T_104
    ,_decoded_decoded_orMatrixOutputs_T_103,_decoded_decoded_orMatrixOutputs_T_102,
    _decoded_decoded_orMatrixOutputs_T_101,_decoded_decoded_orMatrixOutputs_T_100,
    decoded_decoded_orMatrixOutputs_hi_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [7:0] decoded_decoded_orMatrixOutputs_hi_hi_hi_lo = {_decoded_decoded_orMatrixOutputs_T_115,
    _decoded_decoded_orMatrixOutputs_T_114,_decoded_decoded_orMatrixOutputs_T_113,_decoded_decoded_orMatrixOutputs_T_112
    ,_decoded_decoded_orMatrixOutputs_T_111,_decoded_decoded_orMatrixOutputs_T_110,
    _decoded_decoded_orMatrixOutputs_T_109,_decoded_decoded_orMatrixOutputs_T_108}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [30:0] decoded_decoded_orMatrixOutputs_hi_hi = {_decoded_decoded_orMatrixOutputs_T_123,
    _decoded_decoded_orMatrixOutputs_T_122,_decoded_decoded_orMatrixOutputs_T_121,_decoded_decoded_orMatrixOutputs_T_120
    ,_decoded_decoded_orMatrixOutputs_T_119,_decoded_decoded_orMatrixOutputs_T_118,
    _decoded_decoded_orMatrixOutputs_T_117,_decoded_decoded_orMatrixOutputs_T_116,
    decoded_decoded_orMatrixOutputs_hi_hi_hi_lo,decoded_decoded_orMatrixOutputs_hi_hi_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [123:0] decoded_decoded_orMatrixOutputs = {decoded_decoded_orMatrixOutputs_hi_hi,
    decoded_decoded_orMatrixOutputs_hi_lo,decoded_decoded_orMatrixOutputs_lo_hi,decoded_decoded_orMatrixOutputs_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [6:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_lo = {decoded_decoded_orMatrixOutputs[6],
    decoded_decoded_orMatrixOutputs[5],decoded_decoded_orMatrixOutputs[4],decoded_decoded_orMatrixOutputs[3],
    decoded_decoded_orMatrixOutputs[2],decoded_decoded_orMatrixOutputs[1],decoded_decoded_orMatrixOutputs[0]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [14:0] decoded_decoded_invMatrixOutputs_lo_lo_lo = {decoded_decoded_orMatrixOutputs[14],
    decoded_decoded_orMatrixOutputs[13],decoded_decoded_orMatrixOutputs[12],decoded_decoded_orMatrixOutputs[11],
    decoded_decoded_orMatrixOutputs[10],decoded_decoded_orMatrixOutputs[9],decoded_decoded_orMatrixOutputs[8],
    decoded_decoded_orMatrixOutputs[7],decoded_decoded_invMatrixOutputs_lo_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [7:0] decoded_decoded_invMatrixOutputs_lo_lo_hi_lo = {decoded_decoded_orMatrixOutputs[22],
    decoded_decoded_orMatrixOutputs[21],decoded_decoded_orMatrixOutputs[20],decoded_decoded_orMatrixOutputs[19],
    decoded_decoded_orMatrixOutputs[18],decoded_decoded_orMatrixOutputs[17],decoded_decoded_orMatrixOutputs[16],
    decoded_decoded_orMatrixOutputs[15]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [30:0] decoded_decoded_invMatrixOutputs_lo_lo = {decoded_decoded_orMatrixOutputs[30],
    decoded_decoded_orMatrixOutputs[29],decoded_decoded_orMatrixOutputs[28],decoded_decoded_orMatrixOutputs[27],
    decoded_decoded_orMatrixOutputs[26],decoded_decoded_orMatrixOutputs[25],decoded_decoded_orMatrixOutputs[24],
    decoded_decoded_orMatrixOutputs[23],decoded_decoded_invMatrixOutputs_lo_lo_hi_lo,
    decoded_decoded_invMatrixOutputs_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [6:0] decoded_decoded_invMatrixOutputs_lo_hi_lo_lo = {decoded_decoded_orMatrixOutputs[37],
    decoded_decoded_orMatrixOutputs[36],decoded_decoded_orMatrixOutputs[35],decoded_decoded_orMatrixOutputs[34],
    decoded_decoded_orMatrixOutputs[33],decoded_decoded_orMatrixOutputs[32],decoded_decoded_orMatrixOutputs[31]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [14:0] decoded_decoded_invMatrixOutputs_lo_hi_lo = {decoded_decoded_orMatrixOutputs[45],
    decoded_decoded_orMatrixOutputs[44],decoded_decoded_orMatrixOutputs[43],decoded_decoded_orMatrixOutputs[42],
    decoded_decoded_orMatrixOutputs[41],decoded_decoded_orMatrixOutputs[40],decoded_decoded_orMatrixOutputs[39],
    decoded_decoded_orMatrixOutputs[38],decoded_decoded_invMatrixOutputs_lo_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [7:0] decoded_decoded_invMatrixOutputs_lo_hi_hi_lo = {decoded_decoded_orMatrixOutputs[53],
    decoded_decoded_orMatrixOutputs[52],decoded_decoded_orMatrixOutputs[51],decoded_decoded_orMatrixOutputs[50],
    decoded_decoded_orMatrixOutputs[49],decoded_decoded_orMatrixOutputs[48],decoded_decoded_orMatrixOutputs[47],
    decoded_decoded_orMatrixOutputs[46]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [30:0] decoded_decoded_invMatrixOutputs_lo_hi = {decoded_decoded_orMatrixOutputs[61],
    decoded_decoded_orMatrixOutputs[60],decoded_decoded_orMatrixOutputs[59],decoded_decoded_orMatrixOutputs[58],
    decoded_decoded_orMatrixOutputs[57],decoded_decoded_orMatrixOutputs[56],decoded_decoded_orMatrixOutputs[55],
    decoded_decoded_orMatrixOutputs[54],decoded_decoded_invMatrixOutputs_lo_hi_hi_lo,
    decoded_decoded_invMatrixOutputs_lo_hi_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [6:0] decoded_decoded_invMatrixOutputs_hi_lo_lo_lo = {decoded_decoded_orMatrixOutputs[68],
    decoded_decoded_orMatrixOutputs[67],decoded_decoded_orMatrixOutputs[66],decoded_decoded_orMatrixOutputs[65],
    decoded_decoded_orMatrixOutputs[64],decoded_decoded_orMatrixOutputs[63],decoded_decoded_orMatrixOutputs[62]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [14:0] decoded_decoded_invMatrixOutputs_hi_lo_lo = {decoded_decoded_orMatrixOutputs[76],
    decoded_decoded_orMatrixOutputs[75],decoded_decoded_orMatrixOutputs[74],decoded_decoded_orMatrixOutputs[73],
    decoded_decoded_orMatrixOutputs[72],decoded_decoded_orMatrixOutputs[71],decoded_decoded_orMatrixOutputs[70],
    decoded_decoded_orMatrixOutputs[69],decoded_decoded_invMatrixOutputs_hi_lo_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [7:0] decoded_decoded_invMatrixOutputs_hi_lo_hi_lo = {decoded_decoded_orMatrixOutputs[84],
    decoded_decoded_orMatrixOutputs[83],decoded_decoded_orMatrixOutputs[82],decoded_decoded_orMatrixOutputs[81],
    decoded_decoded_orMatrixOutputs[80],decoded_decoded_orMatrixOutputs[79],decoded_decoded_orMatrixOutputs[78],
    decoded_decoded_orMatrixOutputs[77]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [30:0] decoded_decoded_invMatrixOutputs_hi_lo = {decoded_decoded_orMatrixOutputs[92],
    decoded_decoded_orMatrixOutputs[91],decoded_decoded_orMatrixOutputs[90],decoded_decoded_orMatrixOutputs[89],
    decoded_decoded_orMatrixOutputs[88],decoded_decoded_orMatrixOutputs[87],decoded_decoded_orMatrixOutputs[86],
    decoded_decoded_orMatrixOutputs[85],decoded_decoded_invMatrixOutputs_hi_lo_hi_lo,
    decoded_decoded_invMatrixOutputs_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [6:0] decoded_decoded_invMatrixOutputs_hi_hi_lo_lo = {decoded_decoded_orMatrixOutputs[99],
    decoded_decoded_orMatrixOutputs[98],decoded_decoded_orMatrixOutputs[97],decoded_decoded_orMatrixOutputs[96],
    decoded_decoded_orMatrixOutputs[95],decoded_decoded_orMatrixOutputs[94],decoded_decoded_orMatrixOutputs[93]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [14:0] decoded_decoded_invMatrixOutputs_hi_hi_lo = {decoded_decoded_orMatrixOutputs[107],
    decoded_decoded_orMatrixOutputs[106],decoded_decoded_orMatrixOutputs[105],decoded_decoded_orMatrixOutputs[104],
    decoded_decoded_orMatrixOutputs[103],decoded_decoded_orMatrixOutputs[102],decoded_decoded_orMatrixOutputs[101],
    decoded_decoded_orMatrixOutputs[100],decoded_decoded_invMatrixOutputs_hi_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [7:0] decoded_decoded_invMatrixOutputs_hi_hi_hi_lo = {decoded_decoded_orMatrixOutputs[115],
    decoded_decoded_orMatrixOutputs[114],decoded_decoded_orMatrixOutputs[113],decoded_decoded_orMatrixOutputs[112],
    decoded_decoded_orMatrixOutputs[111],decoded_decoded_orMatrixOutputs[110],decoded_decoded_orMatrixOutputs[109],
    decoded_decoded_orMatrixOutputs[108]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [30:0] decoded_decoded_invMatrixOutputs_hi_hi = {decoded_decoded_orMatrixOutputs[123],
    decoded_decoded_orMatrixOutputs[122],decoded_decoded_orMatrixOutputs[121],decoded_decoded_orMatrixOutputs[120],
    decoded_decoded_orMatrixOutputs[119],decoded_decoded_orMatrixOutputs[118],decoded_decoded_orMatrixOutputs[117],
    decoded_decoded_orMatrixOutputs[116],decoded_decoded_invMatrixOutputs_hi_hi_hi_lo,
    decoded_decoded_invMatrixOutputs_hi_hi_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [123:0] decoded_decoded_invMatrixOutputs = {decoded_decoded_invMatrixOutputs_hi_hi,
    decoded_decoded_invMatrixOutputs_hi_lo,decoded_decoded_invMatrixOutputs_lo_hi,decoded_decoded_invMatrixOutputs_lo_lo
    }; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire  decoded_0 = decoded_decoded_invMatrixOutputs[123]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_1 = decoded_decoded_invMatrixOutputs[122]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_2 = decoded_decoded_invMatrixOutputs[121]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_3 = decoded_decoded_invMatrixOutputs[120]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_4 = decoded_decoded_invMatrixOutputs[119]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_5 = decoded_decoded_invMatrixOutputs[118]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_6 = decoded_decoded_invMatrixOutputs[117]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_7 = decoded_decoded_invMatrixOutputs[116]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_8 = decoded_decoded_invMatrixOutputs[115]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_9 = decoded_decoded_invMatrixOutputs[114]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_10 = decoded_decoded_invMatrixOutputs[113]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_11 = decoded_decoded_invMatrixOutputs[112]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_12 = decoded_decoded_invMatrixOutputs[111]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_14 = decoded_decoded_invMatrixOutputs[109]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_15 = decoded_decoded_invMatrixOutputs[108]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_103 = decoded_decoded_invMatrixOutputs[20]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_104 = decoded_decoded_invMatrixOutputs[19]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_105 = decoded_decoded_invMatrixOutputs[18]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_107 = decoded_decoded_invMatrixOutputs[16]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_108 = decoded_decoded_invMatrixOutputs[15]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_109 = decoded_decoded_invMatrixOutputs[14]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_110 = decoded_decoded_invMatrixOutputs[13]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_111 = decoded_decoded_invMatrixOutputs[12]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_112 = decoded_decoded_invMatrixOutputs[11]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_113 = decoded_decoded_invMatrixOutputs[10]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_114 = decoded_decoded_invMatrixOutputs[9]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_115 = decoded_decoded_invMatrixOutputs[8]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_116 = decoded_decoded_invMatrixOutputs[7]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_117 = decoded_decoded_invMatrixOutputs[6]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_118 = decoded_decoded_invMatrixOutputs[5]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_120 = decoded_decoded_invMatrixOutputs[3]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_121 = decoded_decoded_invMatrixOutputs[2]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  decoded_122 = decoded_decoded_invMatrixOutputs[1]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [63:0] _wdata_T_1 = io_rw_cmd[1] ? io_rw_rdata : 64'h0; // @[src/main/scala/rocket/CSR.scala 1695:9]
  wire [63:0] _wdata_T_2 = _wdata_T_1 | io_rw_wdata; // @[src/main/scala/rocket/CSR.scala 1695:30]
  wire [63:0] _wdata_T_5 = &io_rw_cmd[1:0] ? io_rw_wdata : 64'h0; // @[src/main/scala/rocket/CSR.scala 1695:45]
  wire [63:0] _wdata_T_6 = ~_wdata_T_5; // @[src/main/scala/rocket/CSR.scala 1695:41]
  wire [63:0] wdata = _wdata_T_2 & _wdata_T_6; // @[src/main/scala/rocket/CSR.scala 1695:39]
  wire  insn_cease = system_insn & decoded_invMatrixOutputs[5]; // @[src/main/scala/rocket/CSR.scala 894:83]
  wire  insn_wfi = system_insn & decoded_invMatrixOutputs[4]; // @[src/main/scala/rocket/CSR.scala 894:83]
  wire [11:0] addr_1 = io_decode_0_inst[31:20]; // @[src/main/scala/rocket/CSR.scala 898:27]
  wire [31:0] decoded_invInputs_1 = ~io_decode_0_inst; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  decoded_andMatrixInput_0_7 = decoded_invInputs_1[20]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_1_7 = decoded_invInputs_1[21]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_2_6 = decoded_invInputs_1[22]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_3_6 = decoded_invInputs_1[23]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_4_6 = decoded_invInputs_1[24]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_5_6 = decoded_invInputs_1[25]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_6_6 = decoded_invInputs_1[26]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_7_6 = decoded_invInputs_1[27]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_8_6 = decoded_invInputs_1[28]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_9_6 = decoded_invInputs_1[29]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_10_3 = decoded_invInputs_1[30]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_11_3 = decoded_invInputs_1[31]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [5:0] decoded_lo_6 = {decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_8_6,
    decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _decoded_T_14 = {decoded_andMatrixInput_0_7,decoded_andMatrixInput_1_7,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_lo_6}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_15 = &_decoded_T_14; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_8 = io_decode_0_inst[20]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [11:0] _decoded_T_16 = {decoded_andMatrixInput_0_8,decoded_andMatrixInput_1_7,decoded_andMatrixInput_2_6,
    decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_lo_6}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_17 = &_decoded_T_16; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_9 = io_decode_0_inst[0]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_7_8 = io_decode_0_inst[28]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _decoded_T_18 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_2_6,decoded_andMatrixInput_3_6,
    decoded_andMatrixInput_4_6,decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,
    decoded_andMatrixInput_7_8,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_19 = &_decoded_T_18; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_10 = io_decode_0_inst[22]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _decoded_T_20 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,
    decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,
    decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_21 = &_decoded_T_20; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_1_11 = io_decode_0_inst[1]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_2_10 = decoded_invInputs_1[2]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_3_10 = decoded_invInputs_1[3]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_4_10 = io_decode_0_inst[4]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_5_10 = io_decode_0_inst[5]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_6_10 = io_decode_0_inst[6]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  decoded_andMatrixInput_7_10 = decoded_invInputs_1[7]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_8_10 = decoded_invInputs_1[8]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_9_10 = decoded_invInputs_1[9]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  decoded_andMatrixInput_10_5 = io_decode_0_inst[25]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] decoded_lo_10 = {decoded_andMatrixInput_9_10,decoded_andMatrixInput_10_5,decoded_andMatrixInput_6_6,
    decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,decoded_andMatrixInput_9_6,decoded_andMatrixInput_10_3,
    decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [16:0] _decoded_T_22 = {decoded_andMatrixInput_0_9,decoded_andMatrixInput_1_11,decoded_andMatrixInput_2_10,
    decoded_andMatrixInput_3_10,decoded_andMatrixInput_4_10,decoded_andMatrixInput_5_10,decoded_andMatrixInput_6_10,
    decoded_andMatrixInput_7_10,decoded_andMatrixInput_8_10,decoded_lo_10}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_23 = &_decoded_T_22; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_7_11 = io_decode_0_inst[29]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _decoded_T_24 = {decoded_andMatrixInput_0_10,decoded_andMatrixInput_3_6,decoded_andMatrixInput_4_6,
    decoded_andMatrixInput_5_6,decoded_andMatrixInput_6_6,decoded_andMatrixInput_7_6,decoded_andMatrixInput_7_8,
    decoded_andMatrixInput_7_11,decoded_andMatrixInput_10_3,decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_25 = &_decoded_T_24; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_13 = io_decode_0_inst[30]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [1:0] _decoded_T_26 = {decoded_andMatrixInput_0_13,decoded_andMatrixInput_11_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_27 = &_decoded_T_26; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  _decoded_orMatrixOutputs_T_7 = |_decoded_T_23; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_orMatrixOutputs_T_8 = |_decoded_T_21; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_orMatrixOutputs_T_9 = |_decoded_T_25; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _decoded_orMatrixOutputs_T_10 = {_decoded_T_19,_decoded_T_27}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _decoded_orMatrixOutputs_T_11 = |_decoded_orMatrixOutputs_T_10; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_orMatrixOutputs_T_12 = |_decoded_T_17; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_orMatrixOutputs_T_13 = |_decoded_T_15; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [8:0] decoded_orMatrixOutputs_1 = {_decoded_orMatrixOutputs_T_13,_decoded_orMatrixOutputs_T_12,
    _decoded_orMatrixOutputs_T_11,_decoded_orMatrixOutputs_T_9,_decoded_orMatrixOutputs_T_8,_decoded_orMatrixOutputs_T_7
    ,1'h0,2'h0}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [8:0] decoded_invMatrixOutputs_1 = {decoded_orMatrixOutputs_1[8],decoded_orMatrixOutputs_1[7],
    decoded_orMatrixOutputs_1[6],decoded_orMatrixOutputs_1[5],decoded_orMatrixOutputs_1[4],decoded_orMatrixOutputs_1[3],
    decoded_orMatrixOutputs_1[2],decoded_orMatrixOutputs_1[1],decoded_orMatrixOutputs_1[0]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire  is_ret = decoded_invMatrixOutputs_1[6]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  is_wfi = decoded_invMatrixOutputs_1[4]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  is_sfence = decoded_invMatrixOutputs_1[3]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  is_hfence_gvma = decoded_invMatrixOutputs_1[1]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  is_hlsv = decoded_invMatrixOutputs_1[0]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  _is_counter_T_2 = addr_1 >= 12'hc00 & addr_1 < 12'hc20; // @[src/main/scala/util/package.scala 205:55]
  wire  _is_counter_T_5 = addr_1 >= 12'hc80 & addr_1 < 12'hca0; // @[src/main/scala/util/package.scala 205:55]
  wire  is_counter = _is_counter_T_2 | _is_counter_T_5; // @[src/main/scala/rocket/CSR.scala 905:81]
  wire  _allow_wfi_T = reg_mstatus_prv > 2'h1; // @[src/main/scala/rocket/CSR.scala 907:61]
  wire  allow_wfi = reg_mstatus_prv > 2'h1 | ~reg_mstatus_tw; // @[src/main/scala/rocket/CSR.scala 907:71]
  wire  allow_sfence_vma = _allow_wfi_T | ~reg_mstatus_tvm; // @[src/main/scala/rocket/CSR.scala 908:70]
  wire  _allow_hfence_vvma_T_1 = reg_mstatus_prv >= 2'h1; // @[src/main/scala/rocket/CSR.scala 909:88]
  wire  allow_sret = _allow_wfi_T | ~reg_mstatus_tsr; // @[src/main/scala/rocket/CSR.scala 911:72]
  wire [4:0] counter_addr = addr_1[4:0]; // @[src/main/scala/rocket/CSR.scala 912:28]
  wire [31:0] _allow_counter_T_1 = read_mcounteren >> counter_addr; // @[src/main/scala/rocket/CSR.scala 913:70]
  wire [31:0] _allow_counter_T_7 = read_scounteren >> counter_addr; // @[src/main/scala/rocket/CSR.scala 914:75]
  wire  _allow_counter_T_9 = _allow_hfence_vvma_T_1 | _allow_counter_T_7[0]; // @[src/main/scala/rocket/CSR.scala 914:57]
  wire  allow_counter = (_allow_wfi_T | _allow_counter_T_1[0]) & _allow_counter_T_9; // @[src/main/scala/rocket/CSR.scala 913:86]
  wire [11:0] io_decode_0_fp_csr_invInputs = ~addr_1; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  csr_addr_legal = reg_mstatus_prv >= addr_1[9:8]; // @[src/main/scala/rocket/CSR.scala 920:42]
  wire  _csr_exists_T_15 = addr_1 == 12'hb02; // @[src/main/scala/rocket/CSR.scala 900:93]
  wire  _csr_exists_T_113 = addr_1 == 12'h180; // @[src/main/scala/rocket/CSR.scala 900:93]
  wire  _csr_exists_T_138 = addr_1 == 12'h301 | addr_1 == 12'h300 | addr_1 == 12'h305 | addr_1 == 12'h344 | addr_1 == 12'h304
     | addr_1 == 12'h340 | addr_1 == 12'h341 | addr_1 == 12'h343 | addr_1 == 12'h342 | addr_1 == 12'hf14 | addr_1 == 12'h7b0
     | addr_1 == 12'h7b1 | addr_1 == 12'h7b2 | addr_1 == 12'h320 | addr_1 == 12'hb00 | _csr_exists_T_15; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_153 = _csr_exists_T_138 | addr_1 == 12'h323 | addr_1 == 12'hb03 | addr_1 == 12'hc03 | addr_1 == 12'h324
     | addr_1 == 12'hb04 | addr_1 == 12'hc04 | addr_1 == 12'h325 | addr_1 == 12'hb05 | addr_1 == 12'hc05 | addr_1 == 12'h326
     | addr_1 == 12'hb06 | addr_1 == 12'hc06 | addr_1 == 12'h327 | addr_1 == 12'hb07 | addr_1 == 12'hc07; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_168 = _csr_exists_T_153 | addr_1 == 12'h328 | addr_1 == 12'hb08 | addr_1 == 12'hc08 | addr_1 == 12'h329
     | addr_1 == 12'hb09 | addr_1 == 12'hc09 | addr_1 == 12'h32a | addr_1 == 12'hb0a | addr_1 == 12'hc0a | addr_1 == 12'h32b
     | addr_1 == 12'hb0b | addr_1 == 12'hc0b | addr_1 == 12'h32c | addr_1 == 12'hb0c | addr_1 == 12'hc0c; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_183 = _csr_exists_T_168 | addr_1 == 12'h32d | addr_1 == 12'hb0d | addr_1 == 12'hc0d | addr_1 == 12'h32e
     | addr_1 == 12'hb0e | addr_1 == 12'hc0e | addr_1 == 12'h32f | addr_1 == 12'hb0f | addr_1 == 12'hc0f | addr_1 == 12'h330
     | addr_1 == 12'hb10 | addr_1 == 12'hc10 | addr_1 == 12'h331 | addr_1 == 12'hb11 | addr_1 == 12'hc11; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_198 = _csr_exists_T_183 | addr_1 == 12'h332 | addr_1 == 12'hb12 | addr_1 == 12'hc12 | addr_1 == 12'h333
     | addr_1 == 12'hb13 | addr_1 == 12'hc13 | addr_1 == 12'h334 | addr_1 == 12'hb14 | addr_1 == 12'hc14 | addr_1 == 12'h335
     | addr_1 == 12'hb15 | addr_1 == 12'hc15 | addr_1 == 12'h336 | addr_1 == 12'hb16 | addr_1 == 12'hc16; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_213 = _csr_exists_T_198 | addr_1 == 12'h337 | addr_1 == 12'hb17 | addr_1 == 12'hc17 | addr_1 == 12'h338
     | addr_1 == 12'hb18 | addr_1 == 12'hc18 | addr_1 == 12'h339 | addr_1 == 12'hb19 | addr_1 == 12'hc19 | addr_1 == 12'h33a
     | addr_1 == 12'hb1a | addr_1 == 12'hc1a | addr_1 == 12'h33b | addr_1 == 12'hb1b | addr_1 == 12'hc1b; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_228 = _csr_exists_T_213 | addr_1 == 12'h33c | addr_1 == 12'hb1c | addr_1 == 12'hc1c | addr_1 == 12'h33d
     | addr_1 == 12'hb1d | addr_1 == 12'hc1d | addr_1 == 12'h33e | addr_1 == 12'hb1e | addr_1 == 12'hc1e | addr_1 == 12'h33f
     | addr_1 == 12'hb1f | addr_1 == 12'hc1f | addr_1 == 12'h306 | addr_1 == 12'hc00 | addr_1 == 12'hc02; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _csr_exists_T_243 = _csr_exists_T_228 | addr_1 == 12'h30a | addr_1 == 12'h100 | addr_1 == 12'h144 | addr_1 == 12'h104
     | addr_1 == 12'h140 | addr_1 == 12'h142 | addr_1 == 12'h143 | addr_1 == 12'h180 | addr_1 == 12'h141 | addr_1 == 12'h105
     | addr_1 == 12'h106 | addr_1 == 12'h303 | addr_1 == 12'h302 | addr_1 == 12'h10a | addr_1 == 12'hf12; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  csr_exists = _csr_exists_T_243 | addr_1 == 12'hf11 | addr_1 == 12'hf13 | addr_1 == 12'hf15; // @[src/main/scala/rocket/CSR.scala 900:111]
  wire  _io_decode_0_read_illegal_T = ~csr_addr_legal; // @[src/main/scala/rocket/CSR.scala 923:28]
  wire  _io_decode_0_read_illegal_T_1 = ~csr_exists; // @[src/main/scala/rocket/CSR.scala 924:7]
  wire  _io_decode_0_read_illegal_T_2 = ~csr_addr_legal | _io_decode_0_read_illegal_T_1; // @[src/main/scala/rocket/CSR.scala 923:44]
  wire  _io_decode_0_read_illegal_T_6 = ~allow_sfence_vma; // @[src/main/scala/rocket/CSR.scala 925:59]
  wire  _io_decode_0_read_illegal_T_7 = (_csr_exists_T_113 | addr_1 == 12'h680) & ~allow_sfence_vma; // @[src/main/scala/rocket/CSR.scala 925:56]
  wire  _io_decode_0_read_illegal_T_8 = _io_decode_0_read_illegal_T_2 | _io_decode_0_read_illegal_T_7; // @[src/main/scala/rocket/CSR.scala 924:19]
  wire  _io_decode_0_read_illegal_T_10 = is_counter & ~allow_counter; // @[src/main/scala/rocket/CSR.scala 926:18]
  wire  _io_decode_0_read_illegal_T_11 = _io_decode_0_read_illegal_T_8 | _io_decode_0_read_illegal_T_10; // @[src/main/scala/rocket/CSR.scala 925:78]
  wire  io_decode_0_read_illegal_andMatrixInput_0 = addr_1[10]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  io_decode_0_read_illegal_andMatrixInput_1 = io_decode_0_fp_csr_invInputs[11]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [1:0] _io_decode_0_read_illegal_T_12 = {io_decode_0_read_illegal_andMatrixInput_0,
    io_decode_0_read_illegal_andMatrixInput_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _io_decode_0_read_illegal_T_13 = &_io_decode_0_read_illegal_T_12; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  io_decode_0_read_illegal_orMatrixOutputs = |_io_decode_0_read_illegal_T_13; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _io_decode_0_read_illegal_T_16 = io_decode_0_read_illegal_orMatrixOutputs & _T_244; // @[src/main/scala/rocket/CSR.scala 927:42]
  wire  _io_decode_0_read_illegal_T_17 = _io_decode_0_read_illegal_T_11 | _io_decode_0_read_illegal_T_16; // @[src/main/scala/rocket/CSR.scala 926:36]
  wire  _io_decode_0_read_illegal_T_21 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[src/main/scala/rocket/CSR.scala 929:21]
  wire [11:0] io_decode_0_write_flush_addr_m = addr_1 | 12'h300; // @[src/main/scala/rocket/CSR.scala 932:25]
  wire  _io_decode_0_system_illegal_T_4 = is_wfi & ~allow_wfi; // @[src/main/scala/rocket/CSR.scala 936:14]
  wire  _io_decode_0_system_illegal_T_5 = _io_decode_0_read_illegal_T & ~is_hlsv | _io_decode_0_system_illegal_T_4; // @[src/main/scala/rocket/CSR.scala 935:58]
  wire  _io_decode_0_system_illegal_T_7 = is_ret & ~allow_sret; // @[src/main/scala/rocket/CSR.scala 937:14]
  wire  _io_decode_0_system_illegal_T_8 = _io_decode_0_system_illegal_T_5 | _io_decode_0_system_illegal_T_7; // @[src/main/scala/rocket/CSR.scala 936:28]
  wire  _io_decode_0_system_illegal_T_14 = is_ret & io_decode_0_read_illegal_andMatrixInput_0 & addr_1[7] & _T_244; // @[src/main/scala/rocket/CSR.scala 938:37]
  wire  _io_decode_0_system_illegal_T_15 = _io_decode_0_system_illegal_T_8 | _io_decode_0_system_illegal_T_14; // @[src/main/scala/rocket/CSR.scala 937:29]
  wire  _io_decode_0_system_illegal_T_18 = (is_sfence | is_hfence_gvma) & _io_decode_0_read_illegal_T_6; // @[src/main/scala/rocket/CSR.scala 939:37]
  wire [11:0] _debugTVec_T = insn_break ? 12'h800 : 12'h808; // @[src/main/scala/rocket/CSR.scala 968:37]
  wire [11:0] debugTVec = reg_debug ? _debugTVec_T : 12'h800; // @[src/main/scala/rocket/CSR.scala 968:22]
  wire [63:0] notDebugTVec_base = delegate ? read_stvec : read_mtvec; // @[src/main/scala/rocket/CSR.scala 977:19]
  wire [7:0] notDebugTVec_interruptOffset = {cause[5:0], 2'h0}; // @[src/main/scala/rocket/CSR.scala 978:59]
  wire [63:0] notDebugTVec_interruptVec = {notDebugTVec_base[63:8],notDebugTVec_interruptOffset}; // @[src/main/scala/rocket/CSR.scala 979:27]
  wire  notDebugTVec_doVector = notDebugTVec_base[0] & cause[63] & cause_lsbs[7:6] == 2'h0; // @[src/main/scala/rocket/CSR.scala 980:55]
  wire [63:0] _notDebugTVec_T_1 = {notDebugTVec_base[63:2], 2'h0}; // @[src/main/scala/rocket/CSR.scala 981:56]
  wire [63:0] notDebugTVec = notDebugTVec_doVector ? notDebugTVec_interruptVec : _notDebugTVec_T_1; // @[src/main/scala/rocket/CSR.scala 981:8]
  wire [63:0] tvec = trapToDebug ? {{52'd0}, debugTVec} : notDebugTVec; // @[src/main/scala/rocket/CSR.scala 994:17]
  wire [1:0] _T_212 = insn_ret + insn_call; // @[src/main/scala/rocket/CSR.scala 1020:18]
  wire [1:0] _T_214 = insn_break + io_exception; // @[src/main/scala/rocket/CSR.scala 1020:18]
  wire [2:0] _T_216 = _T_212 + _T_214; // @[src/main/scala/rocket/CSR.scala 1020:18]
  wire  _T_220 = ~reset; // @[src/main/scala/rocket/CSR.scala 1020:9]
  wire  line_1043_clock;
  wire  line_1043_reset;
  wire  line_1043_valid;
  reg  line_1043_valid_reg;
  wire  _T_221 = ~(_T_216 <= 3'h1); // @[src/main/scala/rocket/CSR.scala 1020:9]
  wire  line_1044_clock;
  wire  line_1044_reset;
  wire  line_1044_valid;
  reg  line_1044_valid_reg;
  wire  _T_225 = insn_wfi & _io_interrupt_T & _T_244; // @[src/main/scala/rocket/CSR.scala 1022:36]
  wire  line_1045_clock;
  wire  line_1045_reset;
  wire  line_1045_valid;
  reg  line_1045_valid_reg;
  wire  _GEN_86 = insn_wfi & _io_interrupt_T & _T_244 | reg_wfi; // @[src/main/scala/rocket/CSR.scala 1022:{51,61} 581:54]
  wire  _T_228 = |pending_interrupts | exception; // @[src/main/scala/rocket/CSR.scala 1023:55]
  wire  line_1046_clock;
  wire  line_1046_reset;
  wire  line_1046_valid;
  reg  line_1046_valid_reg;
  wire  _T_230 = io_retire | exception; // @[src/main/scala/rocket/CSR.scala 1026:22]
  wire  line_1047_clock;
  wire  line_1047_reset;
  wire  line_1047_valid;
  reg  line_1047_valid_reg;
  wire  _GEN_88 = io_retire | exception | reg_singleStepped; // @[src/main/scala/rocket/CSR.scala 1026:{36,56} 492:30]
  wire  line_1048_clock;
  wire  line_1048_reset;
  wire  line_1048_valid;
  reg  line_1048_valid_reg;
  wire  line_1049_clock;
  wire  line_1049_reset;
  wire  line_1049_valid;
  reg  line_1049_valid_reg;
  wire  line_1050_clock;
  wire  line_1050_reset;
  wire  line_1050_valid;
  reg  line_1050_valid_reg;
  wire  _T_243 = ~(~reg_singleStepped | ~io_retire); // @[src/main/scala/rocket/CSR.scala 1029:9]
  wire  line_1051_clock;
  wire  line_1051_reset;
  wire  line_1051_valid;
  reg  line_1051_valid_reg;
  wire [39:0] _epc_T = ~io_pc; // @[src/main/scala/rocket/CSR.scala 1716:28]
  wire [39:0] _epc_T_1 = _epc_T | 40'h1; // @[src/main/scala/rocket/CSR.scala 1716:31]
  wire [39:0] epc = ~_epc_T_1; // @[src/main/scala/rocket/CSR.scala 1716:26]
  wire [39:0] tval = insn_break ? epc : io_tval; // @[src/main/scala/rocket/CSR.scala 1032:17]
  wire  line_1052_clock;
  wire  line_1052_reset;
  wire  line_1052_valid;
  reg  line_1052_valid_reg;
  wire  line_1053_clock;
  wire  line_1053_reset;
  wire  line_1053_valid;
  reg  line_1053_valid_reg;
  wire  line_1054_clock;
  wire  line_1054_reset;
  wire  line_1054_valid;
  reg  line_1054_valid_reg;
  wire [1:0] _reg_dcsr_cause_T = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[src/main/scala/rocket/CSR.scala 1040:90]
  wire [1:0] _reg_dcsr_cause_T_1 = causeIsDebugInt ? 2'h3 : _reg_dcsr_cause_T; // @[src/main/scala/rocket/CSR.scala 1040:58]
  wire [2:0] _reg_dcsr_cause_T_2 = reg_singleStepped ? 3'h4 : {{1'd0}, _reg_dcsr_cause_T_1}; // @[src/main/scala/rocket/CSR.scala 1040:30]
  wire  _GEN_91 = ~reg_debug | reg_debug; // @[src/main/scala/rocket/CSR.scala 1036:25 1038:19 488:26]
  wire [39:0] _GEN_92 = ~reg_debug ? epc : reg_dpc; // @[src/main/scala/rocket/CSR.scala 1036:25 1039:17 489:20]
  wire [1:0] _GEN_94 = ~reg_debug ? reg_mstatus_prv : reg_dcsr_prv; // @[src/main/scala/rocket/CSR.scala 1036:25 1041:22 409:25]
  wire  line_1055_clock;
  wire  line_1055_reset;
  wire  line_1055_valid;
  reg  line_1055_valid_reg;
  wire  line_1056_clock;
  wire  line_1056_reset;
  wire  line_1056_valid;
  reg  line_1056_valid_reg;
  wire  line_1057_clock;
  wire  line_1057_reset;
  wire  line_1057_valid;
  reg  line_1057_valid_reg;
  wire [39:0] _GEN_108 = delegate ? epc : reg_sepc; // @[src/main/scala/rocket/CSR.scala 1064:35 1069:16 575:21]
  wire [63:0] _GEN_109 = delegate ? cause : reg_scause; // @[src/main/scala/rocket/CSR.scala 1064:35 1070:18 576:23]
  wire [39:0] _GEN_110 = delegate ? tval : reg_stval; // @[src/main/scala/rocket/CSR.scala 1064:35 1071:17 577:22]
  wire  _GEN_112 = delegate ? reg_mstatus_sie : reg_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 1064:35 1073:24 401:28]
  wire [1:0] _GEN_113 = delegate ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp}; // @[src/main/scala/rocket/CSR.scala 1064:35 1074:23 401:28]
  wire  _GEN_114 = delegate ? 1'h0 : reg_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 1064:35 1075:23 401:28]
  wire [39:0] _GEN_118 = delegate ? reg_mepc : epc; // @[src/main/scala/rocket/CSR.scala 1064:35 1081:16 511:21]
  wire [63:0] _GEN_119 = delegate ? reg_mcause : cause; // @[src/main/scala/rocket/CSR.scala 1064:35 1082:18 512:27]
  wire [39:0] _GEN_120 = delegate ? reg_mtval : tval; // @[src/main/scala/rocket/CSR.scala 1064:35 1083:17 513:22]
  wire  _GEN_122 = delegate ? reg_mstatus_mpie : reg_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 1064:35 1085:24 401:28]
  wire [1:0] _GEN_123 = delegate ? reg_mstatus_mpp : reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 1064:35 1086:23 401:28]
  wire  _GEN_124 = delegate & reg_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 1064:35 1087:23 401:28]
  wire  _GEN_185 = trapToDebug ? _GEN_91 : reg_debug; // @[src/main/scala/rocket/CSR.scala 1035:24 488:26]
  wire [39:0] _GEN_186 = trapToDebug ? _GEN_92 : reg_dpc; // @[src/main/scala/rocket/CSR.scala 1035:24 489:20]
  wire [1:0] _GEN_188 = trapToDebug ? _GEN_94 : reg_dcsr_prv; // @[src/main/scala/rocket/CSR.scala 1035:24 409:25]
  wire [39:0] _GEN_205 = trapToDebug ? reg_sepc : _GEN_108; // @[src/main/scala/rocket/CSR.scala 1035:24 575:21]
  wire [63:0] _GEN_206 = trapToDebug ? reg_scause : _GEN_109; // @[src/main/scala/rocket/CSR.scala 1035:24 576:23]
  wire [39:0] _GEN_207 = trapToDebug ? reg_stval : _GEN_110; // @[src/main/scala/rocket/CSR.scala 1035:24 577:22]
  wire  _GEN_209 = trapToDebug ? reg_mstatus_spie : _GEN_112; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire [1:0] _GEN_210 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_113; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire  _GEN_211 = trapToDebug ? reg_mstatus_sie : _GEN_114; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire [39:0] _GEN_214 = trapToDebug ? reg_mepc : _GEN_118; // @[src/main/scala/rocket/CSR.scala 1035:24 511:21]
  wire [63:0] _GEN_215 = trapToDebug ? reg_mcause : _GEN_119; // @[src/main/scala/rocket/CSR.scala 1035:24 512:27]
  wire [39:0] _GEN_216 = trapToDebug ? reg_mtval : _GEN_120; // @[src/main/scala/rocket/CSR.scala 1035:24 513:22]
  wire  _GEN_218 = trapToDebug ? reg_mstatus_mpie : _GEN_122; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire [1:0] _GEN_219 = trapToDebug ? reg_mstatus_mpp : _GEN_123; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire  _GEN_220 = trapToDebug ? reg_mstatus_mie : _GEN_124; // @[src/main/scala/rocket/CSR.scala 1035:24 401:28]
  wire  _GEN_222 = exception ? _GEN_185 : reg_debug; // @[src/main/scala/rocket/CSR.scala 1034:20 488:26]
  wire [39:0] _GEN_223 = exception ? _GEN_186 : reg_dpc; // @[src/main/scala/rocket/CSR.scala 1034:20 489:20]
  wire [1:0] _GEN_225 = exception ? _GEN_188 : reg_dcsr_prv; // @[src/main/scala/rocket/CSR.scala 1034:20 409:25]
  wire [39:0] _GEN_242 = exception ? _GEN_205 : reg_sepc; // @[src/main/scala/rocket/CSR.scala 1034:20 575:21]
  wire [63:0] _GEN_243 = exception ? _GEN_206 : reg_scause; // @[src/main/scala/rocket/CSR.scala 1034:20 576:23]
  wire [39:0] _GEN_244 = exception ? _GEN_207 : reg_stval; // @[src/main/scala/rocket/CSR.scala 1034:20 577:22]
  wire  _GEN_246 = exception ? _GEN_209 : reg_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire [1:0] _GEN_247 = exception ? _GEN_210 : {{1'd0}, reg_mstatus_spp}; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire  _GEN_248 = exception ? _GEN_211 : reg_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire [39:0] _GEN_251 = exception ? _GEN_214 : reg_mepc; // @[src/main/scala/rocket/CSR.scala 1034:20 511:21]
  wire [63:0] _GEN_252 = exception ? _GEN_215 : reg_mcause; // @[src/main/scala/rocket/CSR.scala 1034:20 512:27]
  wire [39:0] _GEN_253 = exception ? _GEN_216 : reg_mtval; // @[src/main/scala/rocket/CSR.scala 1034:20 513:22]
  wire  _GEN_255 = exception ? _GEN_218 : reg_mstatus_mpie; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire [1:0] _GEN_256 = exception ? _GEN_219 : reg_mstatus_mpp; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire  _GEN_257 = exception ? _GEN_220 : reg_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 1034:20 401:28]
  wire  line_1058_clock;
  wire  line_1058_reset;
  wire  line_1058_valid;
  reg  line_1058_valid_reg;
  wire  line_1059_clock;
  wire  line_1059_reset;
  wire  line_1059_valid;
  reg  line_1059_valid_reg;
  wire  line_1060_clock;
  wire  line_1060_reset;
  wire  line_1060_valid;
  reg  line_1060_valid_reg;
  wire  line_1061_clock;
  wire  line_1061_reset;
  wire  line_1061_valid;
  reg  line_1061_valid_reg;
  wire  line_1062_clock;
  wire  line_1062_reset;
  wire  line_1062_valid;
  reg  line_1062_valid_reg;
  wire [39:0] _GEN_279 = io_rw_addr[10] & io_rw_addr[7] ? _T_35 : _T_23; // @[src/main/scala/rocket/CSR.scala 1131:66 1135:15]
  wire  _GEN_281 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_257 : reg_mstatus_mpie; // @[src/main/scala/rocket/CSR.scala 1131:66]
  wire  _GEN_282 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_255 : 1'h1; // @[src/main/scala/rocket/CSR.scala 1131:66]
  wire [1:0] _GEN_283 = io_rw_addr[10] & io_rw_addr[7] ? _GEN_256 : 2'h0; // @[src/main/scala/rocket/CSR.scala 1131:66]
  wire  _GEN_285 = ~io_rw_addr[9] ? reg_mstatus_spie : _GEN_248; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire  _GEN_286 = ~io_rw_addr[9] | _GEN_246; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire [1:0] _GEN_287 = ~io_rw_addr[9] ? 2'h0 : _GEN_247; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire [39:0] _GEN_290 = ~io_rw_addr[9] ? _T_50 : _GEN_279; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire  _GEN_297 = ~io_rw_addr[9] ? _GEN_257 : _GEN_281; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire  _GEN_298 = ~io_rw_addr[9] ? _GEN_255 : _GEN_282; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire [1:0] _GEN_299 = ~io_rw_addr[9] ? _GEN_256 : _GEN_283; // @[src/main/scala/rocket/CSR.scala 1114:48]
  wire  _T_380 = ret_prv <= 2'h1; // @[src/main/scala/rocket/CSR.scala 1152:34]
  wire  line_1063_clock;
  wire  line_1063_reset;
  wire  line_1063_valid;
  reg  line_1063_valid_reg;
  wire  _GEN_301 = ret_prv <= 2'h1 ? 1'h0 : reg_mstatus_mprv; // @[src/main/scala/rocket/CSR.scala 1152:46 1153:24 401:28]
  wire  _GEN_302 = insn_ret ? _GEN_285 : _GEN_248; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire  _GEN_303 = insn_ret ? _GEN_286 : _GEN_246; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire [1:0] _GEN_304 = insn_ret ? _GEN_287 : _GEN_247; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire [63:0] _GEN_306 = insn_ret ? {{24'd0}, _GEN_290} : tvec; // @[src/main/scala/rocket/CSR.scala 1112:19 995:11]
  wire  _GEN_313 = insn_ret ? _GEN_297 : _GEN_257; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire  _GEN_314 = insn_ret ? _GEN_298 : _GEN_255; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire [1:0] _GEN_315 = insn_ret ? _GEN_299 : _GEN_256; // @[src/main/scala/rocket/CSR.scala 1112:19]
  wire  _GEN_318 = insn_ret ? _GEN_301 : reg_mstatus_mprv; // @[src/main/scala/rocket/CSR.scala 1112:19 401:28]
  reg  io_status_cease_r; // @[src/main/scala/rocket/CSR.scala 1159:31]
  wire  line_1064_clock;
  wire  line_1064_reset;
  wire  line_1064_valid;
  reg  line_1064_valid_reg;
  wire [63:0] _io_rw_rdata_T = decoded_0 ? reg_misa : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_1 = decoded_1 ? read_mstatus : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_2 = decoded_2 ? read_mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _io_rw_rdata_T_3 = decoded_3 ? read_mip : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_4 = decoded_4 ? reg_mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_5 = decoded_5 ? reg_mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_6 = decoded_6 ? _T_26 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_7 = decoded_7 ? _T_29 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_8 = decoded_8 ? reg_mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_rw_rdata_T_9 = decoded_9 & io_hartid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_rw_rdata_T_10 = decoded_10 ? _T_30 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_11 = decoded_11 ? _T_38 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_12 = decoded_12 ? reg_dscratch0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_14 = decoded_14 ? value_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_15 = decoded_15 ? value : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_rw_rdata_T_103 = decoded_103 ? read_mcounteren : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_104 = decoded_104 ? value_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_105 = decoded_105 ? value : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_107 = decoded_107 ? _sstatus_T[63:0] : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_108 = decoded_108 ? read_sip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_109 = decoded_109 ? read_sie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_110 = decoded_110 ? reg_sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_111 = decoded_111 ? reg_scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_112 = decoded_112 ? _T_44 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_113 = decoded_113 ? _T_45 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_114 = decoded_114 ? _T_53 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_115 = decoded_115 ? read_stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_rw_rdata_T_116 = decoded_116 ? read_scounteren : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_117 = decoded_117 ? read_mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_118 = decoded_118 ? read_medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_120 = decoded_120 ? 64'h1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_122 = decoded_122 ? 64'h20181004 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_124 = _io_rw_rdata_T | _io_rw_rdata_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_125 = _io_rw_rdata_T_124 | _io_rw_rdata_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_474 = {{48'd0}, _io_rw_rdata_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_126 = _io_rw_rdata_T_125 | _GEN_474; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_127 = _io_rw_rdata_T_126 | _io_rw_rdata_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_128 = _io_rw_rdata_T_127 | _io_rw_rdata_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_129 = _io_rw_rdata_T_128 | _io_rw_rdata_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_130 = _io_rw_rdata_T_129 | _io_rw_rdata_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_131 = _io_rw_rdata_T_130 | _io_rw_rdata_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_475 = {{63'd0}, _io_rw_rdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_132 = _io_rw_rdata_T_131 | _GEN_475; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_476 = {{32'd0}, _io_rw_rdata_T_10}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_133 = _io_rw_rdata_T_132 | _GEN_476; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_134 = _io_rw_rdata_T_133 | _io_rw_rdata_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_135 = _io_rw_rdata_T_134 | _io_rw_rdata_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_137 = _io_rw_rdata_T_135 | _io_rw_rdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_138 = _io_rw_rdata_T_137 | _io_rw_rdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_477 = {{32'd0}, _io_rw_rdata_T_103}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_226 = _io_rw_rdata_T_138 | _GEN_477; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_227 = _io_rw_rdata_T_226 | _io_rw_rdata_T_104; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_228 = _io_rw_rdata_T_227 | _io_rw_rdata_T_105; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_230 = _io_rw_rdata_T_228 | _io_rw_rdata_T_107; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_231 = _io_rw_rdata_T_230 | _io_rw_rdata_T_108; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_232 = _io_rw_rdata_T_231 | _io_rw_rdata_T_109; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_233 = _io_rw_rdata_T_232 | _io_rw_rdata_T_110; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_234 = _io_rw_rdata_T_233 | _io_rw_rdata_T_111; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_235 = _io_rw_rdata_T_234 | _io_rw_rdata_T_112; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_236 = _io_rw_rdata_T_235 | _io_rw_rdata_T_113; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_237 = _io_rw_rdata_T_236 | _io_rw_rdata_T_114; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_238 = _io_rw_rdata_T_237 | _io_rw_rdata_T_115; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_478 = {{32'd0}, _io_rw_rdata_T_116}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_239 = _io_rw_rdata_T_238 | _GEN_478; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_240 = _io_rw_rdata_T_239 | _io_rw_rdata_T_117; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_241 = _io_rw_rdata_T_240 | _io_rw_rdata_T_118; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_rw_rdata_T_243 = _io_rw_rdata_T_241 | _io_rw_rdata_T_120; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_384 = io_rw_cmd == 3'h5; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_385 = io_rw_cmd == 3'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_386 = io_rw_cmd == 3'h7; // @[src/main/scala/util/package.scala 16:47]
  wire  _csr_wen_T_4 = _T_385 | _T_386 | _T_384; // @[src/main/scala/util/package.scala 73:59]
  wire  csr_wen = _csr_wen_T_4 & ~io_rw_stall; // @[src/main/scala/rocket/CSR.scala 1222:56]
  wire  line_1065_clock;
  wire  line_1065_reset;
  wire  line_1065_valid;
  reg  line_1065_valid_reg;
  wire  line_1066_clock;
  wire  line_1066_reset;
  wire  line_1066_valid;
  reg  line_1066_valid_reg;
  wire [104:0] _new_mstatus_WIRE = {{41'd0}, wdata}; // @[src/main/scala/rocket/CSR.scala 1229:{39,39}]
  wire  new_mstatus_sie = _new_mstatus_WIRE[1]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_mie = _new_mstatus_WIRE[3]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_spie = _new_mstatus_WIRE[5]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_mpie = _new_mstatus_WIRE[7]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_spp = _new_mstatus_WIRE[8]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire [1:0] new_mstatus_mpp = _new_mstatus_WIRE[12:11]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire [1:0] new_mstatus_fs = _new_mstatus_WIRE[14:13]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_mprv = _new_mstatus_WIRE[17]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_sum = _new_mstatus_WIRE[18]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_mxr = _new_mstatus_WIRE[19]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_tvm = _new_mstatus_WIRE[20]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_tw = _new_mstatus_WIRE[21]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire  new_mstatus_tsr = _new_mstatus_WIRE[22]; // @[src/main/scala/rocket/CSR.scala 1229:39]
  wire [1:0] _reg_mstatus_fs_T_1 = |new_mstatus_fs ? 2'h3 : 2'h0; // @[src/main/scala/rocket/CSR.scala 1720:66]
  wire [1:0] _GEN_326 = decoded_1 ? {{1'd0}, new_mstatus_spp} : _GEN_304; // @[src/main/scala/rocket/CSR.scala 1228:39 1237:27]
  wire  line_1067_clock;
  wire  line_1067_reset;
  wire  line_1067_valid;
  reg  line_1067_valid_reg;
  wire  f = wdata[5]; // @[src/main/scala/rocket/CSR.scala 1259:20]
  wire  _T_1527 = ~io_pc[1] | wdata[2]; // @[src/main/scala/rocket/CSR.scala 1261:45]
  wire  line_1068_clock;
  wire  line_1068_reset;
  wire  line_1068_valid;
  reg  line_1068_valid_reg;
  wire [63:0] _reg_misa_T = ~wdata; // @[src/main/scala/rocket/CSR.scala 1263:25]
  wire  _reg_misa_T_1 = ~f; // @[src/main/scala/rocket/CSR.scala 1263:35]
  wire [3:0] _reg_misa_T_2 = {_reg_misa_T_1, 3'h0}; // @[src/main/scala/rocket/CSR.scala 1263:38]
  wire [63:0] _GEN_479 = {{60'd0}, _reg_misa_T_2}; // @[src/main/scala/rocket/CSR.scala 1263:32]
  wire [63:0] _reg_misa_T_3 = _reg_misa_T | _GEN_479; // @[src/main/scala/rocket/CSR.scala 1263:32]
  wire [63:0] _reg_misa_T_4 = ~_reg_misa_T_3; // @[src/main/scala/rocket/CSR.scala 1263:23]
  wire [63:0] _reg_misa_T_5 = _reg_misa_T_4 & 64'h1005; // @[src/main/scala/rocket/CSR.scala 1263:55]
  wire [63:0] _reg_misa_T_7 = reg_misa & 64'hffffffffffffeffa; // @[src/main/scala/rocket/CSR.scala 1263:73]
  wire [63:0] _reg_misa_T_8 = _reg_misa_T_5 | _reg_misa_T_7; // @[src/main/scala/rocket/CSR.scala 1263:62]
  wire  line_1069_clock;
  wire  line_1069_reset;
  wire  line_1069_valid;
  reg  line_1069_valid_reg;
  wire [15:0] _new_mip_T_2 = io_rw_cmd[1] ? _read_hvip_T : 16'h0; // @[src/main/scala/rocket/CSR.scala 1695:9]
  wire [63:0] _GEN_480 = {{48'd0}, _new_mip_T_2}; // @[src/main/scala/rocket/CSR.scala 1695:30]
  wire [63:0] _new_mip_T_3 = _GEN_480 | io_rw_wdata; // @[src/main/scala/rocket/CSR.scala 1695:30]
  wire [63:0] _new_mip_T_8 = _new_mip_T_3 & _wdata_T_6; // @[src/main/scala/rocket/CSR.scala 1695:39]
  wire  new_mip_ssip = _new_mip_T_8[1]; // @[src/main/scala/rocket/CSR.scala 1271:88]
  wire  new_mip_stip = _new_mip_T_8[5]; // @[src/main/scala/rocket/CSR.scala 1271:88]
  wire  new_mip_seip = _new_mip_T_8[9]; // @[src/main/scala/rocket/CSR.scala 1271:88]
  wire  line_1070_clock;
  wire  line_1070_reset;
  wire  line_1070_valid;
  reg  line_1070_valid_reg;
  wire [63:0] _reg_mie_T = wdata & 64'haaa; // @[src/main/scala/rocket/CSR.scala 1281:59]
  wire  line_1071_clock;
  wire  line_1071_reset;
  wire  line_1071_valid;
  reg  line_1071_valid_reg;
  wire [63:0] _reg_mepc_T_1 = _reg_misa_T | 64'h1; // @[src/main/scala/rocket/CSR.scala 1716:31]
  wire [63:0] _reg_mepc_T_2 = ~_reg_mepc_T_1; // @[src/main/scala/rocket/CSR.scala 1716:26]
  wire [63:0] _GEN_342 = decoded_6 ? _reg_mepc_T_2 : {{24'd0}, _GEN_251}; // @[src/main/scala/rocket/CSR.scala 1282:{40,51}]
  wire  line_1072_clock;
  wire  line_1072_reset;
  wire  line_1072_valid;
  reg  line_1072_valid_reg;
  wire  line_1073_clock;
  wire  line_1073_reset;
  wire  line_1073_valid;
  reg  line_1073_valid_reg;
  wire [63:0] _GEN_344 = decoded_2 ? wdata : {{32'd0}, reg_mtvec}; // @[src/main/scala/rocket/CSR.scala 1285:{40,52} 518:31]
  wire  line_1074_clock;
  wire  line_1074_reset;
  wire  line_1074_valid;
  reg  line_1074_valid_reg;
  wire  line_1075_clock;
  wire  line_1075_reset;
  wire  line_1075_valid;
  reg  line_1075_valid_reg;
  wire [63:0] _GEN_346 = decoded_7 ? wdata : {{24'd0}, _GEN_253}; // @[src/main/scala/rocket/CSR.scala 1287:{40,52}]
  wire  line_1076_clock;
  wire  line_1076_reset;
  wire  line_1076_valid;
  reg  line_1076_valid_reg;
  wire [63:0] _GEN_347 = decoded_14 ? wdata : {{57'd0}, nextSmall_1}; // @[src/main/scala/rocket/CSR.scala 1713:31 src/main/scala/util/Counters.scala 67:11]
  wire  line_1077_clock;
  wire  line_1077_reset;
  wire  line_1077_valid;
  reg  line_1077_valid_reg;
  wire [63:0] _GEN_349 = decoded_15 ? wdata : {{57'd0}, nextSmall}; // @[src/main/scala/rocket/CSR.scala 1713:31 src/main/scala/util/Counters.scala 67:11]
  wire  line_1078_clock;
  wire  line_1078_reset;
  wire  line_1078_valid;
  reg  line_1078_valid_reg;
  wire [1:0] new_dcsr_prv = wdata[1:0]; // @[src/main/scala/rocket/CSR.scala 1322:38]
  wire  new_dcsr_step = wdata[2]; // @[src/main/scala/rocket/CSR.scala 1322:38]
  wire  new_dcsr_ebreaku = wdata[12]; // @[src/main/scala/rocket/CSR.scala 1322:38]
  wire  new_dcsr_ebreaks = wdata[13]; // @[src/main/scala/rocket/CSR.scala 1322:38]
  wire  new_dcsr_ebreakm = wdata[15]; // @[src/main/scala/rocket/CSR.scala 1322:38]
  wire  line_1079_clock;
  wire  line_1079_reset;
  wire  line_1079_valid;
  reg  line_1079_valid_reg;
  wire [63:0] _GEN_356 = decoded_11 ? _reg_mepc_T_2 : {{24'd0}, _GEN_223}; // @[src/main/scala/rocket/CSR.scala 1330:{42,52}]
  wire  line_1080_clock;
  wire  line_1080_reset;
  wire  line_1080_valid;
  reg  line_1080_valid_reg;
  wire  line_1081_clock;
  wire  line_1081_reset;
  wire  line_1081_valid;
  reg  line_1081_valid_reg;
  wire [1:0] _GEN_360 = decoded_107 ? {{1'd0}, new_mstatus_spp} : _GEN_326; // @[src/main/scala/rocket/CSR.scala 1341:41 1345:25]
  wire  line_1082_clock;
  wire  line_1082_reset;
  wire  line_1082_valid;
  reg  line_1082_valid_reg;
  wire [63:0] _new_sip_T = ~read_mideleg; // @[src/main/scala/rocket/CSR.scala 1354:36]
  wire [63:0] _new_sip_T_1 = _GEN_464 & _new_sip_T; // @[src/main/scala/rocket/CSR.scala 1354:34]
  wire [63:0] _new_sip_T_2 = wdata & read_mideleg; // @[src/main/scala/rocket/CSR.scala 1354:60]
  wire [63:0] _new_sip_T_3 = _new_sip_T_1 | _new_sip_T_2; // @[src/main/scala/rocket/CSR.scala 1354:51]
  wire  new_sip_ssip = _new_sip_T_3[1]; // @[src/main/scala/rocket/CSR.scala 1354:85]
  wire  line_1083_clock;
  wire  line_1083_reset;
  wire  line_1083_valid;
  reg  line_1083_valid_reg;
  wire [43:0] new_satp_ppn = wdata[43:0]; // @[src/main/scala/rocket/CSR.scala 1359:40]
  wire [3:0] new_satp_mode = wdata[63:60]; // @[src/main/scala/rocket/CSR.scala 1359:40]
  wire  _T_1530 = new_satp_mode == 4'h0; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_1531 = new_satp_mode == 4'h8; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_1532 = _T_1530 | _T_1531; // @[src/main/scala/util/package.scala 73:59]
  wire  line_1084_clock;
  wire  line_1084_reset;
  wire  line_1084_valid;
  reg  line_1084_valid_reg;
  wire [3:0] _reg_satp_mode_T = new_satp_mode & 4'h8; // @[src/main/scala/rocket/CSR.scala 1361:44]
  wire  line_1085_clock;
  wire  line_1085_reset;
  wire  line_1085_valid;
  reg  line_1085_valid_reg;
  wire [63:0] _reg_mie_T_1 = ~sie_mask; // @[src/main/scala/rocket/CSR.scala 1367:66]
  wire [63:0] _reg_mie_T_2 = reg_mie & _reg_mie_T_1; // @[src/main/scala/rocket/CSR.scala 1367:64]
  wire [63:0] _reg_mie_T_3 = wdata & sie_mask; // @[src/main/scala/rocket/CSR.scala 1367:86]
  wire [63:0] _reg_mie_T_4 = _reg_mie_T_2 | _reg_mie_T_3; // @[src/main/scala/rocket/CSR.scala 1367:77]
  wire  line_1086_clock;
  wire  line_1086_reset;
  wire  line_1086_valid;
  reg  line_1086_valid_reg;
  wire  line_1087_clock;
  wire  line_1087_reset;
  wire  line_1087_valid;
  reg  line_1087_valid_reg;
  wire [63:0] _GEN_372 = decoded_114 ? _reg_mepc_T_2 : {{24'd0}, _GEN_242}; // @[src/main/scala/rocket/CSR.scala 1369:{42,53}]
  wire  line_1088_clock;
  wire  line_1088_reset;
  wire  line_1088_valid;
  reg  line_1088_valid_reg;
  wire [63:0] _GEN_373 = decoded_115 ? wdata : {{25'd0}, reg_stvec}; // @[src/main/scala/rocket/CSR.scala 1370:{42,54} 579:22]
  wire  line_1089_clock;
  wire  line_1089_reset;
  wire  line_1089_valid;
  reg  line_1089_valid_reg;
  wire  line_1090_clock;
  wire  line_1090_reset;
  wire  line_1090_valid;
  reg  line_1090_valid_reg;
  wire [63:0] _GEN_375 = decoded_112 ? wdata : {{24'd0}, _GEN_244}; // @[src/main/scala/rocket/CSR.scala 1372:{42,54}]
  wire  line_1091_clock;
  wire  line_1091_reset;
  wire  line_1091_valid;
  reg  line_1091_valid_reg;
  wire  line_1092_clock;
  wire  line_1092_reset;
  wire  line_1092_valid;
  reg  line_1092_valid_reg;
  wire  line_1093_clock;
  wire  line_1093_reset;
  wire  line_1093_valid;
  reg  line_1093_valid_reg;
  wire [63:0] _GEN_378 = decoded_116 ? wdata : {{32'd0}, reg_scounteren}; // @[src/main/scala/rocket/CSR.scala 1375:{44,61} 541:22]
  wire  line_1094_clock;
  wire  line_1094_reset;
  wire  line_1094_valid;
  reg  line_1094_valid_reg;
  wire [63:0] _GEN_379 = decoded_103 ? wdata : {{32'd0}, reg_mcounteren}; // @[src/main/scala/rocket/CSR.scala 1451:{44,61} 537:22]
  wire  line_1095_clock;
  wire  line_1095_reset;
  wire  line_1095_valid;
  reg  line_1095_valid_reg;
  wire  line_1096_clock;
  wire  line_1096_reset;
  wire  line_1096_valid;
  reg  line_1096_valid_reg;
  wire  line_1097_clock;
  wire  line_1097_reset;
  wire  line_1097_valid;
  reg  line_1097_valid_reg;
  wire [1:0] _GEN_390 = csr_wen ? _GEN_360 : _GEN_304; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_405 = csr_wen ? _GEN_342 : {{24'd0}, _GEN_251}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_407 = csr_wen ? _GEN_344 : {{32'd0}, reg_mtvec}; // @[src/main/scala/rocket/CSR.scala 1224:18 518:31]
  wire [63:0] _GEN_409 = csr_wen ? _GEN_346 : {{24'd0}, _GEN_253}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_410 = csr_wen ? _GEN_347 : {{57'd0}, nextSmall_1}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_412 = csr_wen ? _GEN_349 : {{57'd0}, nextSmall}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_419 = csr_wen ? _GEN_356 : {{24'd0}, _GEN_223}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_424 = csr_wen ? _GEN_372 : {{24'd0}, _GEN_242}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_425 = csr_wen ? _GEN_373 : {{25'd0}, reg_stvec}; // @[src/main/scala/rocket/CSR.scala 1224:18 579:22]
  wire [63:0] _GEN_427 = csr_wen ? _GEN_375 : {{24'd0}, _GEN_244}; // @[src/main/scala/rocket/CSR.scala 1224:18]
  wire [63:0] _GEN_430 = csr_wen ? _GEN_378 : {{32'd0}, reg_scounteren}; // @[src/main/scala/rocket/CSR.scala 1224:18 541:22]
  wire [63:0] _GEN_431 = csr_wen ? _GEN_379 : {{32'd0}, reg_mcounteren}; // @[src/main/scala/rocket/CSR.scala 1224:18 537:22]
  wire  line_1098_clock;
  wire  line_1098_reset;
  wire  line_1098_valid;
  reg  line_1098_valid_reg;
  wire  line_1099_clock;
  wire  line_1099_reset;
  wire  line_1099_valid;
  reg  line_1099_valid_reg;
  wire  line_1100_clock;
  wire  line_1100_reset;
  wire  line_1100_valid;
  reg  line_1100_valid_reg;
  wire [2:0] _io_trace_0_priv_T = {reg_debug,reg_mstatus_prv}; // @[src/main/scala/rocket/CSR.scala 1629:18]
  wire [63:0] _difftest_interrupt_T_2 = exception & cause[63] ? cause : 64'h0; // @[src/main/scala/rocket/CSR.scala 1640:34]
  wire [63:0] _difftest_exception_T_3 = exception & _causeIsDebugTrigger_T_1 ? cause : 64'h0; // @[src/main/scala/rocket/CSR.scala 1641:34]
  reg [63:0] cycleCnt; // @[src/main/scala/rocket/CSR.scala 1647:27]
  wire [63:0] _cycleCnt_T_1 = cycleCnt + 64'h1; // @[src/main/scala/rocket/CSR.scala 1648:26]
  wire  _difftest_hasTrap_T_2 = io_trace_0_valid & ~(io_trace_0_exception | io_trace_0_interrupt); // @[src/main/scala/rocket/CSR.scala 236:30]
  wire [31:0] _difftest_hasTrap_T_3 = io_trace_0_insn & 32'h707f; // @[src/main/scala/rocket/CSR.scala 237:31]
  wire  _difftest_hasTrap_T_4 = 32'h6b == _difftest_hasTrap_T_3; // @[src/main/scala/rocket/CSR.scala 237:31]
  wire [1:0] _GEN_484 = reset ? 2'h0 : _GEN_390; // @[src/main/scala/rocket/CSR.scala 401:{28,28}]
  wire [63:0] _GEN_485 = reset ? 64'h0 : _GEN_407; // @[src/main/scala/rocket/CSR.scala 518:{31,31}]
  wire [63:0] _GEN_486 = reset ? 64'h0 : _GEN_431; // @[src/main/scala/rocket/CSR.scala 537:{22,22}]
  wire [63:0] _GEN_487 = reset ? 64'h0 : _GEN_430; // @[src/main/scala/rocket/CSR.scala 541:{22,22}]
  wire [63:0] _GEN_488 = reset ? 64'h0 : _GEN_412; // @[src/main/scala/util/Counters.scala 45:{41,41}]
  wire [63:0] _GEN_489 = reset ? 64'h0 : _GEN_410; // @[src/main/scala/util/Counters.scala 45:{41,41}]
  DelayReg_2 difftest_delayer ( // @[difftest/src/main/scala/util/Delayer.scala 54:15]
    .clock(difftest_delayer_clock),
    .reset(difftest_delayer_reset),
    .i_valid(difftest_delayer_i_valid),
    .i_interrupt(difftest_delayer_i_interrupt),
    .i_exception(difftest_delayer_i_exception),
    .i_exceptionPC(difftest_delayer_i_exceptionPC),
    .i_exceptionInst(difftest_delayer_i_exceptionInst),
    .o_valid(difftest_delayer_o_valid),
    .o_interrupt(difftest_delayer_o_interrupt),
    .o_exception(difftest_delayer_o_exception),
    .o_exceptionPC(difftest_delayer_o_exceptionPC),
    .o_exceptionInst(difftest_delayer_o_exceptionInst)
  );
  DummyDPICWrapper_2 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_interrupt(difftest_module_io_bits_interrupt),
    .io_bits_exception(difftest_module_io_bits_exception),
    .io_bits_exceptionPC(difftest_module_io_bits_exceptionPC),
    .io_bits_exceptionInst(difftest_module_io_bits_exceptionInst)
  );
  DummyDPICWrapper_3 difftest_module_1 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_1_clock),
    .reset(difftest_module_1_reset),
    .io_bits_hasTrap(difftest_module_1_io_bits_hasTrap),
    .io_bits_cycleCnt(difftest_module_1_io_bits_cycleCnt),
    .io_bits_instrCnt(difftest_module_1_io_bits_instrCnt),
    .io_bits_pc(difftest_module_1_io_bits_pc)
  );
  GEN_w1_line #(.COVER_INDEX(1041)) line_1041 (
    .clock(line_1041_clock),
    .reset(line_1041_reset),
    .valid(line_1041_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1042)) line_1042 (
    .clock(line_1042_clock),
    .reset(line_1042_reset),
    .valid(line_1042_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1043)) line_1043 (
    .clock(line_1043_clock),
    .reset(line_1043_reset),
    .valid(line_1043_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1044)) line_1044 (
    .clock(line_1044_clock),
    .reset(line_1044_reset),
    .valid(line_1044_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1045)) line_1045 (
    .clock(line_1045_clock),
    .reset(line_1045_reset),
    .valid(line_1045_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1046)) line_1046 (
    .clock(line_1046_clock),
    .reset(line_1046_reset),
    .valid(line_1046_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1047)) line_1047 (
    .clock(line_1047_clock),
    .reset(line_1047_reset),
    .valid(line_1047_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1048)) line_1048 (
    .clock(line_1048_clock),
    .reset(line_1048_reset),
    .valid(line_1048_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1049)) line_1049 (
    .clock(line_1049_clock),
    .reset(line_1049_reset),
    .valid(line_1049_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1050)) line_1050 (
    .clock(line_1050_clock),
    .reset(line_1050_reset),
    .valid(line_1050_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1051)) line_1051 (
    .clock(line_1051_clock),
    .reset(line_1051_reset),
    .valid(line_1051_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1052)) line_1052 (
    .clock(line_1052_clock),
    .reset(line_1052_reset),
    .valid(line_1052_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1053)) line_1053 (
    .clock(line_1053_clock),
    .reset(line_1053_reset),
    .valid(line_1053_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1054)) line_1054 (
    .clock(line_1054_clock),
    .reset(line_1054_reset),
    .valid(line_1054_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1055)) line_1055 (
    .clock(line_1055_clock),
    .reset(line_1055_reset),
    .valid(line_1055_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1056)) line_1056 (
    .clock(line_1056_clock),
    .reset(line_1056_reset),
    .valid(line_1056_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1057)) line_1057 (
    .clock(line_1057_clock),
    .reset(line_1057_reset),
    .valid(line_1057_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1058)) line_1058 (
    .clock(line_1058_clock),
    .reset(line_1058_reset),
    .valid(line_1058_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1059)) line_1059 (
    .clock(line_1059_clock),
    .reset(line_1059_reset),
    .valid(line_1059_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1060)) line_1060 (
    .clock(line_1060_clock),
    .reset(line_1060_reset),
    .valid(line_1060_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1061)) line_1061 (
    .clock(line_1061_clock),
    .reset(line_1061_reset),
    .valid(line_1061_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1062)) line_1062 (
    .clock(line_1062_clock),
    .reset(line_1062_reset),
    .valid(line_1062_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1063)) line_1063 (
    .clock(line_1063_clock),
    .reset(line_1063_reset),
    .valid(line_1063_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1064)) line_1064 (
    .clock(line_1064_clock),
    .reset(line_1064_reset),
    .valid(line_1064_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1065)) line_1065 (
    .clock(line_1065_clock),
    .reset(line_1065_reset),
    .valid(line_1065_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1066)) line_1066 (
    .clock(line_1066_clock),
    .reset(line_1066_reset),
    .valid(line_1066_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1067)) line_1067 (
    .clock(line_1067_clock),
    .reset(line_1067_reset),
    .valid(line_1067_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1068)) line_1068 (
    .clock(line_1068_clock),
    .reset(line_1068_reset),
    .valid(line_1068_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1069)) line_1069 (
    .clock(line_1069_clock),
    .reset(line_1069_reset),
    .valid(line_1069_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1070)) line_1070 (
    .clock(line_1070_clock),
    .reset(line_1070_reset),
    .valid(line_1070_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1071)) line_1071 (
    .clock(line_1071_clock),
    .reset(line_1071_reset),
    .valid(line_1071_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1072)) line_1072 (
    .clock(line_1072_clock),
    .reset(line_1072_reset),
    .valid(line_1072_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1073)) line_1073 (
    .clock(line_1073_clock),
    .reset(line_1073_reset),
    .valid(line_1073_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1074)) line_1074 (
    .clock(line_1074_clock),
    .reset(line_1074_reset),
    .valid(line_1074_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1075)) line_1075 (
    .clock(line_1075_clock),
    .reset(line_1075_reset),
    .valid(line_1075_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1076)) line_1076 (
    .clock(line_1076_clock),
    .reset(line_1076_reset),
    .valid(line_1076_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1077)) line_1077 (
    .clock(line_1077_clock),
    .reset(line_1077_reset),
    .valid(line_1077_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1078)) line_1078 (
    .clock(line_1078_clock),
    .reset(line_1078_reset),
    .valid(line_1078_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1079)) line_1079 (
    .clock(line_1079_clock),
    .reset(line_1079_reset),
    .valid(line_1079_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1080)) line_1080 (
    .clock(line_1080_clock),
    .reset(line_1080_reset),
    .valid(line_1080_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1081)) line_1081 (
    .clock(line_1081_clock),
    .reset(line_1081_reset),
    .valid(line_1081_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1082)) line_1082 (
    .clock(line_1082_clock),
    .reset(line_1082_reset),
    .valid(line_1082_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1083)) line_1083 (
    .clock(line_1083_clock),
    .reset(line_1083_reset),
    .valid(line_1083_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1084)) line_1084 (
    .clock(line_1084_clock),
    .reset(line_1084_reset),
    .valid(line_1084_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1085)) line_1085 (
    .clock(line_1085_clock),
    .reset(line_1085_reset),
    .valid(line_1085_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1086)) line_1086 (
    .clock(line_1086_clock),
    .reset(line_1086_reset),
    .valid(line_1086_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1087)) line_1087 (
    .clock(line_1087_clock),
    .reset(line_1087_reset),
    .valid(line_1087_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1088)) line_1088 (
    .clock(line_1088_clock),
    .reset(line_1088_reset),
    .valid(line_1088_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1089)) line_1089 (
    .clock(line_1089_clock),
    .reset(line_1089_reset),
    .valid(line_1089_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1090)) line_1090 (
    .clock(line_1090_clock),
    .reset(line_1090_reset),
    .valid(line_1090_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1091)) line_1091 (
    .clock(line_1091_clock),
    .reset(line_1091_reset),
    .valid(line_1091_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1092)) line_1092 (
    .clock(line_1092_clock),
    .reset(line_1092_reset),
    .valid(line_1092_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1093)) line_1093 (
    .clock(line_1093_clock),
    .reset(line_1093_reset),
    .valid(line_1093_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1094)) line_1094 (
    .clock(line_1094_clock),
    .reset(line_1094_reset),
    .valid(line_1094_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1095)) line_1095 (
    .clock(line_1095_clock),
    .reset(line_1095_reset),
    .valid(line_1095_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1096)) line_1096 (
    .clock(line_1096_clock),
    .reset(line_1096_reset),
    .valid(line_1096_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1097)) line_1097 (
    .clock(line_1097_clock),
    .reset(line_1097_reset),
    .valid(line_1097_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1098)) line_1098 (
    .clock(line_1098_clock),
    .reset(line_1098_reset),
    .valid(line_1098_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1099)) line_1099 (
    .clock(line_1099_clock),
    .reset(line_1099_reset),
    .valid(line_1099_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1100)) line_1100 (
    .clock(line_1100_clock),
    .reset(line_1100_reset),
    .valid(line_1100_valid)
  );
  assign line_1041_clock = clock;
  assign line_1041_reset = reset;
  assign line_1041_valid = nextSmall[6] ^ line_1041_valid_reg;
  assign line_1042_clock = clock;
  assign line_1042_reset = reset;
  assign line_1042_valid = nextSmall_1[6] ^ line_1042_valid_reg;
  assign line_1043_clock = clock;
  assign line_1043_reset = reset;
  assign line_1043_valid = _T_220 ^ line_1043_valid_reg;
  assign line_1044_clock = clock;
  assign line_1044_reset = reset;
  assign line_1044_valid = _T_221 ^ line_1044_valid_reg;
  assign line_1045_clock = clock;
  assign line_1045_reset = reset;
  assign line_1045_valid = _T_225 ^ line_1045_valid_reg;
  assign line_1046_clock = clock;
  assign line_1046_reset = reset;
  assign line_1046_valid = _T_228 ^ line_1046_valid_reg;
  assign line_1047_clock = clock;
  assign line_1047_reset = reset;
  assign line_1047_valid = _T_230 ^ line_1047_valid_reg;
  assign line_1048_clock = clock;
  assign line_1048_reset = reset;
  assign line_1048_valid = _io_interrupt_T ^ line_1048_valid_reg;
  assign line_1049_clock = clock;
  assign line_1049_reset = reset;
  assign line_1049_valid = _T_220 ^ line_1049_valid_reg;
  assign line_1050_clock = clock;
  assign line_1050_reset = reset;
  assign line_1050_valid = _T_220 ^ line_1050_valid_reg;
  assign line_1051_clock = clock;
  assign line_1051_reset = reset;
  assign line_1051_valid = _T_243 ^ line_1051_valid_reg;
  assign line_1052_clock = clock;
  assign line_1052_reset = reset;
  assign line_1052_valid = exception ^ line_1052_valid_reg;
  assign line_1053_clock = clock;
  assign line_1053_reset = reset;
  assign line_1053_valid = trapToDebug ^ line_1053_valid_reg;
  assign line_1054_clock = clock;
  assign line_1054_reset = reset;
  assign line_1054_valid = _T_244 ^ line_1054_valid_reg;
  assign line_1055_clock = clock;
  assign line_1055_reset = reset;
  assign line_1055_valid = trapToDebug ^ line_1055_valid_reg;
  assign line_1056_clock = clock;
  assign line_1056_reset = reset;
  assign line_1056_valid = delegate ^ line_1056_valid_reg;
  assign line_1057_clock = clock;
  assign line_1057_reset = reset;
  assign line_1057_valid = delegate ^ line_1057_valid_reg;
  assign line_1058_clock = clock;
  assign line_1058_reset = reset;
  assign line_1058_valid = insn_ret ^ line_1058_valid_reg;
  assign line_1059_clock = clock;
  assign line_1059_reset = reset;
  assign line_1059_valid = _T_368 ^ line_1059_valid_reg;
  assign line_1060_clock = clock;
  assign line_1060_reset = reset;
  assign line_1060_valid = _T_368 ^ line_1060_valid_reg;
  assign line_1061_clock = clock;
  assign line_1061_reset = reset;
  assign line_1061_valid = _T_374 ^ line_1061_valid_reg;
  assign line_1062_clock = clock;
  assign line_1062_reset = reset;
  assign line_1062_valid = _T_374 ^ line_1062_valid_reg;
  assign line_1063_clock = clock;
  assign line_1063_reset = reset;
  assign line_1063_valid = _T_380 ^ line_1063_valid_reg;
  assign line_1064_clock = clock;
  assign line_1064_reset = reset;
  assign line_1064_valid = insn_cease ^ line_1064_valid_reg;
  assign line_1065_clock = clock;
  assign line_1065_reset = reset;
  assign line_1065_valid = csr_wen ^ line_1065_valid_reg;
  assign line_1066_clock = clock;
  assign line_1066_reset = reset;
  assign line_1066_valid = decoded_1 ^ line_1066_valid_reg;
  assign line_1067_clock = clock;
  assign line_1067_reset = reset;
  assign line_1067_valid = decoded_0 ^ line_1067_valid_reg;
  assign line_1068_clock = clock;
  assign line_1068_reset = reset;
  assign line_1068_valid = _T_1527 ^ line_1068_valid_reg;
  assign line_1069_clock = clock;
  assign line_1069_reset = reset;
  assign line_1069_valid = decoded_3 ^ line_1069_valid_reg;
  assign line_1070_clock = clock;
  assign line_1070_reset = reset;
  assign line_1070_valid = decoded_4 ^ line_1070_valid_reg;
  assign line_1071_clock = clock;
  assign line_1071_reset = reset;
  assign line_1071_valid = decoded_6 ^ line_1071_valid_reg;
  assign line_1072_clock = clock;
  assign line_1072_reset = reset;
  assign line_1072_valid = decoded_5 ^ line_1072_valid_reg;
  assign line_1073_clock = clock;
  assign line_1073_reset = reset;
  assign line_1073_valid = decoded_2 ^ line_1073_valid_reg;
  assign line_1074_clock = clock;
  assign line_1074_reset = reset;
  assign line_1074_valid = decoded_8 ^ line_1074_valid_reg;
  assign line_1075_clock = clock;
  assign line_1075_reset = reset;
  assign line_1075_valid = decoded_7 ^ line_1075_valid_reg;
  assign line_1076_clock = clock;
  assign line_1076_reset = reset;
  assign line_1076_valid = decoded_14 ^ line_1076_valid_reg;
  assign line_1077_clock = clock;
  assign line_1077_reset = reset;
  assign line_1077_valid = decoded_15 ^ line_1077_valid_reg;
  assign line_1078_clock = clock;
  assign line_1078_reset = reset;
  assign line_1078_valid = decoded_10 ^ line_1078_valid_reg;
  assign line_1079_clock = clock;
  assign line_1079_reset = reset;
  assign line_1079_valid = decoded_11 ^ line_1079_valid_reg;
  assign line_1080_clock = clock;
  assign line_1080_reset = reset;
  assign line_1080_valid = decoded_12 ^ line_1080_valid_reg;
  assign line_1081_clock = clock;
  assign line_1081_reset = reset;
  assign line_1081_valid = decoded_107 ^ line_1081_valid_reg;
  assign line_1082_clock = clock;
  assign line_1082_reset = reset;
  assign line_1082_valid = decoded_108 ^ line_1082_valid_reg;
  assign line_1083_clock = clock;
  assign line_1083_reset = reset;
  assign line_1083_valid = decoded_113 ^ line_1083_valid_reg;
  assign line_1084_clock = clock;
  assign line_1084_reset = reset;
  assign line_1084_valid = _T_1532 ^ line_1084_valid_reg;
  assign line_1085_clock = clock;
  assign line_1085_reset = reset;
  assign line_1085_valid = decoded_109 ^ line_1085_valid_reg;
  assign line_1086_clock = clock;
  assign line_1086_reset = reset;
  assign line_1086_valid = decoded_110 ^ line_1086_valid_reg;
  assign line_1087_clock = clock;
  assign line_1087_reset = reset;
  assign line_1087_valid = decoded_114 ^ line_1087_valid_reg;
  assign line_1088_clock = clock;
  assign line_1088_reset = reset;
  assign line_1088_valid = decoded_115 ^ line_1088_valid_reg;
  assign line_1089_clock = clock;
  assign line_1089_reset = reset;
  assign line_1089_valid = decoded_111 ^ line_1089_valid_reg;
  assign line_1090_clock = clock;
  assign line_1090_reset = reset;
  assign line_1090_valid = decoded_112 ^ line_1090_valid_reg;
  assign line_1091_clock = clock;
  assign line_1091_reset = reset;
  assign line_1091_valid = decoded_117 ^ line_1091_valid_reg;
  assign line_1092_clock = clock;
  assign line_1092_reset = reset;
  assign line_1092_valid = decoded_118 ^ line_1092_valid_reg;
  assign line_1093_clock = clock;
  assign line_1093_reset = reset;
  assign line_1093_valid = decoded_116 ^ line_1093_valid_reg;
  assign line_1094_clock = clock;
  assign line_1094_reset = reset;
  assign line_1094_valid = decoded_103 ^ line_1094_valid_reg;
  assign line_1095_clock = clock;
  assign line_1095_reset = reset;
  assign line_1095_valid = decoded_120 ^ line_1095_valid_reg;
  assign line_1096_clock = clock;
  assign line_1096_reset = reset;
  assign line_1096_valid = decoded_121 ^ line_1096_valid_reg;
  assign line_1097_clock = clock;
  assign line_1097_reset = reset;
  assign line_1097_valid = decoded_122 ^ line_1097_valid_reg;
  assign line_1098_clock = clock;
  assign line_1098_reset = reset;
  assign line_1098_valid = reset ^ line_1098_valid_reg;
  assign line_1099_clock = clock;
  assign line_1099_reset = reset;
  assign line_1099_valid = reset ^ line_1099_valid_reg;
  assign line_1100_clock = clock;
  assign line_1100_reset = reset;
  assign line_1100_valid = reset ^ line_1100_valid_reg;
  assign io_rw_rdata = _io_rw_rdata_T_243 | _io_rw_rdata_T_122; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_decode_0_fp_illegal = io_status_fs == 2'h0 | ~reg_misa[5]; // @[src/main/scala/rocket/CSR.scala 916:91]
  assign io_decode_0_fp_csr = 1'h0; // @[src/main/scala/rocket/Decode.scala 58:116]
  assign io_decode_0_rocc_illegal = io_status_xs == 2'h0 | ~reg_misa[23]; // @[src/main/scala/rocket/CSR.scala 919:93]
  assign io_decode_0_read_illegal = _io_decode_0_read_illegal_T_17 | _io_decode_0_read_illegal_T_21; // @[src/main/scala/rocket/CSR.scala 928:68]
  assign io_decode_0_write_illegal = &addr_1[11:10]; // @[src/main/scala/rocket/CSR.scala 930:41]
  assign io_decode_0_write_flush = ~(io_decode_0_write_flush_addr_m >= 12'h340 & io_decode_0_write_flush_addr_m <= 12'h343
    ); // @[src/main/scala/rocket/CSR.scala 933:7]
  assign io_decode_0_system_illegal = _io_decode_0_system_illegal_T_15 | _io_decode_0_system_illegal_T_18; // @[src/main/scala/rocket/CSR.scala 938:51]
  assign io_csr_stall = reg_wfi | io_status_cease; // @[src/main/scala/rocket/CSR.scala 1158:27]
  assign io_rw_stall = 1'h0; // @[src/main/scala/rocket/CSR.scala 809:{33,47}]
  assign io_eret = _exception_T | insn_ret; // @[src/main/scala/rocket/CSR.scala 999:38]
  assign io_singleStep = reg_dcsr_step & _T_244; // @[src/main/scala/rocket/CSR.scala 1000:34]
  assign io_status_debug = reg_debug; // @[src/main/scala/rocket/CSR.scala 1003:19]
  assign io_status_cease = io_status_cease_r; // @[src/main/scala/rocket/CSR.scala 1159:19]
  assign io_status_wfi = reg_wfi; // @[src/main/scala/rocket/CSR.scala 1160:17]
  assign io_status_isa = reg_misa[31:0]; // @[src/main/scala/rocket/CSR.scala 1004:17]
  assign io_status_dprv = reg_mstatus_mprv & _T_244 ? reg_mstatus_mpp : reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 1007:24]
  assign io_status_dv = 1'h0; // @[src/main/scala/rocket/CSR.scala 1008:39]
  assign io_status_prv = reg_mstatus_prv; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_v = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_sd = &io_status_fs | &io_status_xs | &io_status_vs; // @[src/main/scala/rocket/CSR.scala 1002:58]
  assign io_status_zero2 = 23'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mpv = 1'h0; // @[src/main/scala/rocket/CSR.scala 1010:17]
  assign io_status_gva = reg_mstatus_gva; // @[src/main/scala/rocket/CSR.scala 1011:17]
  assign io_status_mbe = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_sbe = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_sxl = 2'h2; // @[src/main/scala/rocket/CSR.scala 1006:17]
  assign io_status_uxl = 2'h2; // @[src/main/scala/rocket/CSR.scala 1005:17]
  assign io_status_sd_rv32 = 1'h0; // @[src/main/scala/rocket/CSR.scala 1009:39]
  assign io_status_zero1 = 8'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_tsr = reg_mstatus_tsr; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_tw = reg_mstatus_tw; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_tvm = reg_mstatus_tvm; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mxr = reg_mstatus_mxr; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_sum = reg_mstatus_sum; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mprv = reg_mstatus_mprv; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_xs = 2'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_fs = reg_mstatus_fs; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mpp = reg_mstatus_mpp; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_vs = 2'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_spp = reg_mstatus_spp; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_ube = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_spie = reg_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_upie = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_mie = reg_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_hie = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_sie = reg_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_status_uie = 1'h0; // @[src/main/scala/rocket/CSR.scala 1001:13]
  assign io_ptbr_mode = reg_satp_mode; // @[src/main/scala/rocket/CSR.scala 996:11]
  assign io_ptbr_ppn = reg_satp_ppn; // @[src/main/scala/rocket/CSR.scala 996:11]
  assign io_evec = _GEN_306[39:0];
  assign io_time = {large_1,small_1}; // @[src/main/scala/util/Counters.scala 55:30]
  assign io_interrupt = (anyInterrupt & ~io_singleStep | reg_singleStepped) & ~(reg_debug | io_status_cease); // @[src/main/scala/rocket/CSR.scala 626:73]
  assign io_interrupt_cause = 64'h8000000000000000 + _GEN_465; // @[src/main/scala/rocket/CSR.scala 625:63]
  assign io_csrr_counter = decoded_14 | decoded_104; // @[src/main/scala/rocket/CSR.scala 1220:48]
  assign io_trace_0_valid = io_retire > 1'h0 | io_trace_0_exception; // @[src/main/scala/rocket/CSR.scala 1626:32]
  assign io_trace_0_iaddr = io_pc; // @[src/main/scala/rocket/CSR.scala 1628:13]
  assign io_trace_0_insn = io_inst_0; // @[src/main/scala/rocket/CSR.scala 1627:12]
  assign io_trace_0_exception = insn_call | insn_break | io_exception; // @[src/main/scala/rocket/CSR.scala 1019:43]
  assign io_trace_0_interrupt = cause[63]; // @[src/main/scala/rocket/CSR.scala 1631:25]
  assign io_difftest_privilegeMode = {{61'd0}, _io_trace_0_priv_T}; // @[src/main/scala/rocket/CSR.scala 1660:29]
  assign io_difftest_mstatus = _read_mstatus_T[63:0]; // @[src/main/scala/util/package.scala 155:13]
  assign io_difftest_sstatus = _sstatus_T[63:0]; // @[src/main/scala/rocket/CSR.scala 774:{37,37}]
  assign io_difftest_mepc = {_T_25,_T_23}; // @[src/main/scala/util/package.scala 124:15]
  assign io_difftest_sepc = {_T_52,_T_50}; // @[src/main/scala/util/package.scala 124:15]
  assign io_difftest_mtval = {_T_28,reg_mtval}; // @[src/main/scala/util/package.scala 124:15]
  assign io_difftest_stval = {_T_43,reg_stval}; // @[src/main/scala/util/package.scala 124:15]
  assign io_difftest_mtvec = {32'h0,_read_mtvec_T_5}; // @[src/main/scala/util/package.scala 130:15]
  assign io_difftest_stvec = {_read_stvec_T_7,_read_stvec_T_5}; // @[src/main/scala/util/package.scala 124:15]
  assign io_difftest_mcause = reg_mcause; // @[src/main/scala/rocket/CSR.scala 1669:22]
  assign io_difftest_scause = reg_scause; // @[src/main/scala/rocket/CSR.scala 1670:22]
  assign io_difftest_satp = {hi_7,reg_satp_ppn}; // @[src/main/scala/rocket/CSR.scala 1671:32]
  assign io_difftest_mip = {{48'd0}, _read_hvip_T}; // @[src/main/scala/rocket/CSR.scala 1672:19]
  assign io_difftest_mie = reg_mie; // @[src/main/scala/rocket/CSR.scala 1673:19]
  assign io_difftest_mscratch = reg_mscratch; // @[src/main/scala/rocket/CSR.scala 1674:24]
  assign io_difftest_sscratch = reg_sscratch; // @[src/main/scala/rocket/CSR.scala 1675:24]
  assign io_difftest_mideleg = reg_mideleg & 64'h222; // @[src/main/scala/rocket/CSR.scala 504:38]
  assign io_difftest_medeleg = reg_medeleg & 64'hb15d; // @[src/main/scala/rocket/CSR.scala 508:38]
  assign io_snapshot_minstret = {large_,small_}; // @[src/main/scala/util/Counters.scala 55:30]
  assign io_snapshot_mcycle = {large_1,small_1}; // @[src/main/scala/util/Counters.scala 55:30]
  assign difftest_delayer_clock = clock;
  assign difftest_delayer_reset = reset;
  assign difftest_delayer_i_valid = insn_call | insn_break | io_exception; // @[src/main/scala/rocket/CSR.scala 1019:43]
  assign difftest_delayer_i_interrupt = _difftest_interrupt_T_2[31:0]; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1640:28]
  assign difftest_delayer_i_exception = _difftest_exception_T_3[31:0]; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1641:28]
  assign difftest_delayer_i_exceptionPC = {{24'd0}, io_pc}; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1642:28]
  assign difftest_delayer_i_exceptionInst = io_inst_0; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1643:28]
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 158:15]
  assign difftest_module_io_bits_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_io_bits_interrupt = difftest_delayer_o_interrupt; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_io_bits_exception = difftest_delayer_o_exception; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_io_bits_exceptionPC = difftest_delayer_o_exceptionPC; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_io_bits_exceptionInst = difftest_delayer_o_exceptionInst; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_1_clock = clock;
  assign difftest_module_1_reset = reset;
  assign difftest_module_1_io_bits_hasTrap = _difftest_hasTrap_T_2 & _difftest_hasTrap_T_4; // @[src/main/scala/rocket/CSR.scala 1651:47]
  assign difftest_module_1_io_bits_cycleCnt = cycleCnt; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1653:23]
  assign difftest_module_1_io_bits_instrCnt = {large_,small_}; // @[src/main/scala/util/Counters.scala 55:30]
  assign difftest_module_1_io_bits_pc = {{24'd0}, io_pc}; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/CSR.scala 1656:23]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_prv <= 2'h3; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (new_prv == 2'h2) begin // @[src/main/scala/rocket/CSR.scala 1699:29]
      reg_mstatus_prv <= 2'h0;
    end else if (insn_ret) begin // @[src/main/scala/rocket/CSR.scala 1112:19]
      if (~io_rw_addr[9]) begin // @[src/main/scala/rocket/CSR.scala 1114:48]
        reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
      end else begin
        reg_mstatus_prv <= _GEN_276;
      end
    end else if (exception) begin // @[src/main/scala/rocket/CSR.scala 1034:20]
      reg_mstatus_prv <= _GEN_190;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_gva <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (exception) begin // @[src/main/scala/rocket/CSR.scala 1034:20]
      if (!(trapToDebug)) begin // @[src/main/scala/rocket/CSR.scala 1035:24]
        if (!(delegate)) begin // @[src/main/scala/rocket/CSR.scala 1064:35]
          reg_mstatus_gva <= io_gva; // @[src/main/scala/rocket/CSR.scala 1080:23]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_tsr <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_tsr <= new_mstatus_tsr; // @[src/main/scala/rocket/CSR.scala 1241:27]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_tw <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_tw <= new_mstatus_tw; // @[src/main/scala/rocket/CSR.scala 1240:26]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_tvm <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_tvm <= new_mstatus_tvm; // @[src/main/scala/rocket/CSR.scala 1246:27]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_mxr <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_107) begin // @[src/main/scala/rocket/CSR.scala 1341:41]
        reg_mstatus_mxr <= new_mstatus_mxr; // @[src/main/scala/rocket/CSR.scala 1349:27]
      end else if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_mxr <= new_mstatus_mxr; // @[src/main/scala/rocket/CSR.scala 1244:27]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_sum <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_107) begin // @[src/main/scala/rocket/CSR.scala 1341:41]
        reg_mstatus_sum <= new_mstatus_sum; // @[src/main/scala/rocket/CSR.scala 1350:27]
      end else if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_sum <= new_mstatus_sum; // @[src/main/scala/rocket/CSR.scala 1245:27]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_mprv <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_mprv <= new_mstatus_mprv; // @[src/main/scala/rocket/CSR.scala 1234:26]
      end else begin
        reg_mstatus_mprv <= _GEN_318;
      end
    end else begin
      reg_mstatus_mprv <= _GEN_318;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_fs <= 2'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_107) begin // @[src/main/scala/rocket/CSR.scala 1341:41]
        reg_mstatus_fs <= _reg_mstatus_fs_T_1; // @[src/main/scala/rocket/CSR.scala 1346:24]
      end else if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_fs <= _reg_mstatus_fs_T_1; // @[src/main/scala/rocket/CSR.scala 1254:55]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_mpp <= 2'h3; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        if (new_mstatus_mpp == 2'h2) begin // @[src/main/scala/rocket/CSR.scala 1699:29]
          reg_mstatus_mpp <= 2'h0;
        end else begin
          reg_mstatus_mpp <= new_mstatus_mpp;
        end
      end else begin
        reg_mstatus_mpp <= _GEN_315;
      end
    end else begin
      reg_mstatus_mpp <= _GEN_315;
    end
    reg_mstatus_spp <= _GEN_484[0]; // @[src/main/scala/rocket/CSR.scala 401:{28,28}]
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_mpie <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_mpie <= new_mstatus_mpie; // @[src/main/scala/rocket/CSR.scala 1231:24]
      end else begin
        reg_mstatus_mpie <= _GEN_314;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_314;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_spie <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_107) begin // @[src/main/scala/rocket/CSR.scala 1341:41]
        reg_mstatus_spie <= new_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 1344:26]
      end else if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_spie <= new_mstatus_spie; // @[src/main/scala/rocket/CSR.scala 1238:28]
      end else begin
        reg_mstatus_spie <= _GEN_303;
      end
    end else begin
      reg_mstatus_spie <= _GEN_303;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_mie <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_mie <= new_mstatus_mie; // @[src/main/scala/rocket/CSR.scala 1230:23]
      end else begin
        reg_mstatus_mie <= _GEN_313;
      end
    end else begin
      reg_mstatus_mie <= _GEN_313;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 401:28]
      reg_mstatus_sie <= 1'h0; // @[src/main/scala/rocket/CSR.scala 401:28]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_107) begin // @[src/main/scala/rocket/CSR.scala 1341:41]
        reg_mstatus_sie <= new_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 1343:25]
      end else if (decoded_1) begin // @[src/main/scala/rocket/CSR.scala 1228:39]
        reg_mstatus_sie <= new_mstatus_sie; // @[src/main/scala/rocket/CSR.scala 1239:27]
      end else begin
        reg_mstatus_sie <= _GEN_302;
      end
    end else begin
      reg_mstatus_sie <= _GEN_302;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_prv <= 2'h3; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_10) begin // @[src/main/scala/rocket/CSR.scala 1321:38]
        if (new_dcsr_prv == 2'h2) begin // @[src/main/scala/rocket/CSR.scala 1699:29]
          reg_dcsr_prv <= 2'h0;
        end else begin
          reg_dcsr_prv <= new_dcsr_prv;
        end
      end else begin
        reg_dcsr_prv <= _GEN_225;
      end
    end else begin
      reg_dcsr_prv <= _GEN_225;
    end
    if (_io_interrupt_T) begin // @[src/main/scala/rocket/CSR.scala 1027:25]
      reg_singleStepped <= 1'h0; // @[src/main/scala/rocket/CSR.scala 1027:45]
    end else begin
      reg_singleStepped <= _GEN_88;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_ebreakm <= 1'h0; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_10) begin // @[src/main/scala/rocket/CSR.scala 1321:38]
        reg_dcsr_ebreakm <= new_dcsr_ebreakm; // @[src/main/scala/rocket/CSR.scala 1324:26]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_ebreaks <= 1'h0; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_10) begin // @[src/main/scala/rocket/CSR.scala 1321:38]
        reg_dcsr_ebreaks <= new_dcsr_ebreaks; // @[src/main/scala/rocket/CSR.scala 1325:47]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_ebreaku <= 1'h0; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_10) begin // @[src/main/scala/rocket/CSR.scala 1321:38]
        reg_dcsr_ebreaku <= new_dcsr_ebreaku; // @[src/main/scala/rocket/CSR.scala 1326:41]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 488:26]
      reg_debug <= 1'h0; // @[src/main/scala/rocket/CSR.scala 488:26]
    end else if (insn_ret) begin // @[src/main/scala/rocket/CSR.scala 1112:19]
      if (~io_rw_addr[9]) begin // @[src/main/scala/rocket/CSR.scala 1114:48]
        reg_debug <= _GEN_222;
      end else if (io_rw_addr[10] & io_rw_addr[7]) begin // @[src/main/scala/rocket/CSR.scala 1131:66]
        reg_debug <= 1'h0; // @[src/main/scala/rocket/CSR.scala 1134:17]
      end else begin
        reg_debug <= _GEN_222;
      end
    end else begin
      reg_debug <= _GEN_222;
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1562:22]
      reg_mideleg <= 64'h0; // @[src/main/scala/rocket/CSR.scala 1567:20]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_117) begin // @[src/main/scala/rocket/CSR.scala 1373:42]
        reg_mideleg <= wdata; // @[src/main/scala/rocket/CSR.scala 1373:56]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1562:22]
      reg_medeleg <= 64'h0; // @[src/main/scala/rocket/CSR.scala 1568:20]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_118) begin // @[src/main/scala/rocket/CSR.scala 1374:42]
        reg_medeleg <= wdata; // @[src/main/scala/rocket/CSR.scala 1374:56]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_cause <= 3'h0; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (exception) begin // @[src/main/scala/rocket/CSR.scala 1034:20]
      if (trapToDebug) begin // @[src/main/scala/rocket/CSR.scala 1035:24]
        if (~reg_debug) begin // @[src/main/scala/rocket/CSR.scala 1036:25]
          reg_dcsr_cause <= _reg_dcsr_cause_T_2; // @[src/main/scala/rocket/CSR.scala 1040:24]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 409:25]
      reg_dcsr_step <= 1'h0; // @[src/main/scala/rocket/CSR.scala 409:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_10) begin // @[src/main/scala/rocket/CSR.scala 1321:38]
        reg_dcsr_step <= new_dcsr_step; // @[src/main/scala/rocket/CSR.scala 1323:23]
      end
    end
    reg_dpc <= _GEN_419[39:0];
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_12) begin // @[src/main/scala/rocket/CSR.scala 1331:43]
        reg_dscratch0 <= wdata; // @[src/main/scala/rocket/CSR.scala 1331:59]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1562:22]
      reg_mie <= 64'h0; // @[src/main/scala/rocket/CSR.scala 1566:20]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_109) begin // @[src/main/scala/rocket/CSR.scala 1367:42]
        reg_mie <= _reg_mie_T_4; // @[src/main/scala/rocket/CSR.scala 1367:52]
      end else if (decoded_4) begin // @[src/main/scala/rocket/CSR.scala 1281:40]
        reg_mie <= _reg_mie_T; // @[src/main/scala/rocket/CSR.scala 1281:50]
      end
    end
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_3) begin // @[src/main/scala/rocket/CSR.scala 1266:35]
        reg_mip_seip <= new_mip_seip; // @[src/main/scala/rocket/CSR.scala 1275:22]
      end
    end
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_3) begin // @[src/main/scala/rocket/CSR.scala 1266:35]
        reg_mip_stip <= new_mip_stip; // @[src/main/scala/rocket/CSR.scala 1274:22]
      end
    end
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_108) begin // @[src/main/scala/rocket/CSR.scala 1353:37]
        reg_mip_ssip <= new_sip_ssip; // @[src/main/scala/rocket/CSR.scala 1355:22]
      end else if (decoded_3) begin // @[src/main/scala/rocket/CSR.scala 1266:35]
        reg_mip_ssip <= new_mip_ssip; // @[src/main/scala/rocket/CSR.scala 1273:22]
      end
    end
    reg_mepc <= _GEN_405[39:0];
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 512:27]
      reg_mcause <= 64'h0; // @[src/main/scala/rocket/CSR.scala 512:27]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_8) begin // @[src/main/scala/rocket/CSR.scala 1286:40]
        reg_mcause <= wdata; // @[src/main/scala/rocket/CSR.scala 1286:53]
      end else begin
        reg_mcause <= _GEN_252;
      end
    end else begin
      reg_mcause <= _GEN_252;
    end
    reg_mtval <= _GEN_409[39:0];
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_5) begin // @[src/main/scala/rocket/CSR.scala 1283:40]
        reg_mscratch <= wdata; // @[src/main/scala/rocket/CSR.scala 1283:55]
      end
    end
    reg_mtvec <= _GEN_485[31:0]; // @[src/main/scala/rocket/CSR.scala 518:{31,31}]
    reg_mcounteren <= _GEN_486[31:0]; // @[src/main/scala/rocket/CSR.scala 537:{22,22}]
    reg_scounteren <= _GEN_487[31:0]; // @[src/main/scala/rocket/CSR.scala 541:{22,22}]
    reg_sepc <= _GEN_424[39:0];
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_111) begin // @[src/main/scala/rocket/CSR.scala 1371:42]
        reg_scause <= wdata; // @[src/main/scala/rocket/CSR.scala 1371:55]
      end else begin
        reg_scause <= _GEN_243;
      end
    end else begin
      reg_scause <= _GEN_243;
    end
    reg_stval <= _GEN_427[39:0];
    if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_110) begin // @[src/main/scala/rocket/CSR.scala 1368:42]
        reg_sscratch <= wdata; // @[src/main/scala/rocket/CSR.scala 1368:57]
      end
    end
    reg_stvec <= _GEN_425[38:0];
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1562:22]
      reg_satp_mode <= 4'h0; // @[src/main/scala/rocket/CSR.scala 1563:20]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_113) begin // @[src/main/scala/rocket/CSR.scala 1357:38]
        if (_T_1532) begin // @[src/main/scala/rocket/CSR.scala 1360:67]
          reg_satp_mode <= _reg_satp_mode_T; // @[src/main/scala/rocket/CSR.scala 1361:27]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1562:22]
      reg_satp_ppn <= 44'h0; // @[src/main/scala/rocket/CSR.scala 1565:20]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_113) begin // @[src/main/scala/rocket/CSR.scala 1357:38]
        if (_T_1532) begin // @[src/main/scala/rocket/CSR.scala 1360:67]
          reg_satp_ppn <= {{24'd0}, new_satp_ppn[19:0]}; // @[src/main/scala/rocket/CSR.scala 1362:26]
        end
      end
    end
    small_ <= _GEN_488[5:0]; // @[src/main/scala/util/Counters.scala 45:{41,41}]
    if (reset) begin // @[src/main/scala/util/Counters.scala 50:31]
      large_ <= 58'h0; // @[src/main/scala/util/Counters.scala 50:31]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_15) begin // @[src/main/scala/rocket/CSR.scala 1713:31]
        large_ <= wdata[63:6]; // @[src/main/scala/util/Counters.scala 68:23]
      end else begin
        large_ <= _GEN_80;
      end
    end else begin
      large_ <= _GEN_80;
    end
    line_1041_valid_reg <= nextSmall[6];
    line_1042_valid_reg <= nextSmall_1[6];
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 650:25]
      reg_misa <= 64'h8000000000141105; // @[src/main/scala/rocket/CSR.scala 650:25]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_0) begin // @[src/main/scala/rocket/CSR.scala 1257:36]
        if (~io_pc[1] | wdata[2]) begin // @[src/main/scala/rocket/CSR.scala 1261:66]
          reg_misa <= _reg_misa_T_8; // @[src/main/scala/rocket/CSR.scala 1263:20]
        end
      end
    end
    line_1043_valid_reg <= _T_220;
    line_1044_valid_reg <= _T_221;
    line_1045_valid_reg <= _T_225;
    line_1046_valid_reg <= _T_228;
    line_1047_valid_reg <= _T_230;
    line_1048_valid_reg <= _io_interrupt_T;
    line_1049_valid_reg <= _T_220;
    line_1050_valid_reg <= _T_220;
    line_1051_valid_reg <= _T_243;
    line_1052_valid_reg <= exception;
    line_1053_valid_reg <= trapToDebug;
    line_1054_valid_reg <= _T_244;
    line_1055_valid_reg <= trapToDebug;
    line_1056_valid_reg <= delegate;
    line_1057_valid_reg <= delegate;
    line_1058_valid_reg <= insn_ret;
    line_1059_valid_reg <= _T_368;
    line_1060_valid_reg <= _T_368;
    line_1061_valid_reg <= _T_374;
    line_1062_valid_reg <= _T_374;
    line_1063_valid_reg <= _T_380;
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1159:31]
      io_status_cease_r <= 1'h0; // @[src/main/scala/rocket/CSR.scala 1159:31]
    end else begin
      io_status_cease_r <= insn_cease | io_status_cease_r;
    end
    line_1064_valid_reg <= insn_cease;
    line_1065_valid_reg <= csr_wen;
    line_1066_valid_reg <= decoded_1;
    line_1067_valid_reg <= decoded_0;
    line_1068_valid_reg <= _T_1527;
    line_1069_valid_reg <= decoded_3;
    line_1070_valid_reg <= decoded_4;
    line_1071_valid_reg <= decoded_6;
    line_1072_valid_reg <= decoded_5;
    line_1073_valid_reg <= decoded_2;
    line_1074_valid_reg <= decoded_8;
    line_1075_valid_reg <= decoded_7;
    line_1076_valid_reg <= decoded_14;
    line_1077_valid_reg <= decoded_15;
    line_1078_valid_reg <= decoded_10;
    line_1079_valid_reg <= decoded_11;
    line_1080_valid_reg <= decoded_12;
    line_1081_valid_reg <= decoded_107;
    line_1082_valid_reg <= decoded_108;
    line_1083_valid_reg <= decoded_113;
    line_1084_valid_reg <= _T_1532;
    line_1085_valid_reg <= decoded_109;
    line_1086_valid_reg <= decoded_110;
    line_1087_valid_reg <= decoded_114;
    line_1088_valid_reg <= decoded_115;
    line_1089_valid_reg <= decoded_111;
    line_1090_valid_reg <= decoded_112;
    line_1091_valid_reg <= decoded_117;
    line_1092_valid_reg <= decoded_118;
    line_1093_valid_reg <= decoded_116;
    line_1094_valid_reg <= decoded_103;
    line_1095_valid_reg <= decoded_120;
    line_1096_valid_reg <= decoded_121;
    line_1097_valid_reg <= decoded_122;
    line_1098_valid_reg <= reset;
    line_1099_valid_reg <= reset;
    line_1100_valid_reg <= reset;
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 1647:27]
      cycleCnt <= 64'h0; // @[src/main/scala/rocket/CSR.scala 1647:27]
    end else begin
      cycleCnt <= _cycleCnt_T_1; // @[src/main/scala/rocket/CSR.scala 1648:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_T_216 <= 3'h1)) begin
          $fwrite(32'h80000002,
            "Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:1020 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1.U, \"these conditions must be mutually exclusive\")\n"
            ); // @[src/main/scala/rocket/CSR.scala 1020:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_220 & ~(~reg_singleStepped | ~io_retire)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at CSR.scala:1029 assert(!reg_singleStepped || io.retire === 0.U)\n"); // @[src/main/scala/rocket/CSR.scala 1029:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge io_ungated_clock) begin
    if (reset) begin // @[src/main/scala/rocket/CSR.scala 581:54]
      reg_wfi <= 1'h0; // @[src/main/scala/rocket/CSR.scala 581:54]
    end else if (|pending_interrupts | exception) begin // @[src/main/scala/rocket/CSR.scala 1023:69]
      reg_wfi <= 1'h0; // @[src/main/scala/rocket/CSR.scala 1023:79]
    end else begin
      reg_wfi <= _GEN_86;
    end
    small_1 <= _GEN_489[5:0]; // @[src/main/scala/util/Counters.scala 45:{41,41}]
    if (reset) begin // @[src/main/scala/util/Counters.scala 50:31]
      large_1 <= 58'h0; // @[src/main/scala/util/Counters.scala 50:31]
    end else if (csr_wen) begin // @[src/main/scala/rocket/CSR.scala 1224:18]
      if (decoded_14) begin // @[src/main/scala/rocket/CSR.scala 1713:31]
        large_1 <= wdata[63:6]; // @[src/main/scala/util/Counters.scala 68:23]
      end else begin
        large_1 <= _GEN_82;
      end
    end else begin
      large_1 <= _GEN_82;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_gva = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_tsr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_tw = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_tvm = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_mxr = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_sum = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reg_mstatus_spie = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  reg_mstatus_sie = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  reg_singleStepped = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_dcsr_ebreaks = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  reg_debug = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  reg_mideleg = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  reg_medeleg = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_24[0:0];
  _RAND_25 = {2{`RANDOM}};
  reg_dpc = _RAND_25[39:0];
  _RAND_26 = {2{`RANDOM}};
  reg_dscratch0 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  reg_mie = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  reg_mip_seip = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reg_mip_stip = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  reg_mip_ssip = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  reg_mepc = _RAND_31[39:0];
  _RAND_32 = {2{`RANDOM}};
  reg_mcause = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  reg_mtval = _RAND_33[39:0];
  _RAND_34 = {2{`RANDOM}};
  reg_mscratch = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  reg_mtvec = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_mcounteren = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_scounteren = _RAND_37[31:0];
  _RAND_38 = {2{`RANDOM}};
  reg_sepc = _RAND_38[39:0];
  _RAND_39 = {2{`RANDOM}};
  reg_scause = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  reg_stval = _RAND_40[39:0];
  _RAND_41 = {2{`RANDOM}};
  reg_sscratch = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  reg_stvec = _RAND_42[38:0];
  _RAND_43 = {1{`RANDOM}};
  reg_satp_mode = _RAND_43[3:0];
  _RAND_44 = {2{`RANDOM}};
  reg_satp_ppn = _RAND_44[43:0];
  _RAND_45 = {1{`RANDOM}};
  reg_wfi = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  small_ = _RAND_46[5:0];
  _RAND_47 = {2{`RANDOM}};
  large_ = _RAND_47[57:0];
  _RAND_48 = {1{`RANDOM}};
  line_1041_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  small_1 = _RAND_49[5:0];
  _RAND_50 = {2{`RANDOM}};
  large_1 = _RAND_50[57:0];
  _RAND_51 = {1{`RANDOM}};
  line_1042_valid_reg = _RAND_51[0:0];
  _RAND_52 = {2{`RANDOM}};
  reg_misa = _RAND_52[63:0];
  _RAND_53 = {1{`RANDOM}};
  line_1043_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_1044_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_1045_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_1046_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_1047_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_1048_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_1049_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_1050_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_1051_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_1052_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_1053_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_1054_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_1055_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_1056_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_1057_valid_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  line_1058_valid_reg = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  line_1059_valid_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  line_1060_valid_reg = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  line_1061_valid_reg = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  line_1062_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  line_1063_valid_reg = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  io_status_cease_r = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  line_1064_valid_reg = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  line_1065_valid_reg = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  line_1066_valid_reg = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  line_1067_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  line_1068_valid_reg = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  line_1069_valid_reg = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  line_1070_valid_reg = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  line_1071_valid_reg = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  line_1072_valid_reg = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  line_1073_valid_reg = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  line_1074_valid_reg = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  line_1075_valid_reg = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  line_1076_valid_reg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  line_1077_valid_reg = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  line_1078_valid_reg = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  line_1079_valid_reg = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  line_1080_valid_reg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  line_1081_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  line_1082_valid_reg = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  line_1083_valid_reg = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  line_1084_valid_reg = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  line_1085_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  line_1086_valid_reg = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  line_1087_valid_reg = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  line_1088_valid_reg = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  line_1089_valid_reg = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  line_1090_valid_reg = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  line_1091_valid_reg = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  line_1092_valid_reg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  line_1093_valid_reg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  line_1094_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  line_1095_valid_reg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  line_1096_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  line_1097_valid_reg = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  line_1098_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  line_1099_valid_reg = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  line_1100_valid_reg = _RAND_111[0:0];
  _RAND_112 = {2{`RANDOM}};
  cycleCnt = _RAND_112[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_T_216 <= 3'h1); // @[src/main/scala/rocket/CSR.scala 1020:9]
    end
    //
    if (_T_220) begin
      assert(1'h1); // @[src/main/scala/rocket/CSR.scala 1028:9]
    end
    //
    if (_T_220) begin
      assert(~reg_singleStepped | ~io_retire); // @[src/main/scala/rocket/CSR.scala 1029:9]
    end
  end
endmodule
module BreakpointUnit(
  input   clock,
  input   reset
);
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_dw, // @[src/main/scala/rocket/ALU.scala 126:14]
  input  [3:0]  io_fn, // @[src/main/scala/rocket/ALU.scala 126:14]
  input  [63:0] io_in2, // @[src/main/scala/rocket/ALU.scala 126:14]
  input  [63:0] io_in1, // @[src/main/scala/rocket/ALU.scala 126:14]
  output [63:0] io_out, // @[src/main/scala/rocket/ALU.scala 126:14]
  output [63:0] io_adder_out, // @[src/main/scala/rocket/ALU.scala 126:14]
  output        io_cmp_out // @[src/main/scala/rocket/ALU.scala 126:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _in2_inv_T_1 = ~io_in2; // @[src/main/scala/rocket/ALU.scala 139:41]
  wire [63:0] in2_inv = io_fn[3] ? _in2_inv_T_1 : io_in2; // @[src/main/scala/rocket/ALU.scala 139:20]
  wire [63:0] in1_xor_in2 = io_in1 ^ in2_inv; // @[src/main/scala/rocket/ALU.scala 140:28]
  wire [63:0] _io_adder_out_T_1 = io_in1 + in2_inv; // @[src/main/scala/rocket/ALU.scala 141:26]
  wire [63:0] _GEN_2 = {{63'd0}, io_fn[3]}; // @[src/main/scala/rocket/ALU.scala 141:36]
  wire  _slt_T_7 = io_fn[1] ? io_in2[63] : io_in1[63]; // @[src/main/scala/rocket/ALU.scala 146:8]
  wire  slt = io_in1[63] == io_in2[63] ? io_adder_out[63] : _slt_T_7; // @[src/main/scala/rocket/ALU.scala 145:8]
  wire  _io_cmp_out_T_2 = ~io_fn[3]; // @[src/main/scala/rocket/ALU.scala 114:26]
  wire  _io_cmp_out_T_4 = _io_cmp_out_T_2 ? in1_xor_in2 == 64'h0 : slt; // @[src/main/scala/rocket/ALU.scala 147:47]
  wire [31:0] shin_hi_32 = io_fn[3] & io_in1[31] ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/ALU.scala 154:28]
  wire [31:0] shin_hi = io_dw ? io_in1[63:32] : shin_hi_32; // @[src/main/scala/rocket/ALU.scala 155:24]
  wire  _shamt_T_2 = io_in2[5] & io_dw; // @[src/main/scala/rocket/ALU.scala 156:33]
  wire [5:0] shamt = {_shamt_T_2,io_in2[4:0]}; // @[src/main/scala/rocket/ALU.scala 156:22]
  wire [63:0] shin_r = {shin_hi,io_in1[31:0]}; // @[src/main/scala/rocket/ALU.scala 157:18]
  wire  _shin_T_2 = io_fn == 4'h5 | io_fn == 4'hb; // @[src/main/scala/rocket/ALU.scala 159:41]
  wire [63:0] _GEN_3 = {{32'd0}, shin_r[63:32]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_6 = _GEN_3 & 64'hffffffff; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_8 = {shin_r[31:0], 32'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_10 = _shin_T_8 & 64'hffffffff00000000; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _GEN_4 = {{16'd0}, _shin_T_11[63:16]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_16 = _GEN_4 & 64'hffff0000ffff; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_18 = {_shin_T_11[47:0], 16'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_20 = _shin_T_18 & 64'hffff0000ffff0000; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _GEN_5 = {{8'd0}, _shin_T_21[63:8]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_26 = _GEN_5 & 64'hff00ff00ff00ff; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_28 = {_shin_T_21[55:0], 8'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_30 = _shin_T_28 & 64'hff00ff00ff00ff00; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _GEN_6 = {{4'd0}, _shin_T_31[63:4]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_36 = _GEN_6 & 64'hf0f0f0f0f0f0f0f; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_38 = {_shin_T_31[59:0], 4'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_40 = _shin_T_38 & 64'hf0f0f0f0f0f0f0f0; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _GEN_7 = {{2'd0}, _shin_T_41[63:2]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_46 = _GEN_7 & 64'h3333333333333333; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_48 = {_shin_T_41[61:0], 2'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_50 = _shin_T_48 & 64'hcccccccccccccccc; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _GEN_8 = {{1'd0}, _shin_T_51[63:1]}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_56 = _GEN_8 & 64'h5555555555555555; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_58 = {_shin_T_51[62:0], 1'h0}; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_60 = _shin_T_58 & 64'haaaaaaaaaaaaaaaa; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] _shin_T_61 = _shin_T_56 | _shin_T_60; // @[src/main/scala/rocket/ALU.scala 159:83]
  wire [63:0] shin = io_fn == 4'h5 | io_fn == 4'hb ? shin_r : _shin_T_61; // @[src/main/scala/rocket/ALU.scala 159:17]
  wire  _shout_r_T_2 = io_fn[3] & shin[63]; // @[src/main/scala/rocket/ALU.scala 160:41]
  wire [64:0] _shout_r_T_4 = {_shout_r_T_2,shin}; // @[src/main/scala/rocket/ALU.scala 160:63]
  wire [64:0] _shout_r_T_5 = $signed(_shout_r_T_4) >>> shamt; // @[src/main/scala/rocket/ALU.scala 160:70]
  wire [63:0] shout_r = _shout_r_T_5[63:0]; // @[src/main/scala/rocket/ALU.scala 160:79]
  wire [63:0] _GEN_9 = {{32'd0}, shout_r[63:32]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_3 = _GEN_9 & 64'hffffffff; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_5 = {shout_r[31:0], 32'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_7 = _shout_l_T_5 & 64'hffffffff00000000; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _GEN_10 = {{16'd0}, _shout_l_T_8[63:16]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_13 = _GEN_10 & 64'hffff0000ffff; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_15 = {_shout_l_T_8[47:0], 16'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_17 = _shout_l_T_15 & 64'hffff0000ffff0000; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _GEN_11 = {{8'd0}, _shout_l_T_18[63:8]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_23 = _GEN_11 & 64'hff00ff00ff00ff; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_25 = {_shout_l_T_18[55:0], 8'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_27 = _shout_l_T_25 & 64'hff00ff00ff00ff00; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _GEN_12 = {{4'd0}, _shout_l_T_28[63:4]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_33 = _GEN_12 & 64'hf0f0f0f0f0f0f0f; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_35 = {_shout_l_T_28[59:0], 4'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_37 = _shout_l_T_35 & 64'hf0f0f0f0f0f0f0f0; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _GEN_13 = {{2'd0}, _shout_l_T_38[63:2]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_43 = _GEN_13 & 64'h3333333333333333; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_45 = {_shout_l_T_38[61:0], 2'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_47 = _shout_l_T_45 & 64'hcccccccccccccccc; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_48 = _shout_l_T_43 | _shout_l_T_47; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _GEN_14 = {{1'd0}, _shout_l_T_48[63:1]}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_53 = _GEN_14 & 64'h5555555555555555; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_55 = {_shout_l_T_48[62:0], 1'h0}; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_l_T_57 = _shout_l_T_55 & 64'haaaaaaaaaaaaaaaa; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] shout_l = _shout_l_T_53 | _shout_l_T_57; // @[src/main/scala/rocket/ALU.scala 161:24]
  wire [63:0] _shout_T_3 = _shin_T_2 ? shout_r : 64'h0; // @[src/main/scala/rocket/ALU.scala 162:18]
  wire [63:0] _shout_T_5 = io_fn == 4'h1 ? shout_l : 64'h0; // @[src/main/scala/rocket/ALU.scala 163:18]
  wire [63:0] shout = _shout_T_3 | _shout_T_5; // @[src/main/scala/rocket/ALU.scala 162:82]
  wire  _logic_T_1 = io_fn == 4'h6; // @[src/main/scala/rocket/ALU.scala 172:51]
  wire [63:0] _logic_T_3 = io_fn == 4'h4 | io_fn == 4'h6 ? in1_xor_in2 : 64'h0; // @[src/main/scala/rocket/ALU.scala 172:18]
  wire [63:0] _logic_T_7 = io_in1 & io_in2; // @[src/main/scala/rocket/ALU.scala 173:75]
  wire [63:0] _logic_T_8 = _logic_T_1 | io_fn == 4'h7 ? _logic_T_7 : 64'h0; // @[src/main/scala/rocket/ALU.scala 173:18]
  wire [63:0] logic_ = _logic_T_3 | _logic_T_8; // @[src/main/scala/rocket/ALU.scala 172:86]
  wire  _shift_logic_T = io_fn >= 4'hc; // @[src/main/scala/rocket/ALU.scala 111:30]
  wire  _shift_logic_T_1 = _shift_logic_T & slt; // @[src/main/scala/rocket/ALU.scala 175:42]
  wire [63:0] _GEN_15 = {{63'd0}, _shift_logic_T_1}; // @[src/main/scala/rocket/ALU.scala 175:50]
  wire [63:0] _shift_logic_T_2 = _GEN_15 | logic_; // @[src/main/scala/rocket/ALU.scala 175:50]
  wire [63:0] shift_logic = _shift_logic_T_2 | shout; // @[src/main/scala/rocket/ALU.scala 175:58]
  wire [63:0] out = io_fn == 4'h0 | io_fn == 4'ha ? io_adder_out : shift_logic; // @[src/main/scala/rocket/ALU.scala 180:16]
  wire  _T_1 = ~io_dw; // @[src/main/scala/rocket/ALU.scala 185:17]
  wire  line_1101_clock;
  wire  line_1101_reset;
  wire  line_1101_valid;
  reg  line_1101_valid_reg;
  wire [31:0] _io_out_T_1 = out[31] ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/ALU.scala 185:48]
  wire [63:0] _io_out_T_3 = {_io_out_T_1,out[31:0]}; // @[src/main/scala/rocket/ALU.scala 185:43]
  GEN_w1_line #(.COVER_INDEX(1101)) line_1101 (
    .clock(line_1101_clock),
    .reset(line_1101_reset),
    .valid(line_1101_valid)
  );
  assign line_1101_clock = clock;
  assign line_1101_reset = reset;
  assign line_1101_valid = _T_1 ^ line_1101_valid_reg;
  assign io_out = ~io_dw ? _io_out_T_3 : out; // @[src/main/scala/rocket/ALU.scala 182:10 185:{28,37}]
  assign io_adder_out = _io_adder_out_T_1 + _GEN_2; // @[src/main/scala/rocket/ALU.scala 141:36]
  assign io_cmp_out = io_fn[0] ^ _io_cmp_out_T_4; // @[src/main/scala/rocket/ALU.scala 147:42]
  always @(posedge clock) begin
    line_1101_valid_reg <= _T_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1101_valid_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input         io_req_valid, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input  [3:0]  io_req_bits_fn, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input         io_req_bits_dw, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input  [63:0] io_req_bits_in1, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input  [63:0] io_req_bits_in2, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input  [4:0]  io_req_bits_tag, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input         io_kill, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  input         io_resp_ready, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  output        io_resp_valid, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  output [63:0] io_resp_bits_data, // @[src/main/scala/rocket/Multiplier.scala 42:14]
  output [4:0]  io_resp_bits_tag // @[src/main/scala/rocket/Multiplier.scala 42:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [159:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/rocket/Multiplier.scala 48:22]
  reg  req_dw; // @[src/main/scala/rocket/Multiplier.scala 50:16]
  reg [4:0] req_tag; // @[src/main/scala/rocket/Multiplier.scala 50:16]
  reg [6:0] count; // @[src/main/scala/rocket/Multiplier.scala 51:18]
  reg  neg_out; // @[src/main/scala/rocket/Multiplier.scala 54:20]
  reg  isHi; // @[src/main/scala/rocket/Multiplier.scala 55:17]
  reg  resHi; // @[src/main/scala/rocket/Multiplier.scala 56:18]
  reg [64:0] divisor; // @[src/main/scala/rocket/Multiplier.scala 57:20]
  reg [129:0] remainder; // @[src/main/scala/rocket/Multiplier.scala 58:22]
  wire [2:0] decoded_plaInput = io_req_bits_fn[2:0]; // @[src/main/scala/chisel3/util/experimental/decode/decoder.scala 39:16 src/main/scala/chisel3/util/pla.scala 77:22]
  wire [2:0] decoded_invInputs = ~decoded_plaInput; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[0]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  _decoded_T = &decoded_andMatrixInput_0; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[2]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  _decoded_T_1 = &decoded_andMatrixInput_0_1; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_2 = decoded_invInputs[1]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [1:0] _decoded_T_2 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_0_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_3 = &_decoded_T_2; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_3 = decoded_plaInput[0]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_0_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_5 = &_decoded_T_4; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_0_4 = decoded_plaInput[1]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  _decoded_T_6 = &decoded_andMatrixInput_0_4; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  decoded_andMatrixInput_1_2 = decoded_plaInput[2]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [1:0] _decoded_T_7 = {decoded_andMatrixInput_0,decoded_andMatrixInput_1_2}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _decoded_T_8 = &_decoded_T_7; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [1:0] _decoded_orMatrixOutputs_T = {_decoded_T_3,_decoded_T_8}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_orMatrixOutputs_T; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _decoded_orMatrixOutputs_T_2 = {_decoded_T,_decoded_T_3}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_orMatrixOutputs_T_2; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _decoded_orMatrixOutputs_T_4 = {_decoded_T_5,_decoded_T_6}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_orMatrixOutputs_T_4; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_1; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [3:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,
    _decoded_orMatrixOutputs_T_3,_decoded_orMatrixOutputs_T_1}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [3:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1
    ],decoded_orMatrixOutputs[0]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire  cmdMul = decoded_invMatrixOutputs[3]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  cmdHi = decoded_invMatrixOutputs[2]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  lhsSigned = decoded_invMatrixOutputs[1]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  rhsSigned = decoded_invMatrixOutputs[0]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  _T_4 = ~io_req_bits_dw; // @[src/main/scala/rocket/Multiplier.scala 75:60]
  wire  _sign_T_2 = _T_4 ? io_req_bits_in1[31] : io_req_bits_in1[63]; // @[src/main/scala/rocket/Multiplier.scala 78:29]
  wire  lhs_sign = lhsSigned & _sign_T_2; // @[src/main/scala/rocket/Multiplier.scala 78:23]
  wire [31:0] _hi_T = lhs_sign ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/Multiplier.scala 79:29]
  wire [31:0] hi = _T_4 ? _hi_T : io_req_bits_in1[63:32]; // @[src/main/scala/rocket/Multiplier.scala 79:17]
  wire [63:0] lhs_in = {hi,io_req_bits_in1[31:0]}; // @[src/main/scala/rocket/Multiplier.scala 80:9]
  wire  _sign_T_5 = _T_4 ? io_req_bits_in2[31] : io_req_bits_in2[63]; // @[src/main/scala/rocket/Multiplier.scala 78:29]
  wire  rhs_sign = rhsSigned & _sign_T_5; // @[src/main/scala/rocket/Multiplier.scala 78:23]
  wire [31:0] _hi_T_2 = rhs_sign ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/Multiplier.scala 79:29]
  wire [31:0] hi_1 = _T_4 ? _hi_T_2 : io_req_bits_in2[63:32]; // @[src/main/scala/rocket/Multiplier.scala 79:17]
  wire [64:0] subtractor = remainder[128:64] - divisor; // @[src/main/scala/rocket/Multiplier.scala 85:37]
  wire [63:0] result = resHi ? remainder[128:65] : remainder[63:0]; // @[src/main/scala/rocket/Multiplier.scala 86:19]
  wire [63:0] negated_remainder = 64'h0 - result; // @[src/main/scala/rocket/Multiplier.scala 87:27]
  wire  _T_10 = state == 3'h1; // @[src/main/scala/rocket/Multiplier.scala 89:39]
  wire  line_1102_clock;
  wire  line_1102_reset;
  wire  line_1102_valid;
  reg  line_1102_valid_reg;
  wire  line_1103_clock;
  wire  line_1103_reset;
  wire  line_1103_valid;
  reg  line_1103_valid_reg;
  wire [129:0] _GEN_12 = remainder[63] ? {{66'd0}, negated_remainder} : remainder; // @[src/main/scala/rocket/Multiplier.scala 90:27 91:17 58:22]
  wire  line_1104_clock;
  wire  line_1104_reset;
  wire  line_1104_valid;
  reg  line_1104_valid_reg;
  wire [129:0] _GEN_14 = state == 3'h1 ? _GEN_12 : remainder; // @[src/main/scala/rocket/Multiplier.scala 58:22 89:57]
  wire [2:0] _GEN_16 = state == 3'h1 ? 3'h3 : state; // @[src/main/scala/rocket/Multiplier.scala 89:57 96:11 48:22]
  wire  _T_13 = state == 3'h5; // @[src/main/scala/rocket/Multiplier.scala 98:39]
  wire  line_1105_clock;
  wire  line_1105_reset;
  wire  line_1105_valid;
  reg  line_1105_valid_reg;
  wire [2:0] _GEN_18 = state == 3'h5 ? 3'h7 : _GEN_16; // @[src/main/scala/rocket/Multiplier.scala 100:11 98:57]
  wire  _GEN_19 = state == 3'h5 ? 1'h0 : resHi; // @[src/main/scala/rocket/Multiplier.scala 101:11 56:18 98:57]
  wire  _T_14 = state == 3'h2; // @[src/main/scala/rocket/Multiplier.scala 103:39]
  wire  line_1106_clock;
  wire  line_1106_reset;
  wire  line_1106_valid;
  reg  line_1106_valid_reg;
  wire [128:0] mulReg = {remainder[129:65],remainder[63:0]}; // @[src/main/scala/rocket/Multiplier.scala 104:21]
  wire  mplierSign = remainder[64]; // @[src/main/scala/rocket/Multiplier.scala 105:31]
  wire [63:0] mplier = mulReg[63:0]; // @[src/main/scala/rocket/Multiplier.scala 106:24]
  wire [64:0] accum = mulReg[128:64]; // @[src/main/scala/rocket/Multiplier.scala 107:37]
  wire [8:0] _prod_T_2 = {mplierSign,mplier[7:0]}; // @[src/main/scala/rocket/Multiplier.scala 109:60]
  wire [73:0] _prod_T_3 = $signed(_prod_T_2) * $signed(divisor); // @[src/main/scala/rocket/Multiplier.scala 109:67]
  wire [73:0] _GEN_49 = {{9{accum[64]}},accum}; // @[src/main/scala/rocket/Multiplier.scala 109:76]
  wire [73:0] nextMulReg_hi = $signed(_prod_T_3) + $signed(_GEN_49); // @[src/main/scala/rocket/Multiplier.scala 110:25]
  wire [129:0] nextMulReg = {nextMulReg_hi,mplier[63:8]}; // @[src/main/scala/rocket/Multiplier.scala 110:25]
  wire  nextMplierSign = count == 7'h6 & neg_out; // @[src/main/scala/rocket/Multiplier.scala 111:61]
  wire [10:0] _eOutMask_T = count * 4'h8; // @[src/main/scala/rocket/Multiplier.scala 113:54]
  wire [64:0] _eOutMask_T_2 = 65'sh10000000000000000 >>> _eOutMask_T[5:0]; // @[src/main/scala/rocket/Multiplier.scala 113:44]
  wire [63:0] eOutMask = _eOutMask_T_2[63:0]; // @[src/main/scala/rocket/Multiplier.scala 113:91]
  wire  _eOut_T_4 = ~isHi; // @[src/main/scala/rocket/Multiplier.scala 115:7]
  wire  _eOut_T_5 = count != 7'h7 & count != 7'h0 & _eOut_T_4; // @[src/main/scala/rocket/Multiplier.scala 114:91]
  wire [63:0] _eOut_T_6 = ~eOutMask; // @[src/main/scala/rocket/Multiplier.scala 115:26]
  wire [63:0] _eOut_T_7 = mplier & _eOut_T_6; // @[src/main/scala/rocket/Multiplier.scala 115:24]
  wire  eOut = _eOut_T_5 & _eOut_T_7 == 64'h0; // @[src/main/scala/rocket/Multiplier.scala 115:13]
  wire [10:0] _eOutRes_T_2 = 11'h40 - _eOutMask_T; // @[src/main/scala/rocket/Multiplier.scala 116:38]
  wire [128:0] eOutRes = mulReg >> _eOutRes_T_2[5:0]; // @[src/main/scala/rocket/Multiplier.scala 116:27]
  wire [129:0] _nextMulReg1_T_1 = eOut ? {{1'd0}, eOutRes} : nextMulReg; // @[src/main/scala/rocket/Multiplier.scala 117:55]
  wire [128:0] nextMulReg1 = {nextMulReg[128:64],_nextMulReg1_T_1[63:0]}; // @[src/main/scala/rocket/Multiplier.scala 117:26]
  wire [129:0] _remainder_T_2 = {nextMulReg1[128:64],nextMplierSign,nextMulReg1[63:0]}; // @[src/main/scala/rocket/Multiplier.scala 118:21]
  wire [6:0] _count_T_1 = count + 7'h1; // @[src/main/scala/rocket/Multiplier.scala 120:20]
  wire  _T_16 = eOut | count == 7'h7; // @[src/main/scala/rocket/Multiplier.scala 121:16]
  wire  line_1107_clock;
  wire  line_1107_reset;
  wire  line_1107_valid;
  reg  line_1107_valid_reg;
  wire [2:0] _GEN_20 = eOut | count == 7'h7 ? 3'h6 : _GEN_18; // @[src/main/scala/rocket/Multiplier.scala 121:55 122:13]
  wire  _GEN_21 = eOut | count == 7'h7 ? isHi : _GEN_19; // @[src/main/scala/rocket/Multiplier.scala 121:55 123:13]
  wire [2:0] _GEN_24 = state == 3'h2 ? _GEN_20 : _GEN_18; // @[src/main/scala/rocket/Multiplier.scala 103:50]
  wire  _GEN_25 = state == 3'h2 ? _GEN_21 : _GEN_19; // @[src/main/scala/rocket/Multiplier.scala 103:50]
  wire  _T_17 = state == 3'h3; // @[src/main/scala/rocket/Multiplier.scala 126:39]
  wire  line_1108_clock;
  wire  line_1108_reset;
  wire  line_1108_valid;
  reg  line_1108_valid_reg;
  wire  unrolls_less = subtractor[64]; // @[src/main/scala/rocket/Multiplier.scala 130:28]
  wire [63:0] _unrolls_T_2 = unrolls_less ? remainder[127:64] : subtractor[63:0]; // @[src/main/scala/rocket/Multiplier.scala 131:14]
  wire  _unrolls_T_4 = ~unrolls_less; // @[src/main/scala/rocket/Multiplier.scala 131:67]
  wire [128:0] unrolls_0 = {_unrolls_T_2,remainder[63:0],_unrolls_T_4}; // @[src/main/scala/rocket/Multiplier.scala 131:10]
  wire  _T_18 = count == 7'h40; // @[src/main/scala/rocket/Multiplier.scala 135:17]
  wire  line_1109_clock;
  wire  line_1109_reset;
  wire  line_1109_valid;
  reg  line_1109_valid_reg;
  wire [2:0] _state_T = neg_out ? 3'h5 : 3'h7; // @[src/main/scala/rocket/Multiplier.scala 136:19]
  wire [2:0] _GEN_26 = count == 7'h40 ? _state_T : _GEN_24; // @[src/main/scala/rocket/Multiplier.scala 135:42 136:13]
  wire  _divby0_T = count == 7'h0; // @[src/main/scala/rocket/Multiplier.scala 143:24]
  wire  divby0 = count == 7'h0 & _unrolls_T_4; // @[src/main/scala/rocket/Multiplier.scala 143:32]
  wire [31:0] divisorMSB_hi = divisor[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] divisorMSB_lo = divisor[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi = |divisorMSB_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] divisorMSB_hi_1 = divisorMSB_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] divisorMSB_lo_1 = divisorMSB_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_1 = |divisorMSB_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] divisorMSB_hi_2 = divisorMSB_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] divisorMSB_lo_2 = divisorMSB_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_2 = |divisorMSB_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] divisorMSB_hi_3 = divisorMSB_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_3 = divisorMSB_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_3 = |divisorMSB_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_4 = divisorMSB_hi_3[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_5 = divisorMSB_hi_3[3] ? 2'h3 : _divisorMSB_T_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_9 = divisorMSB_lo_3[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_10 = divisorMSB_lo_3[3] ? 2'h3 : _divisorMSB_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_11 = divisorMSB_useHi_3 ? _divisorMSB_T_5 : _divisorMSB_T_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_12 = {divisorMSB_useHi_3,_divisorMSB_T_11}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] divisorMSB_hi_4 = divisorMSB_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_4 = divisorMSB_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_4 = |divisorMSB_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_16 = divisorMSB_hi_4[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_17 = divisorMSB_hi_4[3] ? 2'h3 : _divisorMSB_T_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_21 = divisorMSB_lo_4[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_22 = divisorMSB_lo_4[3] ? 2'h3 : _divisorMSB_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_23 = divisorMSB_useHi_4 ? _divisorMSB_T_17 : _divisorMSB_T_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_24 = {divisorMSB_useHi_4,_divisorMSB_T_23}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _divisorMSB_T_25 = divisorMSB_useHi_2 ? _divisorMSB_T_12 : _divisorMSB_T_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _divisorMSB_T_26 = {divisorMSB_useHi_2,_divisorMSB_T_25}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] divisorMSB_hi_5 = divisorMSB_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] divisorMSB_lo_5 = divisorMSB_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_5 = |divisorMSB_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] divisorMSB_hi_6 = divisorMSB_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_6 = divisorMSB_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_6 = |divisorMSB_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_30 = divisorMSB_hi_6[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_31 = divisorMSB_hi_6[3] ? 2'h3 : _divisorMSB_T_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_35 = divisorMSB_lo_6[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_36 = divisorMSB_lo_6[3] ? 2'h3 : _divisorMSB_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_37 = divisorMSB_useHi_6 ? _divisorMSB_T_31 : _divisorMSB_T_36; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_38 = {divisorMSB_useHi_6,_divisorMSB_T_37}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] divisorMSB_hi_7 = divisorMSB_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_7 = divisorMSB_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_7 = |divisorMSB_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_42 = divisorMSB_hi_7[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_43 = divisorMSB_hi_7[3] ? 2'h3 : _divisorMSB_T_42; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_47 = divisorMSB_lo_7[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_48 = divisorMSB_lo_7[3] ? 2'h3 : _divisorMSB_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_49 = divisorMSB_useHi_7 ? _divisorMSB_T_43 : _divisorMSB_T_48; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_50 = {divisorMSB_useHi_7,_divisorMSB_T_49}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _divisorMSB_T_51 = divisorMSB_useHi_5 ? _divisorMSB_T_38 : _divisorMSB_T_50; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _divisorMSB_T_52 = {divisorMSB_useHi_5,_divisorMSB_T_51}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _divisorMSB_T_53 = divisorMSB_useHi_1 ? _divisorMSB_T_26 : _divisorMSB_T_52; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _divisorMSB_T_54 = {divisorMSB_useHi_1,_divisorMSB_T_53}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] divisorMSB_hi_8 = divisorMSB_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] divisorMSB_lo_8 = divisorMSB_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_8 = |divisorMSB_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] divisorMSB_hi_9 = divisorMSB_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] divisorMSB_lo_9 = divisorMSB_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_9 = |divisorMSB_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] divisorMSB_hi_10 = divisorMSB_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_10 = divisorMSB_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_10 = |divisorMSB_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_58 = divisorMSB_hi_10[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_59 = divisorMSB_hi_10[3] ? 2'h3 : _divisorMSB_T_58; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_63 = divisorMSB_lo_10[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_64 = divisorMSB_lo_10[3] ? 2'h3 : _divisorMSB_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_65 = divisorMSB_useHi_10 ? _divisorMSB_T_59 : _divisorMSB_T_64; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_66 = {divisorMSB_useHi_10,_divisorMSB_T_65}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] divisorMSB_hi_11 = divisorMSB_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_11 = divisorMSB_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_11 = |divisorMSB_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_70 = divisorMSB_hi_11[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_71 = divisorMSB_hi_11[3] ? 2'h3 : _divisorMSB_T_70; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_75 = divisorMSB_lo_11[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_76 = divisorMSB_lo_11[3] ? 2'h3 : _divisorMSB_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_77 = divisorMSB_useHi_11 ? _divisorMSB_T_71 : _divisorMSB_T_76; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_78 = {divisorMSB_useHi_11,_divisorMSB_T_77}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _divisorMSB_T_79 = divisorMSB_useHi_9 ? _divisorMSB_T_66 : _divisorMSB_T_78; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _divisorMSB_T_80 = {divisorMSB_useHi_9,_divisorMSB_T_79}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] divisorMSB_hi_12 = divisorMSB_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] divisorMSB_lo_12 = divisorMSB_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_12 = |divisorMSB_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] divisorMSB_hi_13 = divisorMSB_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_13 = divisorMSB_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_13 = |divisorMSB_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_84 = divisorMSB_hi_13[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_85 = divisorMSB_hi_13[3] ? 2'h3 : _divisorMSB_T_84; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_89 = divisorMSB_lo_13[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_90 = divisorMSB_lo_13[3] ? 2'h3 : _divisorMSB_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_91 = divisorMSB_useHi_13 ? _divisorMSB_T_85 : _divisorMSB_T_90; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_92 = {divisorMSB_useHi_13,_divisorMSB_T_91}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] divisorMSB_hi_14 = divisorMSB_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] divisorMSB_lo_14 = divisorMSB_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  divisorMSB_useHi_14 = |divisorMSB_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _divisorMSB_T_96 = divisorMSB_hi_14[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_97 = divisorMSB_hi_14[3] ? 2'h3 : _divisorMSB_T_96; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_101 = divisorMSB_lo_14[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_102 = divisorMSB_lo_14[3] ? 2'h3 : _divisorMSB_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _divisorMSB_T_103 = divisorMSB_useHi_14 ? _divisorMSB_T_97 : _divisorMSB_T_102; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _divisorMSB_T_104 = {divisorMSB_useHi_14,_divisorMSB_T_103}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _divisorMSB_T_105 = divisorMSB_useHi_12 ? _divisorMSB_T_92 : _divisorMSB_T_104; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _divisorMSB_T_106 = {divisorMSB_useHi_12,_divisorMSB_T_105}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _divisorMSB_T_107 = divisorMSB_useHi_8 ? _divisorMSB_T_80 : _divisorMSB_T_106; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _divisorMSB_T_108 = {divisorMSB_useHi_8,_divisorMSB_T_107}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _divisorMSB_T_109 = divisorMSB_useHi ? _divisorMSB_T_54 : _divisorMSB_T_108; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] divisorMSB = {divisorMSB_useHi,_divisorMSB_T_109}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [31:0] dividendMSB_hi = remainder[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] dividendMSB_lo = remainder[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi = |dividendMSB_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] dividendMSB_hi_1 = dividendMSB_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] dividendMSB_lo_1 = dividendMSB_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_1 = |dividendMSB_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] dividendMSB_hi_2 = dividendMSB_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] dividendMSB_lo_2 = dividendMSB_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_2 = |dividendMSB_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] dividendMSB_hi_3 = dividendMSB_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_3 = dividendMSB_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_3 = |dividendMSB_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_4 = dividendMSB_hi_3[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_5 = dividendMSB_hi_3[3] ? 2'h3 : _dividendMSB_T_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_9 = dividendMSB_lo_3[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_10 = dividendMSB_lo_3[3] ? 2'h3 : _dividendMSB_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_11 = dividendMSB_useHi_3 ? _dividendMSB_T_5 : _dividendMSB_T_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_12 = {dividendMSB_useHi_3,_dividendMSB_T_11}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] dividendMSB_hi_4 = dividendMSB_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_4 = dividendMSB_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_4 = |dividendMSB_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_16 = dividendMSB_hi_4[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_17 = dividendMSB_hi_4[3] ? 2'h3 : _dividendMSB_T_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_21 = dividendMSB_lo_4[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_22 = dividendMSB_lo_4[3] ? 2'h3 : _dividendMSB_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_23 = dividendMSB_useHi_4 ? _dividendMSB_T_17 : _dividendMSB_T_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_24 = {dividendMSB_useHi_4,_dividendMSB_T_23}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _dividendMSB_T_25 = dividendMSB_useHi_2 ? _dividendMSB_T_12 : _dividendMSB_T_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _dividendMSB_T_26 = {dividendMSB_useHi_2,_dividendMSB_T_25}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] dividendMSB_hi_5 = dividendMSB_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] dividendMSB_lo_5 = dividendMSB_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_5 = |dividendMSB_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] dividendMSB_hi_6 = dividendMSB_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_6 = dividendMSB_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_6 = |dividendMSB_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_30 = dividendMSB_hi_6[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_31 = dividendMSB_hi_6[3] ? 2'h3 : _dividendMSB_T_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_35 = dividendMSB_lo_6[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_36 = dividendMSB_lo_6[3] ? 2'h3 : _dividendMSB_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_37 = dividendMSB_useHi_6 ? _dividendMSB_T_31 : _dividendMSB_T_36; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_38 = {dividendMSB_useHi_6,_dividendMSB_T_37}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] dividendMSB_hi_7 = dividendMSB_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_7 = dividendMSB_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_7 = |dividendMSB_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_42 = dividendMSB_hi_7[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_43 = dividendMSB_hi_7[3] ? 2'h3 : _dividendMSB_T_42; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_47 = dividendMSB_lo_7[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_48 = dividendMSB_lo_7[3] ? 2'h3 : _dividendMSB_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_49 = dividendMSB_useHi_7 ? _dividendMSB_T_43 : _dividendMSB_T_48; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_50 = {dividendMSB_useHi_7,_dividendMSB_T_49}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _dividendMSB_T_51 = dividendMSB_useHi_5 ? _dividendMSB_T_38 : _dividendMSB_T_50; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _dividendMSB_T_52 = {dividendMSB_useHi_5,_dividendMSB_T_51}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _dividendMSB_T_53 = dividendMSB_useHi_1 ? _dividendMSB_T_26 : _dividendMSB_T_52; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _dividendMSB_T_54 = {dividendMSB_useHi_1,_dividendMSB_T_53}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] dividendMSB_hi_8 = dividendMSB_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] dividendMSB_lo_8 = dividendMSB_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_8 = |dividendMSB_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] dividendMSB_hi_9 = dividendMSB_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] dividendMSB_lo_9 = dividendMSB_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_9 = |dividendMSB_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] dividendMSB_hi_10 = dividendMSB_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_10 = dividendMSB_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_10 = |dividendMSB_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_58 = dividendMSB_hi_10[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_59 = dividendMSB_hi_10[3] ? 2'h3 : _dividendMSB_T_58; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_63 = dividendMSB_lo_10[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_64 = dividendMSB_lo_10[3] ? 2'h3 : _dividendMSB_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_65 = dividendMSB_useHi_10 ? _dividendMSB_T_59 : _dividendMSB_T_64; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_66 = {dividendMSB_useHi_10,_dividendMSB_T_65}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] dividendMSB_hi_11 = dividendMSB_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_11 = dividendMSB_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_11 = |dividendMSB_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_70 = dividendMSB_hi_11[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_71 = dividendMSB_hi_11[3] ? 2'h3 : _dividendMSB_T_70; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_75 = dividendMSB_lo_11[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_76 = dividendMSB_lo_11[3] ? 2'h3 : _dividendMSB_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_77 = dividendMSB_useHi_11 ? _dividendMSB_T_71 : _dividendMSB_T_76; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_78 = {dividendMSB_useHi_11,_dividendMSB_T_77}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _dividendMSB_T_79 = dividendMSB_useHi_9 ? _dividendMSB_T_66 : _dividendMSB_T_78; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _dividendMSB_T_80 = {dividendMSB_useHi_9,_dividendMSB_T_79}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] dividendMSB_hi_12 = dividendMSB_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] dividendMSB_lo_12 = dividendMSB_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_12 = |dividendMSB_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] dividendMSB_hi_13 = dividendMSB_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_13 = dividendMSB_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_13 = |dividendMSB_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_84 = dividendMSB_hi_13[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_85 = dividendMSB_hi_13[3] ? 2'h3 : _dividendMSB_T_84; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_89 = dividendMSB_lo_13[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_90 = dividendMSB_lo_13[3] ? 2'h3 : _dividendMSB_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_91 = dividendMSB_useHi_13 ? _dividendMSB_T_85 : _dividendMSB_T_90; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_92 = {dividendMSB_useHi_13,_dividendMSB_T_91}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] dividendMSB_hi_14 = dividendMSB_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] dividendMSB_lo_14 = dividendMSB_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  dividendMSB_useHi_14 = |dividendMSB_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _dividendMSB_T_96 = dividendMSB_hi_14[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_97 = dividendMSB_hi_14[3] ? 2'h3 : _dividendMSB_T_96; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_101 = dividendMSB_lo_14[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_102 = dividendMSB_lo_14[3] ? 2'h3 : _dividendMSB_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _dividendMSB_T_103 = dividendMSB_useHi_14 ? _dividendMSB_T_97 : _dividendMSB_T_102; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _dividendMSB_T_104 = {dividendMSB_useHi_14,_dividendMSB_T_103}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _dividendMSB_T_105 = dividendMSB_useHi_12 ? _dividendMSB_T_92 : _dividendMSB_T_104; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _dividendMSB_T_106 = {dividendMSB_useHi_12,_dividendMSB_T_105}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _dividendMSB_T_107 = dividendMSB_useHi_8 ? _dividendMSB_T_80 : _dividendMSB_T_106; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _dividendMSB_T_108 = {dividendMSB_useHi_8,_dividendMSB_T_107}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _dividendMSB_T_109 = dividendMSB_useHi ? _dividendMSB_T_54 : _dividendMSB_T_108; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] dividendMSB = {dividendMSB_useHi,_dividendMSB_T_109}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _eOutPos_T_1 = dividendMSB - divisorMSB; // @[src/main/scala/rocket/Multiplier.scala 149:35]
  wire [5:0] eOutPos = ~_eOutPos_T_1; // @[src/main/scala/rocket/Multiplier.scala 149:21]
  wire  eOut_1 = _divby0_T & ~divby0 & eOutPos >= 6'h1; // @[src/main/scala/rocket/Multiplier.scala 150:43]
  wire  line_1110_clock;
  wire  line_1110_reset;
  wire  line_1110_valid;
  reg  line_1110_valid_reg;
  wire [126:0] _GEN_38 = {{63'd0}, remainder[63:0]}; // @[src/main/scala/rocket/Multiplier.scala 152:39]
  wire [126:0] _remainder_T_4 = _GEN_38 << eOutPos; // @[src/main/scala/rocket/Multiplier.scala 152:39]
  wire [128:0] _GEN_28 = eOut_1 ? {{2'd0}, _remainder_T_4} : unrolls_0; // @[src/main/scala/rocket/Multiplier.scala 134:15 151:19 152:19]
  wire  _T_20 = divby0 & _eOut_T_4; // @[src/main/scala/rocket/Multiplier.scala 156:18]
  wire  line_1111_clock;
  wire  line_1111_reset;
  wire  line_1111_valid;
  reg  line_1111_valid_reg;
  wire  _T_21 = io_resp_ready & io_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_22 = _T_21 | io_kill; // @[src/main/scala/rocket/Multiplier.scala 158:22]
  wire  line_1112_clock;
  wire  line_1112_reset;
  wire  line_1112_valid;
  reg  line_1112_valid_reg;
  wire  _T_23 = io_req_ready & io_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1113_clock;
  wire  line_1113_reset;
  wire  line_1113_valid;
  reg  line_1113_valid_reg;
  wire [2:0] _count_T_8 = cmdMul & _T_4 ? 3'h4 : 3'h0; // @[src/main/scala/rocket/Multiplier.scala 165:38]
  wire [64:0] _divisor_T = {rhs_sign,hi_1,io_req_bits_in2[31:0]}; // @[src/main/scala/rocket/Multiplier.scala 167:19]
  wire [2:0] _outMul_T_1 = state & 3'h1; // @[src/main/scala/rocket/Multiplier.scala 172:23]
  wire  outMul = _outMul_T_1 == 3'h0; // @[src/main/scala/rocket/Multiplier.scala 172:52]
  wire  _loOut_T = ~req_dw; // @[src/main/scala/rocket/Multiplier.scala 75:60]
  wire [31:0] loOut = _loOut_T & outMul ? result[63:32] : result[31:0]; // @[src/main/scala/rocket/Multiplier.scala 173:18]
  wire [31:0] _hiOut_T_3 = loOut[31] ? 32'hffffffff : 32'h0; // @[src/main/scala/rocket/Multiplier.scala 174:39]
  wire [31:0] hiOut = _loOut_T ? _hiOut_T_3 : result[63:32]; // @[src/main/scala/rocket/Multiplier.scala 174:18]
  GEN_w1_line #(.COVER_INDEX(1102)) line_1102 (
    .clock(line_1102_clock),
    .reset(line_1102_reset),
    .valid(line_1102_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1103)) line_1103 (
    .clock(line_1103_clock),
    .reset(line_1103_reset),
    .valid(line_1103_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1104)) line_1104 (
    .clock(line_1104_clock),
    .reset(line_1104_reset),
    .valid(line_1104_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1105)) line_1105 (
    .clock(line_1105_clock),
    .reset(line_1105_reset),
    .valid(line_1105_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1106)) line_1106 (
    .clock(line_1106_clock),
    .reset(line_1106_reset),
    .valid(line_1106_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1107)) line_1107 (
    .clock(line_1107_clock),
    .reset(line_1107_reset),
    .valid(line_1107_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1108)) line_1108 (
    .clock(line_1108_clock),
    .reset(line_1108_reset),
    .valid(line_1108_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1109)) line_1109 (
    .clock(line_1109_clock),
    .reset(line_1109_reset),
    .valid(line_1109_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1110)) line_1110 (
    .clock(line_1110_clock),
    .reset(line_1110_reset),
    .valid(line_1110_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1111)) line_1111 (
    .clock(line_1111_clock),
    .reset(line_1111_reset),
    .valid(line_1111_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1112)) line_1112 (
    .clock(line_1112_clock),
    .reset(line_1112_reset),
    .valid(line_1112_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1113)) line_1113 (
    .clock(line_1113_clock),
    .reset(line_1113_reset),
    .valid(line_1113_valid)
  );
  assign line_1102_clock = clock;
  assign line_1102_reset = reset;
  assign line_1102_valid = _T_10 ^ line_1102_valid_reg;
  assign line_1103_clock = clock;
  assign line_1103_reset = reset;
  assign line_1103_valid = remainder[63] ^ line_1103_valid_reg;
  assign line_1104_clock = clock;
  assign line_1104_reset = reset;
  assign line_1104_valid = divisor[63] ^ line_1104_valid_reg;
  assign line_1105_clock = clock;
  assign line_1105_reset = reset;
  assign line_1105_valid = _T_13 ^ line_1105_valid_reg;
  assign line_1106_clock = clock;
  assign line_1106_reset = reset;
  assign line_1106_valid = _T_14 ^ line_1106_valid_reg;
  assign line_1107_clock = clock;
  assign line_1107_reset = reset;
  assign line_1107_valid = _T_16 ^ line_1107_valid_reg;
  assign line_1108_clock = clock;
  assign line_1108_reset = reset;
  assign line_1108_valid = _T_17 ^ line_1108_valid_reg;
  assign line_1109_clock = clock;
  assign line_1109_reset = reset;
  assign line_1109_valid = _T_18 ^ line_1109_valid_reg;
  assign line_1110_clock = clock;
  assign line_1110_reset = reset;
  assign line_1110_valid = eOut_1 ^ line_1110_valid_reg;
  assign line_1111_clock = clock;
  assign line_1111_reset = reset;
  assign line_1111_valid = _T_20 ^ line_1111_valid_reg;
  assign line_1112_clock = clock;
  assign line_1112_reset = reset;
  assign line_1112_valid = _T_22 ^ line_1112_valid_reg;
  assign line_1113_clock = clock;
  assign line_1113_reset = reset;
  assign line_1113_valid = _T_23 ^ line_1113_valid_reg;
  assign io_req_ready = state == 3'h0; // @[src/main/scala/rocket/Multiplier.scala 179:25]
  assign io_resp_valid = state == 3'h6 | state == 3'h7; // @[src/main/scala/rocket/Multiplier.scala 178:42]
  assign io_resp_bits_data = {hiOut,loOut}; // @[src/main/scala/rocket/Multiplier.scala 177:27]
  assign io_resp_bits_tag = req_tag; // @[src/main/scala/rocket/Multiplier.scala 175:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/rocket/Multiplier.scala 48:22]
      state <= 3'h0; // @[src/main/scala/rocket/Multiplier.scala 48:22]
    end else if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      if (cmdMul) begin // @[src/main/scala/rocket/Multiplier.scala 162:17]
        state <= 3'h2;
      end else if (lhs_sign | rhs_sign) begin // @[src/main/scala/rocket/Multiplier.scala 162:36]
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (_T_21 | io_kill) begin // @[src/main/scala/rocket/Multiplier.scala 158:34]
      state <= 3'h0; // @[src/main/scala/rocket/Multiplier.scala 159:11]
    end else if (state == 3'h3) begin // @[src/main/scala/rocket/Multiplier.scala 126:50]
      state <= _GEN_26;
    end else begin
      state <= _GEN_24;
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      req_dw <= io_req_bits_dw; // @[src/main/scala/rocket/Multiplier.scala 169:9]
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      req_tag <= io_req_bits_tag; // @[src/main/scala/rocket/Multiplier.scala 169:9]
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      count <= {{4'd0}, _count_T_8}; // @[src/main/scala/rocket/Multiplier.scala 165:11]
    end else if (state == 3'h3) begin // @[src/main/scala/rocket/Multiplier.scala 126:50]
      if (eOut_1) begin // @[src/main/scala/rocket/Multiplier.scala 151:19]
        count <= {{1'd0}, eOutPos}; // @[src/main/scala/rocket/Multiplier.scala 153:15]
      end else begin
        count <= _count_T_1; // @[src/main/scala/rocket/Multiplier.scala 141:11]
      end
    end else if (state == 3'h2) begin // @[src/main/scala/rocket/Multiplier.scala 103:50]
      count <= _count_T_1; // @[src/main/scala/rocket/Multiplier.scala 120:11]
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      if (cmdHi) begin // @[src/main/scala/rocket/Multiplier.scala 166:19]
        neg_out <= lhs_sign;
      end else begin
        neg_out <= lhs_sign != rhs_sign;
      end
    end else if (state == 3'h3) begin // @[src/main/scala/rocket/Multiplier.scala 126:50]
      if (divby0 & _eOut_T_4) begin // @[src/main/scala/rocket/Multiplier.scala 156:28]
        neg_out <= 1'h0; // @[src/main/scala/rocket/Multiplier.scala 156:38]
      end
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      isHi <= cmdHi; // @[src/main/scala/rocket/Multiplier.scala 163:10]
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      resHi <= 1'h0; // @[src/main/scala/rocket/Multiplier.scala 164:11]
    end else if (state == 3'h3) begin // @[src/main/scala/rocket/Multiplier.scala 126:50]
      if (count == 7'h40) begin // @[src/main/scala/rocket/Multiplier.scala 135:42]
        resHi <= isHi; // @[src/main/scala/rocket/Multiplier.scala 137:13]
      end else begin
        resHi <= _GEN_25;
      end
    end else begin
      resHi <= _GEN_25;
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      divisor <= _divisor_T; // @[src/main/scala/rocket/Multiplier.scala 167:13]
    end else if (state == 3'h1) begin // @[src/main/scala/rocket/Multiplier.scala 89:57]
      if (divisor[63]) begin // @[src/main/scala/rocket/Multiplier.scala 93:25]
        divisor <= subtractor; // @[src/main/scala/rocket/Multiplier.scala 94:15]
      end
    end
    if (_T_23) begin // @[src/main/scala/rocket/Multiplier.scala 161:22]
      remainder <= {{66'd0}, lhs_in}; // @[src/main/scala/rocket/Multiplier.scala 168:15]
    end else if (state == 3'h3) begin // @[src/main/scala/rocket/Multiplier.scala 126:50]
      remainder <= {{1'd0}, _GEN_28};
    end else if (state == 3'h2) begin // @[src/main/scala/rocket/Multiplier.scala 103:50]
      remainder <= _remainder_T_2; // @[src/main/scala/rocket/Multiplier.scala 118:15]
    end else if (state == 3'h5) begin // @[src/main/scala/rocket/Multiplier.scala 98:57]
      remainder <= {{66'd0}, negated_remainder}; // @[src/main/scala/rocket/Multiplier.scala 99:15]
    end else begin
      remainder <= _GEN_14;
    end
    line_1102_valid_reg <= _T_10;
    line_1103_valid_reg <= remainder[63];
    line_1104_valid_reg <= divisor[63];
    line_1105_valid_reg <= _T_13;
    line_1106_valid_reg <= _T_14;
    line_1107_valid_reg <= _T_16;
    line_1108_valid_reg <= _T_17;
    line_1109_valid_reg <= _T_18;
    line_1110_valid_reg <= eOut_1;
    line_1111_valid_reg <= _T_20;
    line_1112_valid_reg <= _T_22;
    line_1113_valid_reg <= _T_23;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  req_tag = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  neg_out = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isHi = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  resHi = _RAND_6[0:0];
  _RAND_7 = {3{`RANDOM}};
  divisor = _RAND_7[64:0];
  _RAND_8 = {5{`RANDOM}};
  remainder = _RAND_8[129:0];
  _RAND_9 = {1{`RANDOM}};
  line_1102_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1103_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1104_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1105_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1106_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1107_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1108_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1109_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1110_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1111_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1112_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  line_1113_valid_reg = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_4(
  input         clock,
  input         reset,
  input  [63:0] io_bits_value_1, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_2, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_3, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_4, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_5, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_6, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_7, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_8, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_9, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_10, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_11, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_12, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_13, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_14, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_15, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_16, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_17, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_18, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_19, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_20, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_21, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_22, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_23, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_24, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_25, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_26, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_27, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_28, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_29, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_30, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_31 // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_0; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_1; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_2; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_3; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_4; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_5; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_6; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_7; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_8; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_9; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_10; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_11; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_12; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_13; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_14; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_15; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_16; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_17; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_18; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_19; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_20; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_21; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_22; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_23; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_24; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_25; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_26; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_27; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_28; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_29; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_30; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_31; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchIntRegState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_value_0(dpic_io_value_0),
    .io_value_1(dpic_io_value_1),
    .io_value_2(dpic_io_value_2),
    .io_value_3(dpic_io_value_3),
    .io_value_4(dpic_io_value_4),
    .io_value_5(dpic_io_value_5),
    .io_value_6(dpic_io_value_6),
    .io_value_7(dpic_io_value_7),
    .io_value_8(dpic_io_value_8),
    .io_value_9(dpic_io_value_9),
    .io_value_10(dpic_io_value_10),
    .io_value_11(dpic_io_value_11),
    .io_value_12(dpic_io_value_12),
    .io_value_13(dpic_io_value_13),
    .io_value_14(dpic_io_value_14),
    .io_value_15(dpic_io_value_15),
    .io_value_16(dpic_io_value_16),
    .io_value_17(dpic_io_value_17),
    .io_value_18(dpic_io_value_18),
    .io_value_19(dpic_io_value_19),
    .io_value_20(dpic_io_value_20),
    .io_value_21(dpic_io_value_21),
    .io_value_22(dpic_io_value_22),
    .io_value_23(dpic_io_value_23),
    .io_value_24(dpic_io_value_24),
    .io_value_25(dpic_io_value_25),
    .io_value_26(dpic_io_value_26),
    .io_value_27(dpic_io_value_27),
    .io_value_28(dpic_io_value_28),
    .io_value_29(dpic_io_value_29),
    .io_value_30(dpic_io_value_30),
    .io_value_31(dpic_io_value_31),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_value_0 = 64'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_1 = io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_2 = io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_3 = io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_4 = io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_5 = io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_6 = io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_7 = io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_8 = io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_9 = io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_10 = io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_11 = io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_12 = io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_13 = io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_14 = io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_15 = io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_16 = io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_17 = io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_18 = io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_19 = io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_20 = io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_21 = io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_22 = io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_23 = io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_24 = io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_25 = io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_26 = io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_27 = io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_28 = io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_29 = io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_30 = io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_31 = io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_5(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_address, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_address; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestIntWriteback dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_address(dpic_io_address),
    .io_data(dpic_io_data),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_address = io_bits_address; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_6(
  input         clock,
  input         reset,
  input  [63:0] io_bits_privilegeMode, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mcause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_scause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_satp, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mie, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mideleg, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_medeleg // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mcause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_scause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_satp; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mie; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mideleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_medeleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestCSRState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_privilegeMode(dpic_io_privilegeMode),
    .io_mstatus(dpic_io_mstatus),
    .io_sstatus(dpic_io_sstatus),
    .io_mepc(dpic_io_mepc),
    .io_sepc(dpic_io_sepc),
    .io_mtval(dpic_io_mtval),
    .io_stval(dpic_io_stval),
    .io_mtvec(dpic_io_mtvec),
    .io_stvec(dpic_io_stvec),
    .io_mcause(dpic_io_mcause),
    .io_scause(dpic_io_scause),
    .io_satp(dpic_io_satp),
    .io_mip(dpic_io_mip),
    .io_mie(dpic_io_mie),
    .io_mscratch(dpic_io_mscratch),
    .io_sscratch(dpic_io_sscratch),
    .io_mideleg(dpic_io_mideleg),
    .io_medeleg(dpic_io_medeleg),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_privilegeMode = io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mstatus = io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sstatus = io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mepc = io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sepc = io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtval = io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stval = io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtvec = io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stvec = io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mcause = io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_scause = io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_satp = io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mip = io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mie = io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mscratch = io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sscratch = io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mideleg = io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_medeleg = io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_7(
  input         clock,
  input         reset,
  input  [63:0] io_bits_minstret, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mcycle // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_minstret; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mcycle; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestSnapshotCSRState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_minstret(dpic_io_minstret),
    .io_mcycle(dpic_io_mcycle),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_minstret = io_bits_minstret; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mcycle = io_bits_mcycle; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DelayReg_3(
  input         clock,
  input         reset,
  input         i_valid, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input         i_skip, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input         i_rfwen, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input         i_fpwen, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [4:0]  i_wpdest, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [7:0]  i_wdest, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [63:0] i_pc, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [31:0] i_instr, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [7:0]  i_special, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  output        o_valid, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output        o_skip, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output        o_rfwen, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output        o_fpwen, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [4:0]  o_wpdest, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [7:0]  o_wdest, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [63:0] o_pc, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [31:0] o_instr, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [7:0]  o_special // @[difftest/src/main/scala/util/Delayer.scala 24:13]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_skip; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_rfwen; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_fpwen; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [4:0] REG_wpdest; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [7:0] REG_wdest; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_pc; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [31:0] REG_instr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [7:0] REG_special; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  assign o_valid = REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_skip = REG_skip; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_rfwen = REG_rfwen; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_fpwen = REG_fpwen; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_wpdest = REG_wpdest; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_wdest = REG_wdest; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_pc = REG_pc; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_instr = REG_instr; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_special = REG_special; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_valid <= i_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_skip <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_skip <= i_skip; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_rfwen <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_rfwen <= i_rfwen; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_fpwen <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_fpwen <= i_fpwen; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_wpdest <= 5'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_wpdest <= i_wpdest; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_wdest <= 8'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_wdest <= i_wdest; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_pc <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_pc <= i_pc; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_instr <= 32'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_instr <= i_instr; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_special <= 8'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_special <= i_special; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_skip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_rfwen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_fpwen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_wpdest = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  REG_wdest = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  REG_pc = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  REG_instr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  REG_special = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_8(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_skip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_rfwen, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_fpwen, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_wpdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_wdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_instr, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_special // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_skip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isRVC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_rfwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_fpwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_vecwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_wpdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_wdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_instr; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [9:0] dpic_io_robIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_lqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_sqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isLoad; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isStore; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_nFused; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_special; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestInstrCommit dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_skip(dpic_io_skip),
    .io_isRVC(dpic_io_isRVC),
    .io_rfwen(dpic_io_rfwen),
    .io_fpwen(dpic_io_fpwen),
    .io_vecwen(dpic_io_vecwen),
    .io_wpdest(dpic_io_wpdest),
    .io_wdest(dpic_io_wdest),
    .io_pc(dpic_io_pc),
    .io_instr(dpic_io_instr),
    .io_robIdx(dpic_io_robIdx),
    .io_lqIdx(dpic_io_lqIdx),
    .io_sqIdx(dpic_io_sqIdx),
    .io_isLoad(dpic_io_isLoad),
    .io_isStore(dpic_io_isStore),
    .io_nFused(dpic_io_nFused),
    .io_special(dpic_io_special),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_skip = io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isRVC = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_rfwen = io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_fpwen = io_bits_fpwen; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_vecwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wpdest = io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wdest = io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instr = io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_robIdx = 10'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_lqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isLoad = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isStore = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_nFused = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_special = io_bits_special; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DelayReg_4(
  input         clock,
  input         reset,
  input         i_valid, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [4:0]  i_address, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input  [63:0] i_data, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  input         i_nack, // @[difftest/src/main/scala/util/Delayer.scala 23:13]
  output        o_valid, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [4:0]  o_address, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output [63:0] o_data, // @[difftest/src/main/scala/util/Delayer.scala 24:13]
  output        o_nack // @[difftest/src/main/scala/util/Delayer.scala 24:13]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [4:0] REG_address; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg [63:0] REG_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  reg  REG_nack; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
  assign o_valid = REG_valid; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_address = REG_address; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_data = REG_data; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  assign o_nack = REG_nack; // @[difftest/src/main/scala/util/Delayer.scala 32:5]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_valid <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_valid <= i_valid; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_address <= 5'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_address <= i_address; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_data <= 64'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_data <= i_data; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
    if (reset) begin // @[difftest/src/main/scala/util/Delayer.scala 30:16]
      REG_nack <= 1'h0; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end else begin
      REG_nack <= i_nack; // @[difftest/src/main/scala/util/Delayer.scala 30:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_address = _RAND_1[4:0];
  _RAND_2 = {2{`RANDOM}};
  REG_data = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  REG_nack = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_9(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_address, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_nack // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_address; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_nack; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchIntDelayedUpdate dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_address(dpic_io_address),
    .io_data(dpic_io_data),
    .io_nack(dpic_io_nack),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_address = io_bits_address; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_nack = io_bits_nack; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module PlusArgTimeout(
  input         clock,
  input         reset,
  input  [31:0] io_count // @[src/main/scala/util/PlusArg.scala 59:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[src/main/scala/util/PlusArg.scala 62:19]
  wire  _T = plusarg_reader_out > 32'h0; // @[src/main/scala/util/PlusArg.scala 63:13]
  wire  line_1114_clock;
  wire  line_1114_reset;
  wire  line_1114_valid;
  reg  line_1114_valid_reg;
  wire  _T_3 = ~reset; // @[src/main/scala/util/PlusArg.scala 64:12]
  wire  line_1115_clock;
  wire  line_1115_reset;
  wire  line_1115_valid;
  reg  line_1115_valid_reg;
  wire  _T_4 = ~(io_count < plusarg_reader_out); // @[src/main/scala/util/PlusArg.scala 64:12]
  wire  line_1116_clock;
  wire  line_1116_reset;
  wire  line_1116_valid;
  reg  line_1116_valid_reg;
  plusarg_reader #(.DEFAULT(0), .FORMAT("max_core_cycles=%d"), .WIDTH(32)) plusarg_reader ( // @[src/main/scala/util/PlusArg.scala 62:19]
    .out(plusarg_reader_out)
  );
  GEN_w1_line #(.COVER_INDEX(1114)) line_1114 (
    .clock(line_1114_clock),
    .reset(line_1114_reset),
    .valid(line_1114_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1115)) line_1115 (
    .clock(line_1115_clock),
    .reset(line_1115_reset),
    .valid(line_1115_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1116)) line_1116 (
    .clock(line_1116_clock),
    .reset(line_1116_reset),
    .valid(line_1116_valid)
  );
  assign line_1114_clock = clock;
  assign line_1114_reset = reset;
  assign line_1114_valid = _T ^ line_1114_valid_reg;
  assign line_1115_clock = clock;
  assign line_1115_reset = reset;
  assign line_1115_valid = _T_3 ^ line_1115_valid_reg;
  assign line_1116_clock = clock;
  assign line_1116_reset = reset;
  assign line_1116_valid = _T_4 ^ line_1116_valid_reg;
  always @(posedge clock) begin
    line_1114_valid_reg <= _T;
    line_1115_valid_reg <= _T_3;
    line_1116_valid_reg <= _T_4;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~reset & ~(io_count < plusarg_reader_out)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n"
            ); // @[src/main/scala/util/PlusArg.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1114_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1115_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1116_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & ~reset) begin
      assert(io_count < plusarg_reader_out); // @[src/main/scala/util/PlusArg.scala 64:12]
    end
  end
endmodule
module Rocket(
  input         clock,
  input         reset,
  input         io_hartid, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_might_request, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_req_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output [39:0] io_imem_req_bits_pc, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_req_bits_speculative, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_sfence_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_sfence_bits_rs1, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_sfence_bits_rs2, // @[src/main/scala/tile/Core.scala 162:14]
  output [38:0] io_imem_sfence_bits_addr, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_resp_ready, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_imem_resp_valid, // @[src/main/scala/tile/Core.scala 162:14]
  input  [39:0] io_imem_resp_bits_pc, // @[src/main/scala/tile/Core.scala 162:14]
  input  [31:0] io_imem_resp_bits_data, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_imem_resp_bits_xcpt_pf_inst, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_imem_resp_bits_xcpt_ae_inst, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_imem_resp_bits_replay, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_btb_update_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_bht_update_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_flush_icache, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_imem_progress, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_req_ready, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_dmem_req_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output [39:0] io_dmem_req_bits_addr, // @[src/main/scala/tile/Core.scala 162:14]
  output [6:0]  io_dmem_req_bits_tag, // @[src/main/scala/tile/Core.scala 162:14]
  output [4:0]  io_dmem_req_bits_cmd, // @[src/main/scala/tile/Core.scala 162:14]
  output [1:0]  io_dmem_req_bits_size, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_dmem_req_bits_signed, // @[src/main/scala/tile/Core.scala 162:14]
  output [1:0]  io_dmem_req_bits_dprv, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_dmem_req_bits_dv, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_dmem_s1_kill, // @[src/main/scala/tile/Core.scala 162:14]
  output [63:0] io_dmem_s1_data_data, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_nack, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_resp_valid, // @[src/main/scala/tile/Core.scala 162:14]
  input  [6:0]  io_dmem_resp_bits_tag, // @[src/main/scala/tile/Core.scala 162:14]
  input  [63:0] io_dmem_resp_bits_data, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_resp_bits_replay, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_resp_bits_has_data, // @[src/main/scala/tile/Core.scala 162:14]
  input  [63:0] io_dmem_resp_bits_data_word_bypass, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_replay_next, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_ma_ld, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_ma_st, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_pf_ld, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_pf_st, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_ae_ld, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_s2_xcpt_ae_st, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_ordered, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_perf_release, // @[src/main/scala/tile/Core.scala 162:14]
  input         io_dmem_perf_grant, // @[src/main/scala/tile/Core.scala 162:14]
  output [3:0]  io_ptw_ptbr_mode, // @[src/main/scala/tile/Core.scala 162:14]
  output [43:0] io_ptw_ptbr_ppn, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_ptw_sfence_valid, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_ptw_sfence_bits_rs1, // @[src/main/scala/tile/Core.scala 162:14]
  output [1:0]  io_ptw_status_prv, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_ptw_status_mxr, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_ptw_status_sum, // @[src/main/scala/tile/Core.scala 162:14]
  output        io_rocc_cmd_valid // @[src/main/scala/tile/Core.scala 162:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
`endif // RANDOMIZE_REG_INIT
  wire  ibuf_clock; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_reset; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_imem_ready; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_imem_valid; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [39:0] ibuf_io_imem_bits_pc; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [31:0] ibuf_io_imem_bits_data; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_imem_bits_xcpt_pf_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_imem_bits_xcpt_ae_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_imem_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_kill; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [39:0] ibuf_io_pc; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_ready; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_valid; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_xcpt1_gf_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  ibuf_io_inst_0_bits_rvc; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [31:0] ibuf_io_inst_0_bits_inst_bits; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rd; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire [31:0] ibuf_io_inst_0_bits_raw; // @[src/main/scala/rocket/RocketCore.scala 284:20]
  wire  csr_clock; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_reset; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_ungated_clock; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_hartid; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [11:0] csr_io_rw_addr; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [2:0] csr_io_rw_cmd; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_rw_rdata; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_rw_wdata; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [31:0] csr_io_decode_0_inst; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_fp_illegal; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_fp_csr; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_rocc_illegal; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_read_illegal; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_write_illegal; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_write_flush; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_decode_0_system_illegal; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_csr_stall; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_rw_stall; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_eret; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_singleStep; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_debug; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_cease; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_wfi; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [31:0] csr_io_status_isa; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_dprv; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_dv; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_prv; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_v; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_sd; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [22:0] csr_io_status_zero2; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mpv; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_gva; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mbe; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_sbe; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_sxl; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_uxl; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_sd_rv32; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [7:0] csr_io_status_zero1; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_tsr; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_tw; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_tvm; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mxr; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_sum; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mprv; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_xs; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_fs; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_mpp; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [1:0] csr_io_status_vs; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_spp; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mpie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_ube; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_spie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_upie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_mie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_hie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_sie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_status_uie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [3:0] csr_io_ptbr_mode; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [43:0] csr_io_ptbr_ppn; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [39:0] csr_io_evec; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_exception; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_retire; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_cause; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [39:0] csr_io_pc; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [39:0] csr_io_tval; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_gva; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_time; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_interrupt; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_interrupt_cause; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_csrr_counter; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [31:0] csr_io_inst_0; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_trace_0_valid; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [39:0] csr_io_trace_0_iaddr; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [31:0] csr_io_trace_0_insn; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_trace_0_exception; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  csr_io_trace_0_interrupt; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_privilegeMode; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mstatus; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_sstatus; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mepc; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_sepc; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mtval; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_stval; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mtvec; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_stvec; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mcause; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_scause; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_satp; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mip; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mie; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mscratch; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_sscratch; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_mideleg; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_difftest_medeleg; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_snapshot_minstret; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire [63:0] csr_io_snapshot_mcycle; // @[src/main/scala/rocket/RocketCore.scala 313:19]
  wire  bpu_clock; // @[src/main/scala/rocket/RocketCore.scala 351:19]
  wire  bpu_reset; // @[src/main/scala/rocket/RocketCore.scala 351:19]
  wire  alu_clock; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire  alu_reset; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire  alu_io_dw; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire [3:0] alu_io_fn; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire [63:0] alu_io_in2; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire [63:0] alu_io_in1; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire [63:0] alu_io_out; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire [63:0] alu_io_adder_out; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire  alu_io_cmp_out; // @[src/main/scala/rocket/RocketCore.scala 416:19]
  wire  div_clock; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_reset; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_req_ready; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_req_valid; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [3:0] div_io_req_bits_fn; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_req_bits_dw; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [63:0] div_io_req_bits_in1; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [63:0] div_io_req_bits_in2; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [4:0] div_io_req_bits_tag; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_kill; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_resp_ready; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  div_io_resp_valid; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [63:0] div_io_resp_bits_data; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire [4:0] div_io_resp_bits_tag; // @[src/main/scala/rocket/RocketCore.scala 454:19]
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_1_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_1_io_bits_address; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_1_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_2_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_2_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_2_io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_3_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_3_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_3_io_bits_minstret; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_3_io_bits_mcycle; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_delayer_clock; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_reset; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_skip; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_rfwen; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_i_fpwen; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [4:0] difftest_delayer_i_wpdest; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_i_wdest; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_i_pc; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_i_instr; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_i_special; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_skip; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_rfwen; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_o_fpwen; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [4:0] difftest_delayer_o_wpdest; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_o_wdest; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_o_pc; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [31:0] difftest_delayer_o_instr; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [7:0] difftest_delayer_o_special; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_module_4_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_4_io_bits_fpwen; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_4_io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_4_io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_4_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_4_io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_4_io_bits_special; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_delayer_1_clock; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_reset; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_i_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [4:0] difftest_delayer_1_i_address; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_i_data; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_i_nack; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_o_valid; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [4:0] difftest_delayer_1_o_address; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire [63:0] difftest_delayer_1_o_data; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_delayer_1_o_nack; // @[difftest/src/main/scala/util/Delayer.scala 54:15]
  wire  difftest_module_5_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_5_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_5_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_5_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_5_io_bits_address; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_5_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_5_io_bits_nack; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  PlusArgTimeout_clock; // @[src/main/scala/util/PlusArg.scala 89:11]
  wire  PlusArgTimeout_reset; // @[src/main/scala/util/PlusArg.scala 89:11]
  wire [31:0] PlusArgTimeout_io_count; // @[src/main/scala/util/PlusArg.scala 89:11]
  reg  id_reg_pause; // @[src/main/scala/rocket/RocketCore.scala 132:25]
  reg  imem_might_request_reg; // @[src/main/scala/rocket/RocketCore.scala 133:35]
  reg  ex_ctrl_fp; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_branch; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_jal; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_jalr; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_rxs2; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_zbk; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_zkn; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_zks; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [1:0] ex_ctrl_sel_alu2; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [1:0] ex_ctrl_sel_alu1; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [2:0] ex_ctrl_sel_imm; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_alu_dw; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [3:0] ex_ctrl_alu_fn; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [4:0] ex_ctrl_mem_cmd; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_mul; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg [2:0] ex_ctrl_csr; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  ex_ctrl_fence_i; // @[src/main/scala/rocket/RocketCore.scala 219:20]
  reg  mem_ctrl_fp; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_branch; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_jal; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_jalr; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_mul; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg [2:0] mem_ctrl_csr; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  mem_ctrl_fence_i; // @[src/main/scala/rocket/RocketCore.scala 220:21]
  reg  wb_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  wb_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  wb_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  wb_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  wb_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg [2:0] wb_ctrl_csr; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  wb_ctrl_fence_i; // @[src/main/scala/rocket/RocketCore.scala 221:20]
  reg  ex_reg_xcpt_interrupt; // @[src/main/scala/rocket/RocketCore.scala 223:35]
  reg  ex_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 224:35]
  reg  ex_reg_rvc; // @[src/main/scala/rocket/RocketCore.scala 225:35]
  reg  ex_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 227:35]
  reg  ex_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 228:35]
  reg  ex_reg_load_use; // @[src/main/scala/rocket/RocketCore.scala 229:35]
  reg [63:0] ex_reg_cause; // @[src/main/scala/rocket/RocketCore.scala 230:35]
  reg  ex_reg_replay; // @[src/main/scala/rocket/RocketCore.scala 231:26]
  reg [39:0] ex_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 232:22]
  reg [1:0] ex_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 233:28]
  reg [31:0] ex_reg_inst; // @[src/main/scala/rocket/RocketCore.scala 235:24]
  reg [31:0] ex_reg_raw_inst; // @[src/main/scala/rocket/RocketCore.scala 236:28]
  reg  mem_reg_xcpt_interrupt; // @[src/main/scala/rocket/RocketCore.scala 239:36]
  reg  mem_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 240:36]
  reg  mem_reg_rvc; // @[src/main/scala/rocket/RocketCore.scala 241:36]
  reg  mem_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 243:36]
  reg  mem_reg_replay; // @[src/main/scala/rocket/RocketCore.scala 244:36]
  reg  mem_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 245:36]
  reg [63:0] mem_reg_cause; // @[src/main/scala/rocket/RocketCore.scala 246:36]
  reg  mem_reg_slow_bypass; // @[src/main/scala/rocket/RocketCore.scala 247:36]
  reg  mem_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 250:27]
  reg [39:0] mem_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 251:23]
  reg [31:0] mem_reg_inst; // @[src/main/scala/rocket/RocketCore.scala 252:25]
  reg [1:0] mem_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 253:29]
  reg  mem_reg_hls_or_dv; // @[src/main/scala/rocket/RocketCore.scala 254:30]
  reg [31:0] mem_reg_raw_inst; // @[src/main/scala/rocket/RocketCore.scala 255:29]
  reg [63:0] mem_reg_wdata; // @[src/main/scala/rocket/RocketCore.scala 256:26]
  reg [63:0] mem_reg_rs2; // @[src/main/scala/rocket/RocketCore.scala 257:24]
  reg  mem_br_taken; // @[src/main/scala/rocket/RocketCore.scala 258:25]
  reg  wb_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 262:35]
  reg  wb_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 263:35]
  reg  wb_reg_replay; // @[src/main/scala/rocket/RocketCore.scala 264:35]
  reg  wb_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 265:35]
  reg [63:0] wb_reg_cause; // @[src/main/scala/rocket/RocketCore.scala 266:35]
  reg  wb_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 267:26]
  reg [39:0] wb_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 268:22]
  reg [1:0] wb_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 269:28]
  reg  wb_reg_hls_or_dv; // @[src/main/scala/rocket/RocketCore.scala 270:29]
  reg [31:0] wb_reg_inst; // @[src/main/scala/rocket/RocketCore.scala 273:24]
  reg [31:0] wb_reg_raw_inst; // @[src/main/scala/rocket/RocketCore.scala 274:28]
  reg [63:0] wb_reg_wdata; // @[src/main/scala/rocket/RocketCore.scala 275:25]
  wire  replay_wb_common = io_dmem_s2_nack | wb_reg_replay; // @[src/main/scala/rocket/RocketCore.scala 697:42]
  wire  replay_wb_rocc = wb_reg_valid & wb_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 698:37]
  wire  replay_wb = replay_wb_common | replay_wb_rocc; // @[src/main/scala/rocket/RocketCore.scala 700:36]
  wire  _T_92 = wb_reg_valid & wb_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 670:19]
  wire  _T_93 = wb_reg_valid & wb_ctrl_mem & io_dmem_s2_xcpt_ma_st; // @[src/main/scala/rocket/RocketCore.scala 670:34]
  wire  _T_95 = _T_92 & io_dmem_s2_xcpt_ma_ld; // @[src/main/scala/rocket/RocketCore.scala 671:34]
  wire  _T_97 = _T_92 & io_dmem_s2_xcpt_pf_st; // @[src/main/scala/rocket/RocketCore.scala 672:34]
  wire  _T_99 = _T_92 & io_dmem_s2_xcpt_pf_ld; // @[src/main/scala/rocket/RocketCore.scala 673:34]
  wire  _T_105 = _T_92 & io_dmem_s2_xcpt_ae_st; // @[src/main/scala/rocket/RocketCore.scala 676:34]
  wire  _T_107 = _T_92 & io_dmem_s2_xcpt_ae_ld; // @[src/main/scala/rocket/RocketCore.scala 677:34]
  wire  wb_xcpt = wb_reg_xcpt | _T_93 | _T_95 | _T_97 | _T_99 | _T_105 | _T_107; // @[src/main/scala/rocket/RocketCore.scala 1152:26]
  wire  take_pc_wb = replay_wb | wb_xcpt | csr_io_eret | wb_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 701:53]
  wire  _take_pc_mem_T = ~mem_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 570:35]
  wire  _mem_cfi_taken_T = mem_ctrl_branch & mem_br_taken; // @[src/main/scala/rocket/RocketCore.scala 567:40]
  wire  mem_cfi_taken = mem_ctrl_branch & mem_br_taken | mem_ctrl_jalr | mem_ctrl_jal; // @[src/main/scala/rocket/RocketCore.scala 567:74]
  wire  take_pc_mem = mem_reg_valid & ~mem_reg_xcpt & (mem_cfi_taken | mem_reg_sfence); // @[src/main/scala/rocket/RocketCore.scala 570:49]
  wire  take_pc_mem_wb = take_pc_wb | take_pc_mem; // @[src/main/scala/rocket/RocketCore.scala 280:35]
  wire [31:0] id_ctrl_decoder_decoded_plaInput = ibuf_io_inst_0_bits_inst_bits; // @[src/main/scala/chisel3/util/experimental/decode/decoder.scala 39:16 src/main/scala/chisel3/util/pla.scala 77:22]
  wire [31:0] id_ctrl_decoder_decoded_invInputs = ~id_ctrl_decoder_decoded_plaInput; // @[src/main/scala/chisel3/util/pla.scala 78:21]
  wire  id_ctrl_decoder_decoded_andMatrixInput_0 = id_ctrl_decoder_decoded_plaInput[0]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  id_ctrl_decoder_decoded_andMatrixInput_1 = id_ctrl_decoder_decoded_plaInput[1]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  id_ctrl_decoder_decoded_andMatrixInput_2 = id_ctrl_decoder_decoded_invInputs[2]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_3 = id_ctrl_decoder_decoded_invInputs[3]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_4 = id_ctrl_decoder_decoded_invInputs[5]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_5 = id_ctrl_decoder_decoded_invInputs[6]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_6 = id_ctrl_decoder_decoded_invInputs[12]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [6:0] _id_ctrl_decoder_decoded_T = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_1 = &_id_ctrl_decoder_decoded_T; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_4_1 = id_ctrl_decoder_decoded_invInputs[4]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [7:0] _id_ctrl_decoder_decoded_T_2 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_3 = &_id_ctrl_decoder_decoded_T_2; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_1 = id_ctrl_decoder_decoded_invInputs[13]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [7:0] _id_ctrl_decoder_decoded_T_4 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_5 = &_id_ctrl_decoder_decoded_T_4; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_3 = id_ctrl_decoder_decoded_invInputs[14]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [6:0] _id_ctrl_decoder_decoded_T_6 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_7 = &_id_ctrl_decoder_decoded_T_6; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_8 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_9 = &_id_ctrl_decoder_decoded_T_8; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_2_5 = id_ctrl_decoder_decoded_plaInput[2]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  id_ctrl_decoder_decoded_andMatrixInput_3_5 = id_ctrl_decoder_decoded_plaInput[3]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [8:0] _id_ctrl_decoder_decoded_T_10 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_11 = &_id_ctrl_decoder_decoded_T_10; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_3_6 = id_ctrl_decoder_decoded_plaInput[4]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [8:0] _id_ctrl_decoder_decoded_T_12 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_4,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_13 = &_id_ctrl_decoder_decoded_T_12; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] _id_ctrl_decoder_decoded_T_14 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_15 = &_id_ctrl_decoder_decoded_T_14; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] _id_ctrl_decoder_decoded_T_16 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_17 = &_id_ctrl_decoder_decoded_T_16; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_5_9 = id_ctrl_decoder_decoded_plaInput[5]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] _id_ctrl_decoder_decoded_T_18 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_19 = &_id_ctrl_decoder_decoded_T_18; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_20 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_21 = &_id_ctrl_decoder_decoded_T_20; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_9 = id_ctrl_decoder_decoded_invInputs[25]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_10 = id_ctrl_decoder_decoded_invInputs[26]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_11 = id_ctrl_decoder_decoded_invInputs[27]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_12 = id_ctrl_decoder_decoded_invInputs[28]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_13 = id_ctrl_decoder_decoded_invInputs[29]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_14 = id_ctrl_decoder_decoded_invInputs[31]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [6:0] id_ctrl_decoder_decoded_lo_11 = {id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_22 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_23 = &_id_ctrl_decoder_decoded_T_22; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_12 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_9,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_24 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_lo_12}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_25 = &_id_ctrl_decoder_decoded_T_24; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_11_2 = id_ctrl_decoder_decoded_invInputs[30]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [5:0] id_ctrl_decoder_decoded_lo_13 = {id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [12:0] _id_ctrl_decoder_decoded_T_26 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_13}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_27 = &_id_ctrl_decoder_decoded_T_26; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_14 = {id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_28 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_29 = &_id_ctrl_decoder_decoded_T_28; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_15 = {id_ctrl_decoder_decoded_andMatrixInput_9,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_30 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_31 = &_id_ctrl_decoder_decoded_T_30; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_15 = id_ctrl_decoder_decoded_plaInput[6]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] _id_ctrl_decoder_decoded_T_32 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_33 = &_id_ctrl_decoder_decoded_T_32; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_34 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_35 = &_id_ctrl_decoder_decoded_T_34; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_36 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_4_1,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_37 = &_id_ctrl_decoder_decoded_T_36; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_38 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_3,
    id_ctrl_decoder_decoded_andMatrixInput_4_1,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_39 = &_id_ctrl_decoder_decoded_T_38; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [9:0] _id_ctrl_decoder_decoded_T_40 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_41 = &_id_ctrl_decoder_decoded_T_40; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] _id_ctrl_decoder_decoded_T_42 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_43 = &_id_ctrl_decoder_decoded_T_42; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_4_22 = id_ctrl_decoder_decoded_invInputs[7]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_5_22 = id_ctrl_decoder_decoded_invInputs[8]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_6_21 = id_ctrl_decoder_decoded_invInputs[9]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_17 = id_ctrl_decoder_decoded_invInputs[10]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_8_11 = id_ctrl_decoder_decoded_invInputs[11]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_12_5 = id_ctrl_decoder_decoded_invInputs[15]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_13_4 = id_ctrl_decoder_decoded_invInputs[16]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_14_4 = id_ctrl_decoder_decoded_invInputs[17]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_15_1 = id_ctrl_decoder_decoded_invInputs[18]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_16 = id_ctrl_decoder_decoded_invInputs[19]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_17 = id_ctrl_decoder_decoded_invInputs[21]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_18 = id_ctrl_decoder_decoded_invInputs[22]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_19 = id_ctrl_decoder_decoded_invInputs[23]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_20 = id_ctrl_decoder_decoded_invInputs[24]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire [13:0] id_ctrl_decoder_decoded_lo_22 = {id_ctrl_decoder_decoded_andMatrixInput_14_4,
    id_ctrl_decoder_decoded_andMatrixInput_15_1,id_ctrl_decoder_decoded_andMatrixInput_16,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_21 = {id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_8_11,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_12_5,id_ctrl_decoder_decoded_andMatrixInput_13_4}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [27:0] _id_ctrl_decoder_decoded_T_44 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_4_22,
    id_ctrl_decoder_decoded_andMatrixInput_5_22,id_ctrl_decoder_decoded_andMatrixInput_6_21,
    id_ctrl_decoder_decoded_hi_lo_21,id_ctrl_decoder_decoded_lo_22}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_45 = &_id_ctrl_decoder_decoded_T_44; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] id_ctrl_decoder_decoded_lo_23 = {id_ctrl_decoder_decoded_andMatrixInput_13_4,
    id_ctrl_decoder_decoded_andMatrixInput_14_4,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [7:0] id_ctrl_decoder_decoded_hi_lo_22 = {id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_andMatrixInput_6_21,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_andMatrixInput_8_11,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_12_5}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [30:0] _id_ctrl_decoder_decoded_T_46 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_hi_lo_22,id_ctrl_decoder_decoded_lo_23}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_47 = &_id_ctrl_decoder_decoded_T_46; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_19 = id_ctrl_decoder_decoded_plaInput[12]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [9:0] _id_ctrl_decoder_decoded_T_48 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_49 = &_id_ctrl_decoder_decoded_T_48; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_25 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] _id_ctrl_decoder_decoded_T_50 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_25}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_51 = &_id_ctrl_decoder_decoded_T_50; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_52 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_25}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_53 = &_id_ctrl_decoder_decoded_T_52; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_54 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_55 = &_id_ctrl_decoder_decoded_T_54; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_28 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_56 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_28}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_57 = &_id_ctrl_decoder_decoded_T_56; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_58 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_59 = &_id_ctrl_decoder_decoded_T_58; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_60 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_7_1}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_61 = &_id_ctrl_decoder_decoded_T_60; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_62 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_63 = &_id_ctrl_decoder_decoded_T_62; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_64 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_19}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_65 = &_id_ctrl_decoder_decoded_T_64; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_28 = id_ctrl_decoder_decoded_plaInput[13]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] _id_ctrl_decoder_decoded_T_66 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_67 = &_id_ctrl_decoder_decoded_T_66; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_68 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_69 = &_id_ctrl_decoder_decoded_T_68; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [4:0] id_ctrl_decoder_decoded_lo_35 = {id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [10:0] _id_ctrl_decoder_decoded_T_70 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_lo_35}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_71 = &_id_ctrl_decoder_decoded_T_70; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_72 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_73 = &_id_ctrl_decoder_decoded_T_72; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_37 = {id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_74 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_lo_37}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_75 = &_id_ctrl_decoder_decoded_T_74; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_76 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_28}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_77 = &_id_ctrl_decoder_decoded_T_76; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_78 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_79 = &_id_ctrl_decoder_decoded_T_78; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_80 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_7_28}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_81 = &_id_ctrl_decoder_decoded_T_80; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_41 = {id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_82 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_41}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_83 = &_id_ctrl_decoder_decoded_T_82; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_8_27 = id_ctrl_decoder_decoded_plaInput[14]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [8:0] _id_ctrl_decoder_decoded_T_84 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_85 = &_id_ctrl_decoder_decoded_T_84; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_43 = {id_ctrl_decoder_decoded_andMatrixInput_8_27,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] _id_ctrl_decoder_decoded_T_86 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_43}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_87 = &_id_ctrl_decoder_decoded_T_86; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_88 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_89 = &_id_ctrl_decoder_decoded_T_88; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_45 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_90 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_45}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_91 = &_id_ctrl_decoder_decoded_T_90; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_92 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_43}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_93 = &_id_ctrl_decoder_decoded_T_92; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_47 = {id_ctrl_decoder_decoded_andMatrixInput_8_27,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [14:0] _id_ctrl_decoder_decoded_T_94 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_47}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_95 = &_id_ctrl_decoder_decoded_T_94; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_48 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_andMatrixInput_9,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_96 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_48}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_97 = &_id_ctrl_decoder_decoded_T_96; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_49 = {id_ctrl_decoder_decoded_andMatrixInput_8_27,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_98 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_49}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_99 = &_id_ctrl_decoder_decoded_T_98; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_100 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_47}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_101 = &_id_ctrl_decoder_decoded_T_100; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [15:0] _id_ctrl_decoder_decoded_T_102 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_48}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_103 = &_id_ctrl_decoder_decoded_T_102; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_104 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_43}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_105 = &_id_ctrl_decoder_decoded_T_104; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_106 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_107 = &_id_ctrl_decoder_decoded_T_106; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_108 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_109 = &_id_ctrl_decoder_decoded_T_108; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_110 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_111 = &_id_ctrl_decoder_decoded_T_110; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_112 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_113 = &_id_ctrl_decoder_decoded_T_112; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_114 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_lo_43}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_115 = &_id_ctrl_decoder_decoded_T_114; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] _id_ctrl_decoder_decoded_T_116 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_117 = &_id_ctrl_decoder_decoded_T_116; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_118 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_119 = &_id_ctrl_decoder_decoded_T_118; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] _id_ctrl_decoder_decoded_T_120 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_121 = &_id_ctrl_decoder_decoded_T_120; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [9:0] _id_ctrl_decoder_decoded_T_122 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_8_27}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_123 = &_id_ctrl_decoder_decoded_T_122; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_57 = id_ctrl_decoder_decoded_plaInput[25]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [6:0] id_ctrl_decoder_decoded_lo_62 = {id_ctrl_decoder_decoded_andMatrixInput_7_57,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_12,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] _id_ctrl_decoder_decoded_T_124 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_125 = &_id_ctrl_decoder_decoded_T_124; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_126 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_127 = &_id_ctrl_decoder_decoded_T_126; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_128 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_129 = &_id_ctrl_decoder_decoded_T_128; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_130 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_131 = &_id_ctrl_decoder_decoded_T_130; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [13:0] _id_ctrl_decoder_decoded_T_132 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_133 = &_id_ctrl_decoder_decoded_T_132; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_134 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_135 = &_id_ctrl_decoder_decoded_T_134; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] _id_ctrl_decoder_decoded_T_136 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_lo_62}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_137 = &_id_ctrl_decoder_decoded_T_136; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_9_35 = id_ctrl_decoder_decoded_plaInput[27]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] id_ctrl_decoder_decoded_lo_69 = {id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_9_35,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [12:0] _id_ctrl_decoder_decoded_T_138 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_69}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_139 = &_id_ctrl_decoder_decoded_T_138; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_7_65 = id_ctrl_decoder_decoded_invInputs[20]; // @[src/main/scala/chisel3/util/pla.scala 91:29]
  wire  id_ctrl_decoder_decoded_andMatrixInput_13_30 = id_ctrl_decoder_decoded_plaInput[28]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] id_ctrl_decoder_decoded_lo_70 = {id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [16:0] _id_ctrl_decoder_decoded_T_140 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_65,id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_lo_70}
    ; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_141 = &_id_ctrl_decoder_decoded_T_140; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [9:0] id_ctrl_decoder_decoded_hi_71 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_7_65}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [18:0] _id_ctrl_decoder_decoded_T_142 = {id_ctrl_decoder_decoded_hi_71,id_ctrl_decoder_decoded_andMatrixInput_17,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,
    id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_143 = &_id_ctrl_decoder_decoded_T_142; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_18_3 = id_ctrl_decoder_decoded_plaInput[21]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_67 = {id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] id_ctrl_decoder_decoded_lo_72 = {id_ctrl_decoder_decoded_andMatrixInput_14_4,
    id_ctrl_decoder_decoded_andMatrixInput_15_1,id_ctrl_decoder_decoded_andMatrixInput_16,
    id_ctrl_decoder_decoded_andMatrixInput_7_65,id_ctrl_decoder_decoded_andMatrixInput_18_3,
    id_ctrl_decoder_decoded_andMatrixInput_18,id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_67
    }; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [27:0] _id_ctrl_decoder_decoded_T_144 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_6_15,id_ctrl_decoder_decoded_andMatrixInput_4_22,
    id_ctrl_decoder_decoded_andMatrixInput_5_22,id_ctrl_decoder_decoded_andMatrixInput_6_21,
    id_ctrl_decoder_decoded_hi_lo_21,id_ctrl_decoder_decoded_lo_72}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_145 = &_id_ctrl_decoder_decoded_T_144; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [14:0] id_ctrl_decoder_decoded_lo_73 = {id_ctrl_decoder_decoded_andMatrixInput_13_4,
    id_ctrl_decoder_decoded_andMatrixInput_14_4,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_65,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_67}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [30:0] _id_ctrl_decoder_decoded_T_146 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_hi_lo_22,id_ctrl_decoder_decoded_lo_73}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_147 = &_id_ctrl_decoder_decoded_T_146; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_16_6 = id_ctrl_decoder_decoded_plaInput[20]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire  id_ctrl_decoder_decoded_andMatrixInput_18_5 = id_ctrl_decoder_decoded_plaInput[22]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_69 = {id_ctrl_decoder_decoded_andMatrixInput_9,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] id_ctrl_decoder_decoded_lo_74 = {id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_16_6,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18_5,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20,id_ctrl_decoder_decoded_lo_lo_69
    }; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_73 = {id_ctrl_decoder_decoded_andMatrixInput_8_11,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_12_5,
    id_ctrl_decoder_decoded_andMatrixInput_13_4,id_ctrl_decoder_decoded_andMatrixInput_14_4}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [27:0] _id_ctrl_decoder_decoded_T_148 = {id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_andMatrixInput_6_21,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_hi_lo_73,id_ctrl_decoder_decoded_lo_74}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_149 = &_id_ctrl_decoder_decoded_T_148; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_70 = {id_ctrl_decoder_decoded_andMatrixInput_20,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] id_ctrl_decoder_decoded_lo_75 = {id_ctrl_decoder_decoded_andMatrixInput_13_4,
    id_ctrl_decoder_decoded_andMatrixInput_14_4,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_16_6,
    id_ctrl_decoder_decoded_andMatrixInput_17,id_ctrl_decoder_decoded_andMatrixInput_18_5,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_70}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [31:0] _id_ctrl_decoder_decoded_T_150 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_hi_lo_22,id_ctrl_decoder_decoded_lo_75}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_151 = &_id_ctrl_decoder_decoded_T_150; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_76 = {id_ctrl_decoder_decoded_andMatrixInput_6_21,
    id_ctrl_decoder_decoded_andMatrixInput_7_57,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [16:0] _id_ctrl_decoder_decoded_T_152 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_lo_76}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_153 = &_id_ctrl_decoder_decoded_T_152; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [8:0] id_ctrl_decoder_decoded_lo_77 = {id_ctrl_decoder_decoded_andMatrixInput_6_21,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_7_57,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [17:0] _id_ctrl_decoder_decoded_T_154 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_lo_77}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_155 = &_id_ctrl_decoder_decoded_T_154; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [4:0] id_ctrl_decoder_decoded_lo_lo_73 = {id_ctrl_decoder_decoded_andMatrixInput_11,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [9:0] id_ctrl_decoder_decoded_lo_78 = {id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_7_57,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_11_2,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [9:0] id_ctrl_decoder_decoded_hi_78 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_andMatrixInput_6_21}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [19:0] _id_ctrl_decoder_decoded_T_156 = {id_ctrl_decoder_decoded_hi_78,id_ctrl_decoder_decoded_lo_78}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_157 = &_id_ctrl_decoder_decoded_T_156; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [10:0] id_ctrl_decoder_decoded_lo_79 = {id_ctrl_decoder_decoded_andMatrixInput_8_11,
    id_ctrl_decoder_decoded_andMatrixInput_6,id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_7_57,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_lo_lo_73}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [4:0] id_ctrl_decoder_decoded_hi_lo_78 = {id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_andMatrixInput_6_21,id_ctrl_decoder_decoded_andMatrixInput_7_17}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [21:0] _id_ctrl_decoder_decoded_T_158 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_hi_lo_78,id_ctrl_decoder_decoded_lo_79}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_159 = &_id_ctrl_decoder_decoded_T_158; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [6:0] id_ctrl_decoder_decoded_lo_80 = {id_ctrl_decoder_decoded_andMatrixInput_7_28,
    id_ctrl_decoder_decoded_andMatrixInput_6_3,id_ctrl_decoder_decoded_andMatrixInput_9_35,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_13,
    id_ctrl_decoder_decoded_andMatrixInput_11_2,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] _id_ctrl_decoder_decoded_T_160 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_lo_80}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_161 = &_id_ctrl_decoder_decoded_T_160; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_11_43 = id_ctrl_decoder_decoded_plaInput[29]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] id_ctrl_decoder_decoded_lo_81 = {id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_11_43}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _id_ctrl_decoder_decoded_T_162 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_lo_81}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_163 = &_id_ctrl_decoder_decoded_T_162; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_14_36 = id_ctrl_decoder_decoded_plaInput[30]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [7:0] id_ctrl_decoder_decoded_lo_82 = {id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14_36,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_164 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_6,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_82}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_165 = &_id_ctrl_decoder_decoded_T_164; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [5:0] id_ctrl_decoder_decoded_lo_83 = {id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_14_36}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _id_ctrl_decoder_decoded_T_166 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_lo_83}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_167 = &_id_ctrl_decoder_decoded_T_166; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_84 = {id_ctrl_decoder_decoded_andMatrixInput_7_1,
    id_ctrl_decoder_decoded_andMatrixInput_8_27,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14_36,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_168 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_4,id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_19,id_ctrl_decoder_decoded_lo_84}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_169 = &_id_ctrl_decoder_decoded_T_168; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_85 = {id_ctrl_decoder_decoded_andMatrixInput_8_27,
    id_ctrl_decoder_decoded_andMatrixInput_9,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_13,id_ctrl_decoder_decoded_andMatrixInput_14_36,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] _id_ctrl_decoder_decoded_T_170 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_85}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_171 = &_id_ctrl_decoder_decoded_T_170; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [15:0] _id_ctrl_decoder_decoded_T_172 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3_6,id_ctrl_decoder_decoded_andMatrixInput_5_9,
    id_ctrl_decoder_decoded_andMatrixInput_5,id_ctrl_decoder_decoded_andMatrixInput_7_19,
    id_ctrl_decoder_decoded_andMatrixInput_7_1,id_ctrl_decoder_decoded_lo_85}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_173 = &_id_ctrl_decoder_decoded_T_172; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_20_7 = id_ctrl_decoder_decoded_plaInput[24]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_82 = {id_ctrl_decoder_decoded_andMatrixInput_7_57,
    id_ctrl_decoder_decoded_andMatrixInput_10,id_ctrl_decoder_decoded_andMatrixInput_9_35,
    id_ctrl_decoder_decoded_andMatrixInput_13_30,id_ctrl_decoder_decoded_andMatrixInput_11_43,
    id_ctrl_decoder_decoded_andMatrixInput_14_36,id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [13:0] id_ctrl_decoder_decoded_lo_87 = {id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_65,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_andMatrixInput_20_7,
    id_ctrl_decoder_decoded_lo_lo_82}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [27:0] _id_ctrl_decoder_decoded_T_174 = {id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_andMatrixInput_5_22,
    id_ctrl_decoder_decoded_andMatrixInput_6_21,id_ctrl_decoder_decoded_andMatrixInput_7_17,
    id_ctrl_decoder_decoded_hi_lo_73,id_ctrl_decoder_decoded_lo_87}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_175 = &_id_ctrl_decoder_decoded_T_174; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_83 = {id_ctrl_decoder_decoded_andMatrixInput_20_7,
    id_ctrl_decoder_decoded_andMatrixInput_7_57,id_ctrl_decoder_decoded_andMatrixInput_10,
    id_ctrl_decoder_decoded_andMatrixInput_9_35,id_ctrl_decoder_decoded_andMatrixInput_13_30,
    id_ctrl_decoder_decoded_andMatrixInput_11_43,id_ctrl_decoder_decoded_andMatrixInput_14_36,
    id_ctrl_decoder_decoded_andMatrixInput_14}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [15:0] id_ctrl_decoder_decoded_lo_88 = {id_ctrl_decoder_decoded_andMatrixInput_13_4,
    id_ctrl_decoder_decoded_andMatrixInput_14_4,id_ctrl_decoder_decoded_andMatrixInput_15_1,
    id_ctrl_decoder_decoded_andMatrixInput_16,id_ctrl_decoder_decoded_andMatrixInput_7_65,
    id_ctrl_decoder_decoded_andMatrixInput_18_3,id_ctrl_decoder_decoded_andMatrixInput_18,
    id_ctrl_decoder_decoded_andMatrixInput_19,id_ctrl_decoder_decoded_lo_lo_83}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [31:0] _id_ctrl_decoder_decoded_T_176 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2,
    id_ctrl_decoder_decoded_andMatrixInput_3,id_ctrl_decoder_decoded_andMatrixInput_3_6,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_andMatrixInput_6_15,
    id_ctrl_decoder_decoded_andMatrixInput_4_22,id_ctrl_decoder_decoded_hi_lo_22,id_ctrl_decoder_decoded_lo_88}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_177 = &_id_ctrl_decoder_decoded_T_176; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire  id_ctrl_decoder_decoded_andMatrixInput_11_51 = id_ctrl_decoder_decoded_plaInput[31]; // @[src/main/scala/chisel3/util/pla.scala 90:45]
  wire [5:0] id_ctrl_decoder_decoded_lo_89 = {id_ctrl_decoder_decoded_andMatrixInput_5,
    id_ctrl_decoder_decoded_andMatrixInput_7_28,id_ctrl_decoder_decoded_andMatrixInput_6_3,
    id_ctrl_decoder_decoded_andMatrixInput_11,id_ctrl_decoder_decoded_andMatrixInput_12,
    id_ctrl_decoder_decoded_andMatrixInput_11_51}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire [11:0] _id_ctrl_decoder_decoded_T_178 = {id_ctrl_decoder_decoded_andMatrixInput_0,
    id_ctrl_decoder_decoded_andMatrixInput_1,id_ctrl_decoder_decoded_andMatrixInput_2_5,
    id_ctrl_decoder_decoded_andMatrixInput_3_5,id_ctrl_decoder_decoded_andMatrixInput_4_1,
    id_ctrl_decoder_decoded_andMatrixInput_5_9,id_ctrl_decoder_decoded_lo_89}; // @[src/main/scala/chisel3/util/pla.scala 98:53]
  wire  _id_ctrl_decoder_decoded_T_179 = &_id_ctrl_decoder_decoded_T_178; // @[src/main/scala/chisel3/util/pla.scala 98:70]
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T = {_id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_141}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_1 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_2 = |_id_ctrl_decoder_decoded_T_11; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_3 = |_id_ctrl_decoder_decoded_T_49; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_4 = |_id_ctrl_decoder_decoded_T_65; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_5 = |_id_ctrl_decoder_decoded_T_77; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_6 = {_id_ctrl_decoder_decoded_T_45,_id_ctrl_decoder_decoded_T_65
    ,_id_ctrl_decoder_decoded_T_77,_id_ctrl_decoder_decoded_T_145,_id_ctrl_decoder_decoded_T_149,
    _id_ctrl_decoder_decoded_T_153,_id_ctrl_decoder_decoded_T_175}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_7 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_6; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo = {_id_ctrl_decoder_decoded_T_95,
    _id_ctrl_decoder_decoded_T_101,_id_ctrl_decoder_decoded_T_133,_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_141}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [10:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 = {_id_ctrl_decoder_decoded_T_55,
    _id_ctrl_decoder_decoded_T_65,_id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_71,
    _id_ctrl_decoder_decoded_T_77,_id_ctrl_decoder_decoded_T_91,id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1 = {_id_ctrl_decoder_decoded_T_27,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_41,_id_ctrl_decoder_decoded_T_43,
    _id_ctrl_decoder_decoded_T_51}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [21:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_8 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5,
    _id_ctrl_decoder_decoded_T_9,_id_ctrl_decoder_decoded_T_13,_id_ctrl_decoder_decoded_T_15,
    _id_ctrl_decoder_decoded_T_23,id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_1}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_9 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_8; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_10 = {_id_ctrl_decoder_decoded_T_125,
    _id_ctrl_decoder_decoded_T_127,_id_ctrl_decoder_decoded_T_133}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_11 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_10; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_12 = {_id_ctrl_decoder_decoded_T_19,
    _id_ctrl_decoder_decoded_T_161,_id_ctrl_decoder_decoded_T_163}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_13 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_12; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_14 = {_id_ctrl_decoder_decoded_T_141,
    _id_ctrl_decoder_decoded_T_161,_id_ctrl_decoder_decoded_T_167}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_15 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_14; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [3:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_16 = {_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_141,_id_ctrl_decoder_decoded_T_153,_id_ctrl_decoder_decoded_T_179}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_17 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_16; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_18 = |_id_ctrl_decoder_decoded_T_71; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_19 = |_id_ctrl_decoder_decoded_T_153; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_20 = {_id_ctrl_decoder_decoded_T_3,_id_ctrl_decoder_decoded_T_5,
    _id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_143,_id_ctrl_decoder_decoded_T_159}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_21 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_20; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_4 = {_id_ctrl_decoder_decoded_T_105,
    _id_ctrl_decoder_decoded_T_109,_id_ctrl_decoder_decoded_T_123,_id_ctrl_decoder_decoded_T_129,
    _id_ctrl_decoder_decoded_T_135}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [10:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_22 = {_id_ctrl_decoder_decoded_T_51,
    _id_ctrl_decoder_decoded_T_55,_id_ctrl_decoder_decoded_T_61,_id_ctrl_decoder_decoded_T_91,
    _id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_101,id_ctrl_decoder_decoded_orMatrixOutputs_lo_4}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_23 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_22; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [5:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_5 = {_id_ctrl_decoder_decoded_T_131,
    _id_ctrl_decoder_decoded_T_137,_id_ctrl_decoder_decoded_T_165,_id_ctrl_decoder_decoded_T_169,
    _id_ctrl_decoder_decoded_T_171,_id_ctrl_decoder_decoded_T_173}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [11:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_24 = {_id_ctrl_decoder_decoded_T_35,
    _id_ctrl_decoder_decoded_T_81,_id_ctrl_decoder_decoded_T_83,_id_ctrl_decoder_decoded_T_113,
    _id_ctrl_decoder_decoded_T_115,_id_ctrl_decoder_decoded_T_119,id_ctrl_decoder_decoded_orMatrixOutputs_lo_5}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_25 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_24; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [7:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_26 = {_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_73,_id_ctrl_decoder_decoded_T_85,_id_ctrl_decoder_decoded_T_87,
    _id_ctrl_decoder_decoded_T_89,_id_ctrl_decoder_decoded_T_93,_id_ctrl_decoder_decoded_T_99,
    _id_ctrl_decoder_decoded_T_133}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_27 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_26; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_28 = {_id_ctrl_decoder_decoded_T_69,
    _id_ctrl_decoder_decoded_T_75,_id_ctrl_decoder_decoded_T_89,_id_ctrl_decoder_decoded_T_165,
    _id_ctrl_decoder_decoded_T_169,_id_ctrl_decoder_decoded_T_171,_id_ctrl_decoder_decoded_T_173}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_29 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_28; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_12 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5,
    _id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_15,_id_ctrl_decoder_decoded_T_25,
    _id_ctrl_decoder_decoded_T_27,_id_ctrl_decoder_decoded_T_39,_id_ctrl_decoder_decoded_T_43,
    _id_ctrl_decoder_decoded_T_51,_id_ctrl_decoder_decoded_T_59}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [18:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_30 = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_12,
    _id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_77,
    _id_ctrl_decoder_decoded_T_89,_id_ctrl_decoder_decoded_T_91,_id_ctrl_decoder_decoded_T_103,
    _id_ctrl_decoder_decoded_T_139,_id_ctrl_decoder_decoded_T_141,_id_ctrl_decoder_decoded_T_153}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_31 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_30; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [3:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_32 = {_id_ctrl_decoder_decoded_T_33,
    _id_ctrl_decoder_decoded_T_43,_id_ctrl_decoder_decoded_T_107,_id_ctrl_decoder_decoded_T_117}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_33 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_32; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_34 = {_id_ctrl_decoder_decoded_T_15,
    _id_ctrl_decoder_decoded_T_43}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_35 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_34; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [5:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_10 = {_id_ctrl_decoder_decoded_T_57,
    _id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_91,_id_ctrl_decoder_decoded_T_97,
    _id_ctrl_decoder_decoded_T_111,_id_ctrl_decoder_decoded_T_121}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [11:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_36 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5
    ,_id_ctrl_decoder_decoded_T_9,_id_ctrl_decoder_decoded_T_13,_id_ctrl_decoder_decoded_T_41,
    _id_ctrl_decoder_decoded_T_53,id_ctrl_decoder_decoded_orMatrixOutputs_lo_10}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_37 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_36; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6 = {_id_ctrl_decoder_decoded_T_101,
    _id_ctrl_decoder_decoded_T_133,_id_ctrl_decoder_decoded_T_139,_id_ctrl_decoder_decoded_T_141,
    _id_ctrl_decoder_decoded_T_155}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [10:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_11 = {_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_79,_id_ctrl_decoder_decoded_T_89,
    _id_ctrl_decoder_decoded_T_91,_id_ctrl_decoder_decoded_T_95,id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9 = {_id_ctrl_decoder_decoded_T_29,
    _id_ctrl_decoder_decoded_T_39,_id_ctrl_decoder_decoded_T_51,_id_ctrl_decoder_decoded_T_55,
    _id_ctrl_decoder_decoded_T_63}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [21:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_38 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_13,_id_ctrl_decoder_decoded_T_23,
    _id_ctrl_decoder_decoded_T_27,id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_39 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_38; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_40 = {_id_ctrl_decoder_decoded_T_17,
    _id_ctrl_decoder_decoded_T_43}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_41 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_40; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 = {_id_ctrl_decoder_decoded_T_53,
    _id_ctrl_decoder_decoded_T_57,_id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_91,
    _id_ctrl_decoder_decoded_T_97,_id_ctrl_decoder_decoded_T_111,_id_ctrl_decoder_decoded_T_121}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [13:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_42 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_13,_id_ctrl_decoder_decoded_T_15,
    _id_ctrl_decoder_decoded_T_41,_id_ctrl_decoder_decoded_T_43,id_ctrl_decoder_decoded_orMatrixOutputs_lo_12}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_43 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_42; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5,
    _id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_13,_id_ctrl_decoder_decoded_T_15,
    _id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_27,_id_ctrl_decoder_decoded_T_29,
    _id_ctrl_decoder_decoded_T_33,_id_ctrl_decoder_decoded_T_39}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [18:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_44 = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_17,
    _id_ctrl_decoder_decoded_T_51,_id_ctrl_decoder_decoded_T_55,_id_ctrl_decoder_decoded_T_67,
    _id_ctrl_decoder_decoded_T_91,_id_ctrl_decoder_decoded_T_95,_id_ctrl_decoder_decoded_T_101,
    _id_ctrl_decoder_decoded_T_107,_id_ctrl_decoder_decoded_T_117,_id_ctrl_decoder_decoded_T_133}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_45 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_44; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [5:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_15 = {_id_ctrl_decoder_decoded_T_89,
    _id_ctrl_decoder_decoded_T_101,_id_ctrl_decoder_decoded_T_133,_id_ctrl_decoder_decoded_T_139,
    _id_ctrl_decoder_decoded_T_141,_id_ctrl_decoder_decoded_T_157}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [12:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_48 = {_id_ctrl_decoder_decoded_T_19,
    _id_ctrl_decoder_decoded_T_21,_id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_27,
    _id_ctrl_decoder_decoded_T_29,_id_ctrl_decoder_decoded_T_31,_id_ctrl_decoder_decoded_T_71,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_15}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_49 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_48; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_50 = |_id_ctrl_decoder_decoded_T_41; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_51 = |_id_ctrl_decoder_decoded_T_43; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [1:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_52 = {_id_ctrl_decoder_decoded_T_33,
    _id_ctrl_decoder_decoded_T_89}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_53 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_52; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [6:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_11 = {_id_ctrl_decoder_decoded_T_133,
    _id_ctrl_decoder_decoded_T_139,_id_ctrl_decoder_decoded_T_143,_id_ctrl_decoder_decoded_T_147,
    _id_ctrl_decoder_decoded_T_151,_id_ctrl_decoder_decoded_T_159,_id_ctrl_decoder_decoded_T_177}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [14:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 = {_id_ctrl_decoder_decoded_T_59,
    _id_ctrl_decoder_decoded_T_67,_id_ctrl_decoder_decoded_T_71,_id_ctrl_decoder_decoded_T_77,
    _id_ctrl_decoder_decoded_T_89,_id_ctrl_decoder_decoded_T_91,_id_ctrl_decoder_decoded_T_95,
    _id_ctrl_decoder_decoded_T_101,id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_11}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [6:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_14 = {_id_ctrl_decoder_decoded_T_29,
    _id_ctrl_decoder_decoded_T_37,_id_ctrl_decoder_decoded_T_39,_id_ctrl_decoder_decoded_T_43,
    _id_ctrl_decoder_decoded_T_47,_id_ctrl_decoder_decoded_T_51,_id_ctrl_decoder_decoded_T_55}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire [29:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_54 = {_id_ctrl_decoder_decoded_T_1,_id_ctrl_decoder_decoded_T_5
    ,_id_ctrl_decoder_decoded_T_7,_id_ctrl_decoder_decoded_T_11,_id_ctrl_decoder_decoded_T_13,
    _id_ctrl_decoder_decoded_T_15,_id_ctrl_decoder_decoded_T_23,_id_ctrl_decoder_decoded_T_27,
    id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_14,id_ctrl_decoder_decoded_orMatrixOutputs_lo_16}; // @[src/main/scala/chisel3/util/pla.scala 114:19]
  wire  _id_ctrl_decoder_decoded_orMatrixOutputs_T_55 = |_id_ctrl_decoder_decoded_orMatrixOutputs_T_54; // @[src/main/scala/chisel3/util/pla.scala 114:36]
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_12 = {1'h0,_id_ctrl_decoder_decoded_orMatrixOutputs_T_11,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_9,_id_ctrl_decoder_decoded_orMatrixOutputs_T_7,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_5,_id_ctrl_decoder_decoded_orMatrixOutputs_T_4,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_3,_id_ctrl_decoder_decoded_orMatrixOutputs_T_2,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_1,1'h0}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [10:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_15 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_23,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_21,_id_ctrl_decoder_decoded_orMatrixOutputs_T_19,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_18,_id_ctrl_decoder_decoded_orMatrixOutputs_T_17,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_15,_id_ctrl_decoder_decoded_orMatrixOutputs_T_13,1'h0,1'h0,2'h0}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_6 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_33,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_31,_id_ctrl_decoder_decoded_orMatrixOutputs_T_29,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_27,_id_ctrl_decoder_decoded_orMatrixOutputs_T_25}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [10:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15 = {_id_ctrl_decoder_decoded_orMatrixOutputs_T_55,1'h0,1'h0
    ,_id_ctrl_decoder_decoded_orMatrixOutputs_T_53,_id_ctrl_decoder_decoded_orMatrixOutputs_T_51,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_50,_id_ctrl_decoder_decoded_orMatrixOutputs_T_49,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_39,1'h0,2'h0}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [42:0] id_ctrl_decoder_decoded_orMatrixOutputs = {id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_45,_id_ctrl_decoder_decoded_orMatrixOutputs_T_43,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_41,_id_ctrl_decoder_decoded_orMatrixOutputs_T_39,
    _id_ctrl_decoder_decoded_orMatrixOutputs_T_37,_id_ctrl_decoder_decoded_orMatrixOutputs_T_35,
    id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_6,id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_15,
    id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_12}; // @[src/main/scala/chisel3/util/pla.scala 102:36]
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[9],
    id_ctrl_decoder_decoded_orMatrixOutputs[8],id_ctrl_decoder_decoded_orMatrixOutputs[7],
    id_ctrl_decoder_decoded_orMatrixOutputs[6],id_ctrl_decoder_decoded_orMatrixOutputs[5],
    id_ctrl_decoder_decoded_orMatrixOutputs[4],id_ctrl_decoder_decoded_orMatrixOutputs[3],
    id_ctrl_decoder_decoded_orMatrixOutputs[2],id_ctrl_decoder_decoded_orMatrixOutputs[1],
    id_ctrl_decoder_decoded_orMatrixOutputs[0]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[14],
    id_ctrl_decoder_decoded_orMatrixOutputs[13],id_ctrl_decoder_decoded_orMatrixOutputs[12],
    id_ctrl_decoder_decoded_orMatrixOutputs[11],id_ctrl_decoder_decoded_orMatrixOutputs[10]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [20:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[20],
    id_ctrl_decoder_decoded_orMatrixOutputs[19],id_ctrl_decoder_decoded_orMatrixOutputs[18],
    id_ctrl_decoder_decoded_orMatrixOutputs[17],id_ctrl_decoder_decoded_orMatrixOutputs[16],
    id_ctrl_decoder_decoded_orMatrixOutputs[15],id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo,
    id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[25],
    id_ctrl_decoder_decoded_orMatrixOutputs[24],id_ctrl_decoder_decoded_orMatrixOutputs[23],
    id_ctrl_decoder_decoded_orMatrixOutputs[22],id_ctrl_decoder_decoded_orMatrixOutputs[21]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [10:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[31],
    id_ctrl_decoder_decoded_orMatrixOutputs[30],id_ctrl_decoder_decoded_orMatrixOutputs[29],
    id_ctrl_decoder_decoded_orMatrixOutputs[28],id_ctrl_decoder_decoded_orMatrixOutputs[27],
    id_ctrl_decoder_decoded_orMatrixOutputs[26],id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo = {id_ctrl_decoder_decoded_orMatrixOutputs[36],
    id_ctrl_decoder_decoded_orMatrixOutputs[35],id_ctrl_decoder_decoded_orMatrixOutputs[34],
    id_ctrl_decoder_decoded_orMatrixOutputs[33],id_ctrl_decoder_decoded_orMatrixOutputs[32]}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire [42:0] id_ctrl_decoder_decoded_invMatrixOutputs = {id_ctrl_decoder_decoded_orMatrixOutputs[42],
    id_ctrl_decoder_decoded_orMatrixOutputs[41],id_ctrl_decoder_decoded_orMatrixOutputs[40],
    id_ctrl_decoder_decoded_orMatrixOutputs[39],id_ctrl_decoder_decoded_orMatrixOutputs[38],
    id_ctrl_decoder_decoded_orMatrixOutputs[37],id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo,
    id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo,id_ctrl_decoder_decoded_invMatrixOutputs_lo}; // @[src/main/scala/chisel3/util/pla.scala 120:37]
  wire  id_ctrl_decoder_0 = id_ctrl_decoder_decoded_invMatrixOutputs[42]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_1 = id_ctrl_decoder_decoded_invMatrixOutputs[41]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_2 = id_ctrl_decoder_decoded_invMatrixOutputs[40]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_3 = id_ctrl_decoder_decoded_invMatrixOutputs[39]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_4 = id_ctrl_decoder_decoded_invMatrixOutputs[38]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_5 = id_ctrl_decoder_decoded_invMatrixOutputs[37]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_6 = id_ctrl_decoder_decoded_invMatrixOutputs[36]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_7 = id_ctrl_decoder_decoded_invMatrixOutputs[35]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_8 = id_ctrl_decoder_decoded_invMatrixOutputs[34]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_9 = id_ctrl_decoder_decoded_invMatrixOutputs[33]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_10 = id_ctrl_decoder_decoded_invMatrixOutputs[32]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [1:0] id_ctrl_decoder_11 = id_ctrl_decoder_decoded_invMatrixOutputs[31:30]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [1:0] id_ctrl_decoder_12 = id_ctrl_decoder_decoded_invMatrixOutputs[29:28]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [2:0] id_ctrl_decoder_13 = id_ctrl_decoder_decoded_invMatrixOutputs[27:25]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_14 = id_ctrl_decoder_decoded_invMatrixOutputs[24]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [3:0] id_ctrl_decoder_15 = id_ctrl_decoder_decoded_invMatrixOutputs[23:20]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_16 = id_ctrl_decoder_decoded_invMatrixOutputs[19]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [4:0] id_ctrl_decoder_17 = id_ctrl_decoder_decoded_invMatrixOutputs[18:14]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_21 = id_ctrl_decoder_decoded_invMatrixOutputs[10]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_22 = id_ctrl_decoder_decoded_invMatrixOutputs[9]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_23 = id_ctrl_decoder_decoded_invMatrixOutputs[8]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_24 = id_ctrl_decoder_decoded_invMatrixOutputs[7]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [2:0] id_ctrl_decoder_25 = id_ctrl_decoder_decoded_invMatrixOutputs[6:4]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_26 = id_ctrl_decoder_decoded_invMatrixOutputs[3]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_27 = id_ctrl_decoder_decoded_invMatrixOutputs[2]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_28 = id_ctrl_decoder_decoded_invMatrixOutputs[1]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire  id_ctrl_decoder_29 = id_ctrl_decoder_decoded_invMatrixOutputs[0]; // @[src/main/scala/rocket/Decode.scala 53:77]
  wire [4:0] id_raddr2 = ibuf_io_inst_0_bits_inst_rs2; // @[src/main/scala/rocket/RocketCore.scala 298:72]
  wire [4:0] id_raddr1 = ibuf_io_inst_0_bits_inst_rs1; // @[src/main/scala/rocket/RocketCore.scala 298:72]
  wire [4:0] id_waddr = ibuf_io_inst_0_bits_inst_rd; // @[src/main/scala/rocket/RocketCore.scala 298:72]
  reg  id_reg_fence; // @[src/main/scala/rocket/RocketCore.scala 305:29]
  reg [63:0] rf_0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_1; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_2; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_3; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_4; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_5; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_6; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_7; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_8; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_9; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_10; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_11; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_12; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_13; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_14; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_15; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_16; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_17; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_18; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_19; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_20; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_21; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_22; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_23; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_24; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_25; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_26; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_27; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_28; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_29; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  reg [63:0] rf_30; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
  wire [4:0] _id_rs_T_3 = ~id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 1195:39]
  wire  line_1117_clock;
  wire  line_1117_reset;
  wire  line_1117_valid;
  reg  line_1117_valid_reg;
  wire  line_1118_clock;
  wire  line_1118_reset;
  wire  line_1118_valid;
  reg  line_1118_valid_reg;
  wire [63:0] _GEN_124 = 5'h1 == _id_rs_T_3 ? rf_1 : rf_0; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1119_clock;
  wire  line_1119_reset;
  wire  line_1119_valid;
  reg  line_1119_valid_reg;
  wire [63:0] _GEN_125 = 5'h2 == _id_rs_T_3 ? rf_2 : _GEN_124; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1120_clock;
  wire  line_1120_reset;
  wire  line_1120_valid;
  reg  line_1120_valid_reg;
  wire [63:0] _GEN_126 = 5'h3 == _id_rs_T_3 ? rf_3 : _GEN_125; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1121_clock;
  wire  line_1121_reset;
  wire  line_1121_valid;
  reg  line_1121_valid_reg;
  wire [63:0] _GEN_127 = 5'h4 == _id_rs_T_3 ? rf_4 : _GEN_126; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1122_clock;
  wire  line_1122_reset;
  wire  line_1122_valid;
  reg  line_1122_valid_reg;
  wire [63:0] _GEN_128 = 5'h5 == _id_rs_T_3 ? rf_5 : _GEN_127; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1123_clock;
  wire  line_1123_reset;
  wire  line_1123_valid;
  reg  line_1123_valid_reg;
  wire [63:0] _GEN_129 = 5'h6 == _id_rs_T_3 ? rf_6 : _GEN_128; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1124_clock;
  wire  line_1124_reset;
  wire  line_1124_valid;
  reg  line_1124_valid_reg;
  wire [63:0] _GEN_130 = 5'h7 == _id_rs_T_3 ? rf_7 : _GEN_129; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1125_clock;
  wire  line_1125_reset;
  wire  line_1125_valid;
  reg  line_1125_valid_reg;
  wire [63:0] _GEN_131 = 5'h8 == _id_rs_T_3 ? rf_8 : _GEN_130; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1126_clock;
  wire  line_1126_reset;
  wire  line_1126_valid;
  reg  line_1126_valid_reg;
  wire [63:0] _GEN_132 = 5'h9 == _id_rs_T_3 ? rf_9 : _GEN_131; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1127_clock;
  wire  line_1127_reset;
  wire  line_1127_valid;
  reg  line_1127_valid_reg;
  wire [63:0] _GEN_133 = 5'ha == _id_rs_T_3 ? rf_10 : _GEN_132; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1128_clock;
  wire  line_1128_reset;
  wire  line_1128_valid;
  reg  line_1128_valid_reg;
  wire [63:0] _GEN_134 = 5'hb == _id_rs_T_3 ? rf_11 : _GEN_133; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1129_clock;
  wire  line_1129_reset;
  wire  line_1129_valid;
  reg  line_1129_valid_reg;
  wire [63:0] _GEN_135 = 5'hc == _id_rs_T_3 ? rf_12 : _GEN_134; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1130_clock;
  wire  line_1130_reset;
  wire  line_1130_valid;
  reg  line_1130_valid_reg;
  wire [63:0] _GEN_136 = 5'hd == _id_rs_T_3 ? rf_13 : _GEN_135; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1131_clock;
  wire  line_1131_reset;
  wire  line_1131_valid;
  reg  line_1131_valid_reg;
  wire [63:0] _GEN_137 = 5'he == _id_rs_T_3 ? rf_14 : _GEN_136; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1132_clock;
  wire  line_1132_reset;
  wire  line_1132_valid;
  reg  line_1132_valid_reg;
  wire [63:0] _GEN_138 = 5'hf == _id_rs_T_3 ? rf_15 : _GEN_137; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1133_clock;
  wire  line_1133_reset;
  wire  line_1133_valid;
  reg  line_1133_valid_reg;
  wire [63:0] _GEN_139 = 5'h10 == _id_rs_T_3 ? rf_16 : _GEN_138; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1134_clock;
  wire  line_1134_reset;
  wire  line_1134_valid;
  reg  line_1134_valid_reg;
  wire [63:0] _GEN_140 = 5'h11 == _id_rs_T_3 ? rf_17 : _GEN_139; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1135_clock;
  wire  line_1135_reset;
  wire  line_1135_valid;
  reg  line_1135_valid_reg;
  wire [63:0] _GEN_141 = 5'h12 == _id_rs_T_3 ? rf_18 : _GEN_140; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1136_clock;
  wire  line_1136_reset;
  wire  line_1136_valid;
  reg  line_1136_valid_reg;
  wire [63:0] _GEN_142 = 5'h13 == _id_rs_T_3 ? rf_19 : _GEN_141; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1137_clock;
  wire  line_1137_reset;
  wire  line_1137_valid;
  reg  line_1137_valid_reg;
  wire [63:0] _GEN_143 = 5'h14 == _id_rs_T_3 ? rf_20 : _GEN_142; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1138_clock;
  wire  line_1138_reset;
  wire  line_1138_valid;
  reg  line_1138_valid_reg;
  wire [63:0] _GEN_144 = 5'h15 == _id_rs_T_3 ? rf_21 : _GEN_143; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1139_clock;
  wire  line_1139_reset;
  wire  line_1139_valid;
  reg  line_1139_valid_reg;
  wire [63:0] _GEN_145 = 5'h16 == _id_rs_T_3 ? rf_22 : _GEN_144; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1140_clock;
  wire  line_1140_reset;
  wire  line_1140_valid;
  reg  line_1140_valid_reg;
  wire [63:0] _GEN_146 = 5'h17 == _id_rs_T_3 ? rf_23 : _GEN_145; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1141_clock;
  wire  line_1141_reset;
  wire  line_1141_valid;
  reg  line_1141_valid_reg;
  wire [63:0] _GEN_147 = 5'h18 == _id_rs_T_3 ? rf_24 : _GEN_146; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1142_clock;
  wire  line_1142_reset;
  wire  line_1142_valid;
  reg  line_1142_valid_reg;
  wire [63:0] _GEN_148 = 5'h19 == _id_rs_T_3 ? rf_25 : _GEN_147; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1143_clock;
  wire  line_1143_reset;
  wire  line_1143_valid;
  reg  line_1143_valid_reg;
  wire [63:0] _GEN_149 = 5'h1a == _id_rs_T_3 ? rf_26 : _GEN_148; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1144_clock;
  wire  line_1144_reset;
  wire  line_1144_valid;
  reg  line_1144_valid_reg;
  wire [63:0] _GEN_150 = 5'h1b == _id_rs_T_3 ? rf_27 : _GEN_149; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1145_clock;
  wire  line_1145_reset;
  wire  line_1145_valid;
  reg  line_1145_valid_reg;
  wire [63:0] _GEN_151 = 5'h1c == _id_rs_T_3 ? rf_28 : _GEN_150; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1146_clock;
  wire  line_1146_reset;
  wire  line_1146_valid;
  reg  line_1146_valid_reg;
  wire [63:0] _GEN_152 = 5'h1d == _id_rs_T_3 ? rf_29 : _GEN_151; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1147_clock;
  wire  line_1147_reset;
  wire  line_1147_valid;
  reg  line_1147_valid_reg;
  wire [63:0] _GEN_153 = 5'h1e == _id_rs_T_3 ? rf_30 : _GEN_152; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire [4:0] _id_rs_T_8 = ~id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 1195:39]
  wire  line_1148_clock;
  wire  line_1148_reset;
  wire  line_1148_valid;
  reg  line_1148_valid_reg;
  wire  line_1149_clock;
  wire  line_1149_reset;
  wire  line_1149_valid;
  reg  line_1149_valid_reg;
  wire [63:0] _GEN_155 = 5'h1 == _id_rs_T_8 ? rf_1 : rf_0; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1150_clock;
  wire  line_1150_reset;
  wire  line_1150_valid;
  reg  line_1150_valid_reg;
  wire [63:0] _GEN_156 = 5'h2 == _id_rs_T_8 ? rf_2 : _GEN_155; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1151_clock;
  wire  line_1151_reset;
  wire  line_1151_valid;
  reg  line_1151_valid_reg;
  wire [63:0] _GEN_157 = 5'h3 == _id_rs_T_8 ? rf_3 : _GEN_156; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1152_clock;
  wire  line_1152_reset;
  wire  line_1152_valid;
  reg  line_1152_valid_reg;
  wire [63:0] _GEN_158 = 5'h4 == _id_rs_T_8 ? rf_4 : _GEN_157; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1153_clock;
  wire  line_1153_reset;
  wire  line_1153_valid;
  reg  line_1153_valid_reg;
  wire [63:0] _GEN_159 = 5'h5 == _id_rs_T_8 ? rf_5 : _GEN_158; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1154_clock;
  wire  line_1154_reset;
  wire  line_1154_valid;
  reg  line_1154_valid_reg;
  wire [63:0] _GEN_160 = 5'h6 == _id_rs_T_8 ? rf_6 : _GEN_159; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1155_clock;
  wire  line_1155_reset;
  wire  line_1155_valid;
  reg  line_1155_valid_reg;
  wire [63:0] _GEN_161 = 5'h7 == _id_rs_T_8 ? rf_7 : _GEN_160; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1156_clock;
  wire  line_1156_reset;
  wire  line_1156_valid;
  reg  line_1156_valid_reg;
  wire [63:0] _GEN_162 = 5'h8 == _id_rs_T_8 ? rf_8 : _GEN_161; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1157_clock;
  wire  line_1157_reset;
  wire  line_1157_valid;
  reg  line_1157_valid_reg;
  wire [63:0] _GEN_163 = 5'h9 == _id_rs_T_8 ? rf_9 : _GEN_162; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1158_clock;
  wire  line_1158_reset;
  wire  line_1158_valid;
  reg  line_1158_valid_reg;
  wire [63:0] _GEN_164 = 5'ha == _id_rs_T_8 ? rf_10 : _GEN_163; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1159_clock;
  wire  line_1159_reset;
  wire  line_1159_valid;
  reg  line_1159_valid_reg;
  wire [63:0] _GEN_165 = 5'hb == _id_rs_T_8 ? rf_11 : _GEN_164; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1160_clock;
  wire  line_1160_reset;
  wire  line_1160_valid;
  reg  line_1160_valid_reg;
  wire [63:0] _GEN_166 = 5'hc == _id_rs_T_8 ? rf_12 : _GEN_165; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1161_clock;
  wire  line_1161_reset;
  wire  line_1161_valid;
  reg  line_1161_valid_reg;
  wire [63:0] _GEN_167 = 5'hd == _id_rs_T_8 ? rf_13 : _GEN_166; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1162_clock;
  wire  line_1162_reset;
  wire  line_1162_valid;
  reg  line_1162_valid_reg;
  wire [63:0] _GEN_168 = 5'he == _id_rs_T_8 ? rf_14 : _GEN_167; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1163_clock;
  wire  line_1163_reset;
  wire  line_1163_valid;
  reg  line_1163_valid_reg;
  wire [63:0] _GEN_169 = 5'hf == _id_rs_T_8 ? rf_15 : _GEN_168; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1164_clock;
  wire  line_1164_reset;
  wire  line_1164_valid;
  reg  line_1164_valid_reg;
  wire [63:0] _GEN_170 = 5'h10 == _id_rs_T_8 ? rf_16 : _GEN_169; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1165_clock;
  wire  line_1165_reset;
  wire  line_1165_valid;
  reg  line_1165_valid_reg;
  wire [63:0] _GEN_171 = 5'h11 == _id_rs_T_8 ? rf_17 : _GEN_170; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1166_clock;
  wire  line_1166_reset;
  wire  line_1166_valid;
  reg  line_1166_valid_reg;
  wire [63:0] _GEN_172 = 5'h12 == _id_rs_T_8 ? rf_18 : _GEN_171; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1167_clock;
  wire  line_1167_reset;
  wire  line_1167_valid;
  reg  line_1167_valid_reg;
  wire [63:0] _GEN_173 = 5'h13 == _id_rs_T_8 ? rf_19 : _GEN_172; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1168_clock;
  wire  line_1168_reset;
  wire  line_1168_valid;
  reg  line_1168_valid_reg;
  wire [63:0] _GEN_174 = 5'h14 == _id_rs_T_8 ? rf_20 : _GEN_173; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1169_clock;
  wire  line_1169_reset;
  wire  line_1169_valid;
  reg  line_1169_valid_reg;
  wire [63:0] _GEN_175 = 5'h15 == _id_rs_T_8 ? rf_21 : _GEN_174; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1170_clock;
  wire  line_1170_reset;
  wire  line_1170_valid;
  reg  line_1170_valid_reg;
  wire [63:0] _GEN_176 = 5'h16 == _id_rs_T_8 ? rf_22 : _GEN_175; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1171_clock;
  wire  line_1171_reset;
  wire  line_1171_valid;
  reg  line_1171_valid_reg;
  wire [63:0] _GEN_177 = 5'h17 == _id_rs_T_8 ? rf_23 : _GEN_176; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1172_clock;
  wire  line_1172_reset;
  wire  line_1172_valid;
  reg  line_1172_valid_reg;
  wire [63:0] _GEN_178 = 5'h18 == _id_rs_T_8 ? rf_24 : _GEN_177; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1173_clock;
  wire  line_1173_reset;
  wire  line_1173_valid;
  reg  line_1173_valid_reg;
  wire [63:0] _GEN_179 = 5'h19 == _id_rs_T_8 ? rf_25 : _GEN_178; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1174_clock;
  wire  line_1174_reset;
  wire  line_1174_valid;
  reg  line_1174_valid_reg;
  wire [63:0] _GEN_180 = 5'h1a == _id_rs_T_8 ? rf_26 : _GEN_179; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1175_clock;
  wire  line_1175_reset;
  wire  line_1175_valid;
  reg  line_1175_valid_reg;
  wire [63:0] _GEN_181 = 5'h1b == _id_rs_T_8 ? rf_27 : _GEN_180; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1176_clock;
  wire  line_1176_reset;
  wire  line_1176_valid;
  reg  line_1176_valid_reg;
  wire [63:0] _GEN_182 = 5'h1c == _id_rs_T_8 ? rf_28 : _GEN_181; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1177_clock;
  wire  line_1177_reset;
  wire  line_1177_valid;
  reg  line_1177_valid_reg;
  wire [63:0] _GEN_183 = 5'h1d == _id_rs_T_8 ? rf_29 : _GEN_182; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  line_1178_clock;
  wire  line_1178_reset;
  wire  line_1178_valid;
  reg  line_1178_valid_reg;
  wire [63:0] _GEN_184 = 5'h1e == _id_rs_T_8 ? rf_30 : _GEN_183; // @[src/main/scala/rocket/RocketCore.scala 1201:{25,25}]
  wire  _id_csr_en_T = id_ctrl_decoder_25 == 3'h6; // @[src/main/scala/util/package.scala 16:47]
  wire  _id_csr_en_T_1 = id_ctrl_decoder_25 == 3'h7; // @[src/main/scala/util/package.scala 16:47]
  wire  _id_csr_en_T_2 = id_ctrl_decoder_25 == 3'h5; // @[src/main/scala/util/package.scala 16:47]
  wire  _id_csr_en_T_3 = _id_csr_en_T | _id_csr_en_T_1; // @[src/main/scala/util/package.scala 73:59]
  wire  id_csr_en = _id_csr_en_T | _id_csr_en_T_1 | _id_csr_en_T_2; // @[src/main/scala/util/package.scala 73:59]
  wire  id_system_insn = id_ctrl_decoder_25 == 3'h4; // @[src/main/scala/rocket/RocketCore.scala 315:36]
  wire  id_csr_ren = _id_csr_en_T_3 & ibuf_io_inst_0_bits_inst_rs1 == 5'h0; // @[src/main/scala/rocket/RocketCore.scala 316:54]
  wire  _id_csr_flush_T = ~id_csr_ren; // @[src/main/scala/rocket/RocketCore.scala 318:54]
  wire  id_csr_flush = id_system_insn | id_csr_en & ~id_csr_ren & csr_io_decode_0_write_flush; // @[src/main/scala/rocket/RocketCore.scala 318:37]
  wire  _id_illegal_insn_T_4 = (id_ctrl_decoder_22 | id_ctrl_decoder_23) & ~csr_io_status_isa[12]; // @[src/main/scala/rocket/RocketCore.scala 322:34]
  wire  _id_illegal_insn_T_5 = ~id_ctrl_decoder_0 | _id_illegal_insn_T_4; // @[src/main/scala/rocket/RocketCore.scala 321:40]
  wire  _id_illegal_insn_T_8 = id_ctrl_decoder_28 & ~csr_io_status_isa[0]; // @[src/main/scala/rocket/RocketCore.scala 323:17]
  wire  _id_illegal_insn_T_9 = _id_illegal_insn_T_5 | _id_illegal_insn_T_8; // @[src/main/scala/rocket/RocketCore.scala 322:65]
  wire  _id_illegal_insn_T_11 = id_ctrl_decoder_1 & csr_io_decode_0_fp_illegal; // @[src/main/scala/rocket/RocketCore.scala 324:16]
  wire  _id_illegal_insn_T_12 = _id_illegal_insn_T_9 | _id_illegal_insn_T_11; // @[src/main/scala/rocket/RocketCore.scala 323:48]
  wire  _id_illegal_insn_T_15 = id_ctrl_decoder_29 & ~csr_io_status_isa[3]; // @[src/main/scala/rocket/RocketCore.scala 325:16]
  wire  _id_illegal_insn_T_16 = _id_illegal_insn_T_12 | _id_illegal_insn_T_15; // @[src/main/scala/rocket/RocketCore.scala 324:70]
  wire  _id_illegal_insn_T_18 = ~csr_io_status_isa[2]; // @[src/main/scala/rocket/RocketCore.scala 326:33]
  wire  _id_illegal_insn_T_19 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2]; // @[src/main/scala/rocket/RocketCore.scala 326:30]
  wire  _id_illegal_insn_T_20 = _id_illegal_insn_T_16 | _id_illegal_insn_T_19; // @[src/main/scala/rocket/RocketCore.scala 325:47]
  wire  _id_illegal_insn_T_27 = id_ctrl_decoder_2 & csr_io_decode_0_rocc_illegal; // @[src/main/scala/rocket/RocketCore.scala 330:18]
  wire  _id_illegal_insn_T_28 = _id_illegal_insn_T_20 | _id_illegal_insn_T_27; // @[src/main/scala/rocket/RocketCore.scala 329:37]
  wire  _id_illegal_insn_T_32 = id_csr_en & (csr_io_decode_0_read_illegal | _id_csr_flush_T &
    csr_io_decode_0_write_illegal); // @[src/main/scala/rocket/RocketCore.scala 331:15]
  wire  _id_illegal_insn_T_33 = _id_illegal_insn_T_28 | _id_illegal_insn_T_32; // @[src/main/scala/rocket/RocketCore.scala 330:51]
  wire  _id_illegal_insn_T_36 = ~ibuf_io_inst_0_bits_rvc & (id_system_insn & csr_io_decode_0_system_illegal); // @[src/main/scala/rocket/RocketCore.scala 332:31]
  wire  id_illegal_insn = _id_illegal_insn_T_33 | _id_illegal_insn_T_36; // @[src/main/scala/rocket/RocketCore.scala 331:99]
  wire  id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26]; // @[src/main/scala/rocket/RocketCore.scala 338:29]
  wire  id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25]; // @[src/main/scala/rocket/RocketCore.scala 339:29]
  wire [3:0] id_fence_succ = ibuf_io_inst_0_bits_inst_bits[23:20]; // @[src/main/scala/rocket/RocketCore.scala 341:33]
  wire  id_fence_next = id_ctrl_decoder_27 | id_ctrl_decoder_28 & id_amo_aq; // @[src/main/scala/rocket/RocketCore.scala 342:37]
  wire  id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid; // @[src/main/scala/rocket/RocketCore.scala 343:38]
  wire  _T = ~id_mem_busy; // @[src/main/scala/rocket/RocketCore.scala 344:9]
  wire  line_1179_clock;
  wire  line_1179_reset;
  wire  line_1179_valid;
  reg  line_1179_valid_reg;
  wire  _GEN_185 = ~id_mem_busy ? 1'h0 : id_reg_fence; // @[src/main/scala/rocket/RocketCore.scala 344:23 305:29 344:38]
  wire  id_do_fence = id_mem_busy & (id_ctrl_decoder_28 & id_amo_rl | id_ctrl_decoder_26 | id_reg_fence & (
    id_ctrl_decoder_16 | id_ctrl_decoder_2)); // @[src/main/scala/rocket/RocketCore.scala 349:17]
  wire  id_xcpt = csr_io_interrupt | ibuf_io_inst_0_bits_xcpt0_pf_inst | ibuf_io_inst_0_bits_xcpt0_ae_inst |
    ibuf_io_inst_0_bits_xcpt1_pf_inst | ibuf_io_inst_0_bits_xcpt1_gf_inst | ibuf_io_inst_0_bits_xcpt1_ae_inst |
    id_illegal_insn; // @[src/main/scala/rocket/RocketCore.scala 1152:26]
  wire [4:0] _T_11 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 5'h1 : 5'h2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_12 = ibuf_io_inst_0_bits_xcpt1_gf_inst ? 5'h14 : _T_11; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_13 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 5'hc : _T_12; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_14 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 5'h1 : _T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_16 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 5'hc : _T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] ex_waddr = ex_reg_inst[11:7]; // @[src/main/scala/rocket/RocketCore.scala 390:29]
  wire [4:0] mem_waddr = mem_reg_inst[11:7]; // @[src/main/scala/rocket/RocketCore.scala 391:31]
  wire [4:0] wb_waddr = wb_reg_inst[11:7]; // @[src/main/scala/rocket/RocketCore.scala 392:29]
  wire  _T_29 = ex_reg_valid & ex_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 395:19]
  wire  _T_30 = mem_reg_valid & mem_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 396:20]
  wire  _T_32 = mem_reg_valid & mem_ctrl_wxd & ~mem_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 396:36]
  wire  id_bypass_src_0_0 = 5'h0 == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 398:82]
  wire  id_bypass_src_0_1 = _T_29 & ex_waddr == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  wire  id_bypass_src_0_2 = _T_32 & mem_waddr == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  wire  id_bypass_src_0_3 = _T_30 & mem_waddr == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  wire  id_bypass_src_1_0 = 5'h0 == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 398:82]
  wire  id_bypass_src_1_1 = _T_29 & ex_waddr == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  wire  id_bypass_src_1_2 = _T_32 & mem_waddr == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  wire  id_bypass_src_1_3 = _T_30 & mem_waddr == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 398:74]
  reg  ex_reg_rs_bypass_0; // @[src/main/scala/rocket/RocketCore.scala 402:29]
  reg  ex_reg_rs_bypass_1; // @[src/main/scala/rocket/RocketCore.scala 402:29]
  reg [1:0] ex_reg_rs_lsb_0; // @[src/main/scala/rocket/RocketCore.scala 403:26]
  reg [1:0] ex_reg_rs_lsb_1; // @[src/main/scala/rocket/RocketCore.scala 403:26]
  reg [61:0] ex_reg_rs_msb_0; // @[src/main/scala/rocket/RocketCore.scala 404:26]
  reg [61:0] ex_reg_rs_msb_1; // @[src/main/scala/rocket/RocketCore.scala 404:26]
  wire [63:0] _ex_rs_T_1 = ex_reg_rs_lsb_0 == 2'h1 ? mem_reg_wdata : 64'h0; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_3 = ex_reg_rs_lsb_0 == 2'h2 ? wb_reg_wdata : _ex_rs_T_1; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_5 = ex_reg_rs_lsb_0 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_3; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_6 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0}; // @[src/main/scala/rocket/RocketCore.scala 406:69]
  wire [63:0] ex_rs_0 = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[src/main/scala/rocket/RocketCore.scala 406:14]
  wire [63:0] _ex_rs_T_8 = ex_reg_rs_lsb_1 == 2'h1 ? mem_reg_wdata : 64'h0; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_10 = ex_reg_rs_lsb_1 == 2'h2 ? wb_reg_wdata : _ex_rs_T_8; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_12 = ex_reg_rs_lsb_1 == 2'h3 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_10; // @[src/main/scala/util/package.scala 33:76]
  wire [63:0] _ex_rs_T_13 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1}; // @[src/main/scala/rocket/RocketCore.scala 406:69]
  wire [63:0] ex_rs_1 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[src/main/scala/rocket/RocketCore.scala 406:14]
  wire  _ex_imm_sign_T = ex_ctrl_sel_imm == 3'h5; // @[src/main/scala/rocket/RocketCore.scala 1217:24]
  wire  _ex_imm_sign_T_2 = ex_reg_inst[31]; // @[src/main/scala/rocket/RocketCore.scala 1217:49]
  wire  ex_imm_sign = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[src/main/scala/rocket/RocketCore.scala 1217:19]
  wire  _ex_imm_b30_20_T = ex_ctrl_sel_imm == 3'h2; // @[src/main/scala/rocket/RocketCore.scala 1218:26]
  wire [10:0] _ex_imm_b30_20_T_2 = ex_reg_inst[30:20]; // @[src/main/scala/rocket/RocketCore.scala 1218:49]
  wire [7:0] _ex_imm_b19_12_T_4 = ex_reg_inst[19:12]; // @[src/main/scala/rocket/RocketCore.scala 1219:73]
  wire  _ex_imm_b11_T_2 = _ex_imm_b30_20_T | _ex_imm_sign_T; // @[src/main/scala/rocket/RocketCore.scala 1220:33]
  wire  _ex_imm_b11_T_5 = ex_reg_inst[20]; // @[src/main/scala/rocket/RocketCore.scala 1221:44]
  wire  _ex_imm_b11_T_6 = ex_ctrl_sel_imm == 3'h1; // @[src/main/scala/rocket/RocketCore.scala 1222:23]
  wire  _ex_imm_b11_T_8 = ex_reg_inst[7]; // @[src/main/scala/rocket/RocketCore.scala 1222:43]
  wire  _ex_imm_b11_T_9 = ex_ctrl_sel_imm == 3'h1 ? $signed(_ex_imm_b11_T_8) : $signed(ex_imm_sign); // @[src/main/scala/rocket/RocketCore.scala 1222:18]
  wire  _ex_imm_b11_T_10 = ex_ctrl_sel_imm == 3'h3 ? $signed(_ex_imm_b11_T_5) : $signed(_ex_imm_b11_T_9); // @[src/main/scala/rocket/RocketCore.scala 1221:18]
  wire [5:0] ex_imm_b10_5 = _ex_imm_b11_T_2 ? 6'h0 : ex_reg_inst[30:25]; // @[src/main/scala/rocket/RocketCore.scala 1223:20]
  wire  _ex_imm_b4_1_T_1 = ex_ctrl_sel_imm == 3'h0; // @[src/main/scala/rocket/RocketCore.scala 1225:24]
  wire [3:0] _ex_imm_b4_1_T_8 = _ex_imm_sign_T ? ex_reg_inst[19:16] : ex_reg_inst[24:21]; // @[src/main/scala/rocket/RocketCore.scala 1226:19]
  wire [3:0] _ex_imm_b4_1_T_9 = ex_ctrl_sel_imm == 3'h0 | _ex_imm_b11_T_6 ? ex_reg_inst[11:8] : _ex_imm_b4_1_T_8; // @[src/main/scala/rocket/RocketCore.scala 1225:19]
  wire [3:0] ex_imm_b4_1 = _ex_imm_b30_20_T ? 4'h0 : _ex_imm_b4_1_T_9; // @[src/main/scala/rocket/RocketCore.scala 1224:19]
  wire  _ex_imm_b0_T_6 = _ex_imm_sign_T & ex_reg_inst[15]; // @[src/main/scala/rocket/RocketCore.scala 1229:17]
  wire  _ex_imm_b0_T_7 = ex_ctrl_sel_imm == 3'h4 ? ex_reg_inst[20] : _ex_imm_b0_T_6; // @[src/main/scala/rocket/RocketCore.scala 1228:17]
  wire  ex_imm_b0 = _ex_imm_b4_1_T_1 ? ex_reg_inst[7] : _ex_imm_b0_T_7; // @[src/main/scala/rocket/RocketCore.scala 1227:17]
  wire  ex_imm_hi_lo_lo = _ex_imm_b30_20_T | _ex_imm_sign_T ? $signed(1'sh0) : $signed(_ex_imm_b11_T_10); // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [7:0] ex_imm_hi_lo_hi = ex_ctrl_sel_imm != 3'h2 & ex_ctrl_sel_imm != 3'h3 ? $signed({8{ex_imm_sign}}) : $signed(
    _ex_imm_b19_12_T_4); // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [10:0] ex_imm_hi_hi_lo = ex_ctrl_sel_imm == 3'h2 ? $signed(_ex_imm_b30_20_T_2) : $signed({11{ex_imm_sign}}); // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire  ex_imm_hi_hi_hi = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [31:0] ex_imm = {ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_b10_5,ex_imm_b4_1,
    ex_imm_b0}; // @[src/main/scala/rocket/RocketCore.scala 1231:53]
  wire [63:0] _ex_op1_T = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[src/main/scala/rocket/RocketCore.scala 409:24]
  wire [39:0] _ex_op1_T_1 = ex_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 410:24]
  wire [63:0] _ex_op1_T_3 = 2'h1 == ex_ctrl_sel_alu1 ? $signed(_ex_op1_T) : $signed(64'sh0); // @[src/main/scala/rocket/RocketCore.scala 408:48]
  wire [63:0] _ex_op2_T = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[src/main/scala/rocket/RocketCore.scala 412:24]
  wire [3:0] _ex_op2_T_1 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[src/main/scala/rocket/RocketCore.scala 414:19]
  wire [63:0] _ex_op2_T_3 = 2'h2 == ex_ctrl_sel_alu2 ? $signed(_ex_op2_T) : $signed(64'sh0); // @[src/main/scala/rocket/RocketCore.scala 411:48]
  wire [63:0] _ex_op2_T_5 = 2'h3 == ex_ctrl_sel_alu2 ? $signed({{32{ex_imm[31]}},ex_imm}) : $signed(_ex_op2_T_3); // @[src/main/scala/rocket/RocketCore.scala 411:48]
  wire  _T_140 = id_raddr1 != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 840:55]
  wire  _T_141 = id_ctrl_decoder_7 & id_raddr1 != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 840:42]
  wire  _data_hazard_ex_T = id_raddr1 == ex_waddr; // @[src/main/scala/rocket/RocketCore.scala 860:70]
  wire  _T_142 = id_raddr2 != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 841:55]
  wire  _T_143 = id_ctrl_decoder_6 & id_raddr2 != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 841:42]
  wire  _data_hazard_ex_T_2 = id_raddr2 == ex_waddr; // @[src/main/scala/rocket/RocketCore.scala 860:70]
  wire  _T_145 = id_ctrl_decoder_24 & id_waddr != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 842:42]
  wire  _data_hazard_ex_T_4 = id_waddr == ex_waddr; // @[src/main/scala/rocket/RocketCore.scala 860:70]
  wire  _data_hazard_ex_T_7 = _T_141 & _data_hazard_ex_T | _T_143 & _data_hazard_ex_T_2 | _T_145 & _data_hazard_ex_T_4; // @[src/main/scala/rocket/RocketCore.scala 1161:50]
  wire  data_hazard_ex = ex_ctrl_wxd & _data_hazard_ex_T_7; // @[src/main/scala/rocket/RocketCore.scala 860:36]
  wire  ex_cannot_bypass = ex_ctrl_csr != 3'h0 | ex_ctrl_jalr | ex_ctrl_mem | ex_ctrl_mul | ex_ctrl_div | ex_ctrl_fp |
    ex_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 859:123]
  wire  id_ex_hazard = ex_reg_valid & (data_hazard_ex & ex_cannot_bypass); // @[src/main/scala/rocket/RocketCore.scala 862:35]
  wire  _data_hazard_mem_T = id_raddr1 == mem_waddr; // @[src/main/scala/rocket/RocketCore.scala 869:72]
  wire  _data_hazard_mem_T_2 = id_raddr2 == mem_waddr; // @[src/main/scala/rocket/RocketCore.scala 869:72]
  wire  _data_hazard_mem_T_4 = id_waddr == mem_waddr; // @[src/main/scala/rocket/RocketCore.scala 869:72]
  wire  _data_hazard_mem_T_7 = _T_141 & _data_hazard_mem_T | _T_143 & _data_hazard_mem_T_2 | _T_145 &
    _data_hazard_mem_T_4; // @[src/main/scala/rocket/RocketCore.scala 1161:50]
  wire  data_hazard_mem = mem_ctrl_wxd & _data_hazard_mem_T_7; // @[src/main/scala/rocket/RocketCore.scala 869:38]
  wire  mem_cannot_bypass = mem_ctrl_csr != 3'h0 | mem_ctrl_mem & mem_reg_slow_bypass | mem_ctrl_mul | mem_ctrl_div |
    mem_ctrl_fp | mem_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 868:131]
  wire  id_mem_hazard = mem_reg_valid & (data_hazard_mem & mem_cannot_bypass); // @[src/main/scala/rocket/RocketCore.scala 871:37]
  wire  _data_hazard_wb_T = id_raddr1 == wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 875:70]
  wire  _data_hazard_wb_T_2 = id_raddr2 == wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 875:70]
  wire  _data_hazard_wb_T_4 = id_waddr == wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 875:70]
  wire  _data_hazard_wb_T_7 = _T_141 & _data_hazard_wb_T | _T_143 & _data_hazard_wb_T_2 | _T_145 & _data_hazard_wb_T_4; // @[src/main/scala/rocket/RocketCore.scala 1161:50]
  wire  data_hazard_wb = wb_ctrl_wxd & _data_hazard_wb_T_7; // @[src/main/scala/rocket/RocketCore.scala 875:36]
  wire  wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid; // @[src/main/scala/rocket/RocketCore.scala 538:36]
  wire  wb_set_sboard = wb_ctrl_div | wb_dcache_miss | wb_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 696:53]
  wire  id_wb_hazard = wb_reg_valid & (data_hazard_wb & wb_set_sboard); // @[src/main/scala/rocket/RocketCore.scala 877:35]
  reg [31:0] reg_r; // @[src/main/scala/rocket/RocketCore.scala 1179:32]
  wire [31:0] r = {reg_r[31:1], 1'h0}; // @[src/main/scala/rocket/RocketCore.scala 1180:43]
  wire [31:0] _id_sboard_hazard_T = r >> id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 1176:35]
  wire  dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data; // @[src/main/scala/rocket/RocketCore.scala 707:44]
  wire  dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 708:42]
  wire  dmem_resp_xpu = ~io_dmem_resp_bits_tag[0]; // @[src/main/scala/rocket/RocketCore.scala 704:23]
  wire  _T_134 = dmem_resp_replay & dmem_resp_xpu; // @[src/main/scala/rocket/RocketCore.scala 730:26]
  wire  _ll_wen_T = div_io_resp_ready & div_io_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  ll_wen = dmem_resp_replay & dmem_resp_xpu | _ll_wen_T; // @[src/main/scala/rocket/RocketCore.scala 730:44 735:12 713:27]
  wire [4:0] dmem_resp_waddr = io_dmem_resp_bits_tag[5:1]; // @[src/main/scala/rocket/RocketCore.scala 706:46]
  wire [4:0] ll_waddr = dmem_resp_replay & dmem_resp_xpu ? dmem_resp_waddr : div_io_resp_bits_tag; // @[src/main/scala/rocket/RocketCore.scala 730:44 734:14 712:29]
  wire  _id_sboard_hazard_T_3 = ll_wen & ll_waddr == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 852:58]
  wire  _id_sboard_hazard_T_5 = _id_sboard_hazard_T[0] & ~_id_sboard_hazard_T_3; // @[src/main/scala/rocket/RocketCore.scala 855:77]
  wire [31:0] _id_sboard_hazard_T_7 = r >> id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 1176:35]
  wire  _id_sboard_hazard_T_10 = ll_wen & ll_waddr == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 852:58]
  wire  _id_sboard_hazard_T_12 = _id_sboard_hazard_T_7[0] & ~_id_sboard_hazard_T_10; // @[src/main/scala/rocket/RocketCore.scala 855:77]
  wire [31:0] _id_sboard_hazard_T_14 = r >> id_waddr; // @[src/main/scala/rocket/RocketCore.scala 1176:35]
  wire  _id_sboard_hazard_T_17 = ll_wen & ll_waddr == id_waddr; // @[src/main/scala/rocket/RocketCore.scala 852:58]
  wire  _id_sboard_hazard_T_19 = _id_sboard_hazard_T_14[0] & ~_id_sboard_hazard_T_17; // @[src/main/scala/rocket/RocketCore.scala 855:77]
  wire  id_sboard_hazard = _T_141 & _id_sboard_hazard_T_5 | _T_143 & _id_sboard_hazard_T_12 | _T_145 &
    _id_sboard_hazard_T_19; // @[src/main/scala/rocket/RocketCore.scala 1161:50]
  wire  _ctrl_stalld_T_5 = csr_io_singleStep & (ex_reg_valid | mem_reg_valid | wb_reg_valid); // @[src/main/scala/rocket/RocketCore.scala 899:23]
  wire  _ctrl_stalld_T_6 = id_ex_hazard | id_mem_hazard | id_wb_hazard | id_sboard_hazard | _ctrl_stalld_T_5; // @[src/main/scala/rocket/RocketCore.scala 898:71]
  reg  dcache_blocked_blocked; // @[src/main/scala/rocket/RocketCore.scala 890:22]
  wire  _dcache_blocked_T = ~io_dmem_perf_grant; // @[src/main/scala/rocket/RocketCore.scala 892:16]
  wire  dcache_blocked = dcache_blocked_blocked & ~io_dmem_perf_grant; // @[src/main/scala/rocket/RocketCore.scala 892:13]
  wire  _ctrl_stalld_T_13 = id_ctrl_decoder_16 & dcache_blocked; // @[src/main/scala/rocket/RocketCore.scala 902:17]
  wire  _ctrl_stalld_T_14 = _ctrl_stalld_T_6 | _ctrl_stalld_T_13; // @[src/main/scala/rocket/RocketCore.scala 901:32]
  reg  rocc_blocked; // @[src/main/scala/rocket/RocketCore.scala 894:25]
  wire  _ctrl_stalld_T_15 = id_ctrl_decoder_2 & rocc_blocked; // @[src/main/scala/rocket/RocketCore.scala 903:18]
  wire  _ctrl_stalld_T_16 = _ctrl_stalld_T_14 | _ctrl_stalld_T_15; // @[src/main/scala/rocket/RocketCore.scala 902:35]
  wire  wb_wxd = wb_reg_valid & wb_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 695:29]
  wire  _ctrl_stalld_T_17 = ~wb_wxd; // @[src/main/scala/rocket/RocketCore.scala 904:65]
  wire  _ctrl_stalld_T_22 = id_ctrl_decoder_23 & (~(div_io_req_ready | div_io_resp_valid & ~wb_wxd) | div_io_req_valid); // @[src/main/scala/rocket/RocketCore.scala 904:17]
  wire  _ctrl_stalld_T_23 = _ctrl_stalld_T_16 | _ctrl_stalld_T_22; // @[src/main/scala/rocket/RocketCore.scala 903:34]
  wire  _ctrl_stalld_T_26 = _ctrl_stalld_T_23 | id_do_fence; // @[src/main/scala/rocket/RocketCore.scala 905:15]
  wire  _ctrl_stalld_T_27 = _ctrl_stalld_T_26 | csr_io_csr_stall; // @[src/main/scala/rocket/RocketCore.scala 906:17]
  wire  ctrl_stalld = _ctrl_stalld_T_27 | id_reg_pause; // @[src/main/scala/rocket/RocketCore.scala 907:22]
  wire  ctrl_killd = ~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay | take_pc_mem_wb | ctrl_stalld |
    csr_io_interrupt; // @[src/main/scala/rocket/RocketCore.scala 910:104]
  wire  _ex_reg_valid_T = ~ctrl_killd; // @[src/main/scala/rocket/RocketCore.scala 468:19]
  wire  _ex_reg_replay_T = ~take_pc_mem_wb; // @[src/main/scala/rocket/RocketCore.scala 469:20]
  wire  _ex_reg_replay_T_1 = ~take_pc_mem_wb & ibuf_io_inst_0_valid; // @[src/main/scala/rocket/RocketCore.scala 469:29]
  wire  line_1180_clock;
  wire  line_1180_reset;
  wire  line_1180_valid;
  reg  line_1180_valid_reg;
  wire  _T_36 = id_ctrl_decoder_27 & id_fence_succ == 4'h0; // @[src/main/scala/rocket/RocketCore.scala 477:25]
  wire  line_1181_clock;
  wire  line_1181_reset;
  wire  line_1181_valid;
  reg  line_1181_valid_reg;
  wire  _GEN_186 = id_ctrl_decoder_27 & id_fence_succ == 4'h0 | id_reg_pause; // @[src/main/scala/rocket/RocketCore.scala 132:25 477:{51,66}]
  wire  line_1182_clock;
  wire  line_1182_reset;
  wire  line_1182_valid;
  reg  line_1182_valid_reg;
  wire  _GEN_187 = id_fence_next | _GEN_185; // @[src/main/scala/rocket/RocketCore.scala 478:{26,41}]
  wire  line_1183_clock;
  wire  line_1183_reset;
  wire  line_1183_valid;
  reg  line_1183_valid_reg;
  wire [2:0] _T_37 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_gf_inst,
    ibuf_io_inst_0_bits_xcpt1_ae_inst}; // @[src/main/scala/rocket/RocketCore.scala 484:22]
  wire  _T_38 = |_T_37; // @[src/main/scala/rocket/RocketCore.scala 484:29]
  wire  line_1184_clock;
  wire  line_1184_reset;
  wire  line_1184_valid;
  reg  line_1184_valid_reg;
  wire  _GEN_190 = |_T_37 | ibuf_io_inst_0_bits_rvc; // @[src/main/scala/rocket/RocketCore.scala 475:16 484:34 487:20]
  wire [2:0] _T_39 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,1'h0,ibuf_io_inst_0_bits_xcpt0_ae_inst}; // @[src/main/scala/rocket/RocketCore.scala 489:40]
  wire  _T_40 = |_T_39; // @[src/main/scala/rocket/RocketCore.scala 489:47]
  wire  line_1185_clock;
  wire  line_1185_reset;
  wire  line_1185_valid;
  reg  line_1185_valid_reg;
  wire  _GEN_194 = id_xcpt | id_ctrl_decoder_14; // @[src/main/scala/rocket/RocketCore.scala 474:13 479:20 481:22]
  wire  _T_42 = id_ctrl_decoder_17 == 5'h14; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_43 = id_ctrl_decoder_17 == 5'h15; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_44 = id_ctrl_decoder_17 == 5'h16; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_45 = id_ctrl_decoder_17 == 5'h5; // @[src/main/scala/util/package.scala 16:47]
  wire  _T_48 = _T_42 | _T_43 | _T_44 | _T_45; // @[src/main/scala/util/package.scala 73:59]
  wire  line_1186_clock;
  wire  line_1186_reset;
  wire  line_1186_valid;
  reg  line_1186_valid_reg;
  wire [1:0] _ex_reg_mem_size_T_6 = {_T_142,_T_140}; // @[src/main/scala/rocket/RocketCore.scala 499:29]
  wire  do_bypass = id_bypass_src_0_0 | id_bypass_src_0_1 | id_bypass_src_0_2 | id_bypass_src_0_3; // @[src/main/scala/rocket/RocketCore.scala 511:48]
  wire [1:0] _bypass_src_T = id_bypass_src_0_2 ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _bypass_src_T_1 = id_bypass_src_0_1 ? 2'h1 : _bypass_src_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  _T_52 = id_ctrl_decoder_7 & ~do_bypass; // @[src/main/scala/rocket/RocketCore.scala 515:23]
  wire  line_1187_clock;
  wire  line_1187_reset;
  wire  line_1187_valid;
  reg  line_1187_valid_reg;
  wire  _wb_valid_T_2 = ~wb_xcpt; // @[src/main/scala/rocket/RocketCore.scala 739:48]
  wire  wb_valid = wb_reg_valid & ~replay_wb & ~wb_xcpt; // @[src/main/scala/rocket/RocketCore.scala 739:45]
  wire  wb_wen = wb_valid & wb_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 740:25]
  wire  rf_wen = wb_wen | ll_wen; // @[src/main/scala/rocket/RocketCore.scala 741:23]
  wire [4:0] rf_waddr = ll_wen ? ll_waddr : wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 742:21]
  wire  _T_135 = rf_waddr != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 1206:16]
  wire  _T_138 = rf_waddr == id_raddr1; // @[src/main/scala/rocket/RocketCore.scala 1209:20]
  wire [63:0] ll_wdata = div_io_resp_bits_data; // @[src/main/scala/rocket/RocketCore.scala 711:{29,29}]
  wire  _rf_wdata_T_4 = wb_ctrl_csr != 3'h0; // @[src/main/scala/rocket/RocketCore.scala 745:34]
  wire [63:0] _rf_wdata_T_6 = wb_ctrl_csr != 3'h0 ? csr_io_rw_rdata : wb_reg_wdata; // @[src/main/scala/rocket/RocketCore.scala 745:21]
  wire [63:0] _rf_wdata_T_7 = ll_wen ? ll_wdata : _rf_wdata_T_6; // @[src/main/scala/rocket/RocketCore.scala 744:21]
  wire [63:0] rf_wdata = dmem_resp_valid & dmem_resp_xpu & dmem_resp_waddr != 5'h0 ? io_dmem_resp_bits_data :
    _rf_wdata_T_7; // @[src/main/scala/rocket/RocketCore.scala 743:21]
  wire [63:0] _GEN_447 = rf_waddr == id_raddr1 ? rf_wdata : _GEN_153; // @[src/main/scala/rocket/RocketCore.scala 1201:19 1209:{31,39}]
  wire [63:0] _GEN_480 = rf_waddr != 5'h0 ? _GEN_447 : _GEN_153; // @[src/main/scala/rocket/RocketCore.scala 1201:19 1206:25]
  wire [63:0] id_rs_0 = rf_wen ? _GEN_480 : _GEN_153; // @[src/main/scala/rocket/RocketCore.scala 748:17 1201:19]
  wire  do_bypass_1 = id_bypass_src_1_0 | id_bypass_src_1_1 | id_bypass_src_1_2 | id_bypass_src_1_3; // @[src/main/scala/rocket/RocketCore.scala 511:48]
  wire [1:0] _bypass_src_T_2 = id_bypass_src_1_2 ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  _T_54 = id_ctrl_decoder_6 & ~do_bypass_1; // @[src/main/scala/rocket/RocketCore.scala 515:23]
  wire  line_1188_clock;
  wire  line_1188_reset;
  wire  line_1188_valid;
  reg  line_1188_valid_reg;
  wire  _T_139 = rf_waddr == id_raddr2; // @[src/main/scala/rocket/RocketCore.scala 1209:20]
  wire [63:0] _GEN_448 = rf_waddr == id_raddr2 ? rf_wdata : _GEN_184; // @[src/main/scala/rocket/RocketCore.scala 1201:19 1209:{31,39}]
  wire [63:0] _GEN_481 = rf_waddr != 5'h0 ? _GEN_448 : _GEN_184; // @[src/main/scala/rocket/RocketCore.scala 1201:19 1206:25]
  wire [63:0] id_rs_1 = rf_wen ? _GEN_481 : _GEN_184; // @[src/main/scala/rocket/RocketCore.scala 748:17 1201:19]
  wire  line_1189_clock;
  wire  line_1189_reset;
  wire  line_1189_valid;
  reg  line_1189_valid_reg;
  wire [31:0] inst = ibuf_io_inst_0_bits_rvc ? {{16'd0}, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw; // @[src/main/scala/rocket/RocketCore.scala 521:21]
  wire  id_load_use = mem_reg_valid & data_hazard_mem & mem_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 872:51]
  wire  _T_58 = _ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 527:41]
  wire  line_1190_clock;
  wire  line_1190_reset;
  wire  line_1190_valid;
  reg  line_1190_valid_reg;
  wire  ex_pc_valid = ex_reg_valid | ex_reg_replay | ex_reg_xcpt_interrupt; // @[src/main/scala/rocket/RocketCore.scala 537:51]
  wire  _replay_ex_structural_T = ~io_dmem_req_ready; // @[src/main/scala/rocket/RocketCore.scala 539:45]
  wire  _replay_ex_structural_T_3 = ex_ctrl_div & ~div_io_req_ready; // @[src/main/scala/rocket/RocketCore.scala 540:42]
  wire  replay_ex_structural = ex_ctrl_mem & ~io_dmem_req_ready | _replay_ex_structural_T_3; // @[src/main/scala/rocket/RocketCore.scala 539:64]
  wire  replay_ex_load_use = wb_dcache_miss & ex_reg_load_use; // @[src/main/scala/rocket/RocketCore.scala 541:43]
  wire  replay_ex = ex_reg_replay | ex_reg_valid & (replay_ex_structural | replay_ex_load_use); // @[src/main/scala/rocket/RocketCore.scala 542:33]
  wire  ctrl_killx = take_pc_mem_wb | replay_ex | ~ex_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 543:48]
  wire  ex_slow_bypass = ex_ctrl_mem_cmd == 5'h7 | ex_reg_mem_size < 2'h2; // @[src/main/scala/rocket/RocketCore.scala 545:50]
  wire  ex_sfence = ex_ctrl_mem & (ex_ctrl_mem_cmd == 5'h14 | ex_ctrl_mem_cmd == 5'h15 | ex_ctrl_mem_cmd == 5'h16); // @[src/main/scala/rocket/RocketCore.scala 546:44]
  wire  ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 549:28]
  wire  mem_pc_valid = mem_reg_valid | mem_reg_replay | mem_reg_xcpt_interrupt; // @[src/main/scala/rocket/RocketCore.scala 555:54]
  wire  mem_br_target_sign = mem_reg_inst[31]; // @[src/main/scala/rocket/RocketCore.scala 1217:49]
  wire [5:0] mem_br_target_b10_5 = mem_reg_inst[30:25]; // @[src/main/scala/rocket/RocketCore.scala 1223:62]
  wire [3:0] mem_br_target_b4_1 = mem_reg_inst[11:8]; // @[src/main/scala/rocket/RocketCore.scala 1225:57]
  wire  mem_br_target_hi_lo_lo = mem_reg_inst[7]; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [7:0] mem_br_target_hi_lo_hi = {8{mem_br_target_sign}}; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [10:0] mem_br_target_hi_hi_lo = {11{mem_br_target_sign}}; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire  mem_br_target_hi_hi_hi = mem_reg_inst[31]; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [31:0] _mem_br_target_T_3 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi,
    mem_br_target_hi_lo_lo,mem_br_target_b10_5,mem_br_target_b4_1,1'h0}; // @[src/main/scala/rocket/RocketCore.scala 1231:53]
  wire  mem_br_target_hi_lo_lo_1 = mem_reg_inst[20]; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [7:0] mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12]; // @[src/main/scala/rocket/RocketCore.scala 1231:8]
  wire [31:0] _mem_br_target_T_5 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi_1,
    mem_br_target_hi_lo_lo_1,mem_br_target_b10_5,mem_reg_inst[24:21],1'h0}; // @[src/main/scala/rocket/RocketCore.scala 1231:53]
  wire [3:0] _mem_br_target_T_6 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[src/main/scala/rocket/RocketCore.scala 559:8]
  wire [31:0] _mem_br_target_T_7 = mem_ctrl_jal ? $signed(_mem_br_target_T_5) : $signed({{28{_mem_br_target_T_6[3]}},
    _mem_br_target_T_6}); // @[src/main/scala/rocket/RocketCore.scala 558:8]
  wire [31:0] _mem_br_target_T_8 = _mem_cfi_taken_T ? $signed(_mem_br_target_T_3) : $signed(_mem_br_target_T_7); // @[src/main/scala/rocket/RocketCore.scala 557:8]
  wire [39:0] _GEN_519 = {{8{_mem_br_target_T_8[31]}},_mem_br_target_T_8}; // @[src/main/scala/rocket/RocketCore.scala 556:41]
  wire [39:0] mem_br_target = $signed(mem_reg_pc) + $signed(_GEN_519); // @[src/main/scala/rocket/RocketCore.scala 556:41]
  wire [24:0] mem_npc_a = mem_reg_wdata[63:39]; // @[src/main/scala/rocket/RocketCore.scala 1167:23]
  wire  mem_npc_msb = $signed(mem_npc_a) == 25'sh0 | $signed(mem_npc_a) == -25'sh1 ? mem_reg_wdata[39] : ~mem_reg_wdata[
    38]; // @[src/main/scala/rocket/RocketCore.scala 1168:18]
  wire [39:0] _mem_npc_T_3 = {mem_npc_msb,mem_reg_wdata[38:0]}; // @[src/main/scala/rocket/RocketCore.scala 560:106]
  wire [39:0] _mem_npc_T_4 = mem_ctrl_jalr | mem_reg_sfence ? $signed(_mem_npc_T_3) : $signed(mem_br_target); // @[src/main/scala/rocket/RocketCore.scala 560:21]
  wire [39:0] mem_npc = $signed(_mem_npc_T_4) & -40'sh2; // @[src/main/scala/rocket/RocketCore.scala 560:139]
  wire  _mem_wrong_npc_T_3 = ibuf_io_inst_0_valid | ibuf_io_imem_valid ? mem_npc != ibuf_io_pc : 1'h1; // @[src/main/scala/rocket/RocketCore.scala 563:8]
  wire  mem_wrong_npc = ex_pc_valid ? mem_npc != ex_reg_pc : _mem_wrong_npc_T_3; // @[src/main/scala/rocket/RocketCore.scala 562:8]
  wire  mem_npc_misaligned = _id_illegal_insn_T_18 & mem_npc[1] & ~mem_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 564:70]
  wire [63:0] mem_int_wdata = _take_pc_mem_T & (mem_ctrl_jalr ^ mem_npc_misaligned) ? $signed({{24{mem_br_target[39]}},
    mem_br_target}) : $signed(mem_reg_wdata); // @[src/main/scala/rocket/RocketCore.scala 565:119]
  wire  mem_cfi = mem_ctrl_branch | mem_ctrl_jalr | mem_ctrl_jal; // @[src/main/scala/rocket/RocketCore.scala 566:50]
  wire  _mem_reg_valid_T = ~ctrl_killx; // @[src/main/scala/rocket/RocketCore.scala 572:20]
  wire  _T_69 = mem_reg_valid & mem_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 579:23]
  wire  line_1191_clock;
  wire  line_1191_reset;
  wire  line_1191_valid;
  reg  line_1191_valid_reg;
  wire  line_1192_clock;
  wire  line_1192_reset;
  wire  line_1192_valid;
  reg  line_1192_valid_reg;
  wire  line_1193_clock;
  wire  line_1193_reset;
  wire  line_1193_valid;
  reg  line_1193_valid_reg;
  wire  _mem_reg_wdata_T_4 = ~ex_ctrl_zbk & ~ex_ctrl_zkn & ~ex_ctrl_zks; // @[src/main/scala/rocket/RocketCore.scala 603:37]
  wire  _T_72 = ex_ctrl_rxs2 & (ex_ctrl_mem | ex_ctrl_rocc | ex_sfence); // @[src/main/scala/rocket/RocketCore.scala 608:24]
  wire  line_1194_clock;
  wire  line_1194_reset;
  wire  line_1194_valid;
  reg  line_1194_valid_reg;
  wire [1:0] size = ex_ctrl_rocc ? 2'h3 : ex_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 609:21]
  wire [63:0] _mem_reg_rs2_T_4 = {ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[7:0],ex_rs_1[
    7:0],ex_rs_1[7:0]}; // @[src/main/scala/rocket/AMOALU.scala 28:32]
  wire [63:0] _mem_reg_rs2_T_8 = {ex_rs_1[15:0],ex_rs_1[15:0],ex_rs_1[15:0],ex_rs_1[15:0]}; // @[src/main/scala/rocket/AMOALU.scala 28:32]
  wire [63:0] _mem_reg_rs2_T_11 = {ex_rs_1[31:0],ex_rs_1[31:0]}; // @[src/main/scala/rocket/AMOALU.scala 28:32]
  wire [63:0] _mem_reg_rs2_T_12 = size == 2'h2 ? _mem_reg_rs2_T_11 : ex_rs_1; // @[src/main/scala/rocket/AMOALU.scala 28:13]
  wire [63:0] _mem_reg_rs2_T_13 = size == 2'h1 ? _mem_reg_rs2_T_8 : _mem_reg_rs2_T_12; // @[src/main/scala/rocket/AMOALU.scala 28:13]
  wire  _T_73 = ex_ctrl_jalr & csr_io_status_debug; // @[src/main/scala/rocket/RocketCore.scala 612:24]
  wire  line_1195_clock;
  wire  line_1195_reset;
  wire  line_1195_valid;
  reg  line_1195_valid_reg;
  wire  _GEN_263 = ex_ctrl_jalr & csr_io_status_debug | ex_ctrl_fence_i; // @[src/main/scala/rocket/RocketCore.scala 582:14 612:48 614:24]
  wire  _GEN_264 = ex_ctrl_jalr & csr_io_status_debug | ex_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 588:24 612:48 615:26]
  wire  _T_74 = mem_reg_xcpt_interrupt | mem_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 626:29]
  wire  _T_75 = mem_reg_valid & mem_npc_misaligned; // @[src/main/scala/rocket/RocketCore.scala 627:20]
  wire  mem_xcpt = _T_74 | _T_75; // @[src/main/scala/rocket/RocketCore.scala 1152:26]
  wire [3:0] _T_78 = _T_75 ? 4'h0 : 4'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  dcache_kill_mem = _T_30 & io_dmem_replay_next; // @[src/main/scala/rocket/RocketCore.scala 637:55]
  wire  replay_mem = dcache_kill_mem | mem_reg_replay; // @[src/main/scala/rocket/RocketCore.scala 639:37]
  wire  killm_common = dcache_kill_mem | take_pc_wb | mem_reg_xcpt | ~mem_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 640:68]
  reg  div_io_kill_REG; // @[src/main/scala/rocket/RocketCore.scala 641:41]
  wire  ctrl_killm = killm_common | mem_xcpt; // @[src/main/scala/rocket/RocketCore.scala 642:33]
  wire  _wb_reg_valid_T = ~ctrl_killm; // @[src/main/scala/rocket/RocketCore.scala 645:19]
  wire  _wb_reg_replay_T = ~take_pc_wb; // @[src/main/scala/rocket/RocketCore.scala 646:34]
  wire  line_1196_clock;
  wire  line_1196_reset;
  wire  line_1196_valid;
  reg  line_1196_valid_reg;
  wire  _T_91 = mem_ctrl_rocc | mem_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 653:25]
  wire  line_1197_clock;
  wire  line_1197_reset;
  wire  line_1197_valid;
  reg  line_1197_valid_reg;
  wire [2:0] _T_115 = _T_105 ? 3'h7 : 3'h5; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_116 = {{2'd0}, _T_115}; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_118 = _T_99 ? 5'hd : _T_116; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_119 = _T_97 ? 5'hf : _T_118; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_120 = _T_95 ? 5'h4 : _T_119; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _T_121 = _T_93 ? 5'h6 : _T_120; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  line_1198_clock;
  wire  line_1198_reset;
  wire  line_1198_valid;
  reg  line_1198_valid_reg;
  wire  ll_wen_try = div_io_resp_valid | _T_134; // @[src/main/scala/rocket/RocketCore.scala 737:60]
  wire  line_1199_clock;
  wire  line_1199_reset;
  wire  line_1199_valid;
  reg  line_1199_valid_reg;
  wire  line_1200_clock;
  wire  line_1200_reset;
  wire  line_1200_valid;
  reg  line_1200_valid_reg;
  wire [4:0] _T_137 = ~rf_waddr; // @[src/main/scala/rocket/RocketCore.scala 1195:39]
  wire  line_1201_clock;
  wire  line_1201_reset;
  wire  line_1201_valid;
  reg  line_1201_valid_reg;
  wire  line_1202_clock;
  wire  line_1202_reset;
  wire  line_1202_valid;
  reg  line_1202_valid_reg;
  wire  line_1203_clock;
  wire  line_1203_reset;
  wire  line_1203_valid;
  reg  line_1203_valid_reg;
  wire  line_1204_clock;
  wire  line_1204_reset;
  wire  line_1204_valid;
  reg  line_1204_valid_reg;
  wire  line_1205_clock;
  wire  line_1205_reset;
  wire  line_1205_valid;
  reg  line_1205_valid_reg;
  wire  line_1206_clock;
  wire  line_1206_reset;
  wire  line_1206_valid;
  reg  line_1206_valid_reg;
  wire  line_1207_clock;
  wire  line_1207_reset;
  wire  line_1207_valid;
  reg  line_1207_valid_reg;
  wire  line_1208_clock;
  wire  line_1208_reset;
  wire  line_1208_valid;
  reg  line_1208_valid_reg;
  wire  line_1209_clock;
  wire  line_1209_reset;
  wire  line_1209_valid;
  reg  line_1209_valid_reg;
  wire  line_1210_clock;
  wire  line_1210_reset;
  wire  line_1210_valid;
  reg  line_1210_valid_reg;
  wire  line_1211_clock;
  wire  line_1211_reset;
  wire  line_1211_valid;
  reg  line_1211_valid_reg;
  wire  line_1212_clock;
  wire  line_1212_reset;
  wire  line_1212_valid;
  reg  line_1212_valid_reg;
  wire  line_1213_clock;
  wire  line_1213_reset;
  wire  line_1213_valid;
  reg  line_1213_valid_reg;
  wire  line_1214_clock;
  wire  line_1214_reset;
  wire  line_1214_valid;
  reg  line_1214_valid_reg;
  wire  line_1215_clock;
  wire  line_1215_reset;
  wire  line_1215_valid;
  reg  line_1215_valid_reg;
  wire  line_1216_clock;
  wire  line_1216_reset;
  wire  line_1216_valid;
  reg  line_1216_valid_reg;
  wire  line_1217_clock;
  wire  line_1217_reset;
  wire  line_1217_valid;
  reg  line_1217_valid_reg;
  wire  line_1218_clock;
  wire  line_1218_reset;
  wire  line_1218_valid;
  reg  line_1218_valid_reg;
  wire  line_1219_clock;
  wire  line_1219_reset;
  wire  line_1219_valid;
  reg  line_1219_valid_reg;
  wire  line_1220_clock;
  wire  line_1220_reset;
  wire  line_1220_valid;
  reg  line_1220_valid_reg;
  wire  line_1221_clock;
  wire  line_1221_reset;
  wire  line_1221_valid;
  reg  line_1221_valid_reg;
  wire  line_1222_clock;
  wire  line_1222_reset;
  wire  line_1222_valid;
  reg  line_1222_valid_reg;
  wire  line_1223_clock;
  wire  line_1223_reset;
  wire  line_1223_valid;
  reg  line_1223_valid_reg;
  wire  line_1224_clock;
  wire  line_1224_reset;
  wire  line_1224_valid;
  reg  line_1224_valid_reg;
  wire  line_1225_clock;
  wire  line_1225_reset;
  wire  line_1225_valid;
  reg  line_1225_valid_reg;
  wire  line_1226_clock;
  wire  line_1226_reset;
  wire  line_1226_valid;
  reg  line_1226_valid_reg;
  wire  line_1227_clock;
  wire  line_1227_reset;
  wire  line_1227_valid;
  reg  line_1227_valid_reg;
  wire  line_1228_clock;
  wire  line_1228_reset;
  wire  line_1228_valid;
  reg  line_1228_valid_reg;
  wire  line_1229_clock;
  wire  line_1229_reset;
  wire  line_1229_valid;
  reg  line_1229_valid_reg;
  wire  line_1230_clock;
  wire  line_1230_reset;
  wire  line_1230_valid;
  reg  line_1230_valid_reg;
  wire  line_1231_clock;
  wire  line_1231_reset;
  wire  line_1231_valid;
  reg  line_1231_valid_reg;
  wire  line_1232_clock;
  wire  line_1232_reset;
  wire  line_1232_valid;
  reg  line_1232_valid_reg;
  wire  line_1233_clock;
  wire  line_1233_reset;
  wire  line_1233_valid;
  reg  line_1233_valid_reg;
  wire [15:0] _csr_io_inst_0_T_3 = &wb_reg_raw_inst[1:0] ? wb_reg_inst[31:16] : 16'h0; // @[src/main/scala/rocket/RocketCore.scala 768:50]
  wire  tval_dmem_addr = ~wb_reg_xcpt; // @[src/main/scala/rocket/RocketCore.scala 777:24]
  wire  _tval_any_addr_T = wb_reg_cause == 64'h3; // @[src/main/scala/util/package.scala 16:47]
  wire  _tval_any_addr_T_1 = wb_reg_cause == 64'h1; // @[src/main/scala/util/package.scala 16:47]
  wire  _tval_any_addr_T_2 = wb_reg_cause == 64'hc; // @[src/main/scala/util/package.scala 16:47]
  wire  _tval_any_addr_T_3 = wb_reg_cause == 64'h14; // @[src/main/scala/util/package.scala 16:47]
  wire  _tval_any_addr_T_6 = _tval_any_addr_T | _tval_any_addr_T_1 | _tval_any_addr_T_2 | _tval_any_addr_T_3; // @[src/main/scala/util/package.scala 73:59]
  wire  tval_any_addr = tval_dmem_addr | _tval_any_addr_T_6; // @[src/main/scala/rocket/RocketCore.scala 778:38]
  wire  tval_inst = wb_reg_cause == 64'h2; // @[src/main/scala/rocket/RocketCore.scala 780:32]
  wire  tval_valid = wb_xcpt & (tval_any_addr | tval_inst); // @[src/main/scala/rocket/RocketCore.scala 781:28]
  wire [24:0] csr_io_tval_a = wb_reg_wdata[63:39]; // @[src/main/scala/rocket/RocketCore.scala 1167:23]
  wire  csr_io_tval_msb = $signed(csr_io_tval_a) == 25'sh0 | $signed(csr_io_tval_a) == -25'sh1 ? wb_reg_wdata[39] : ~
    wb_reg_wdata[38]; // @[src/main/scala/rocket/RocketCore.scala 1168:18]
  wire [39:0] _csr_io_tval_T_1 = {csr_io_tval_msb,wb_reg_wdata[38:0]}; // @[src/main/scala/rocket/RocketCore.scala 1169:8]
  wire  csr_io_htval_htval_valid_imem = wb_reg_xcpt & _tval_any_addr_T_3; // @[src/main/scala/rocket/RocketCore.scala 785:40]
  wire  _csr_io_htval_T_3 = ~reset; // @[src/main/scala/rocket/RocketCore.scala 787:11]
  wire  line_1234_clock;
  wire  line_1234_reset;
  wire  line_1234_valid;
  reg  line_1234_valid_reg;
  wire  _csr_io_htval_T_4 = ~(~csr_io_htval_htval_valid_imem); // @[src/main/scala/rocket/RocketCore.scala 787:11]
  wire  line_1235_clock;
  wire  line_1235_reset;
  wire  line_1235_valid;
  reg  line_1235_valid_reg;
  wire [2:0] _csr_io_rw_cmd_T = wb_reg_valid ? 3'h0 : 3'h4; // @[src/main/scala/rocket/CSR.scala 185:15]
  wire [2:0] _csr_io_rw_cmd_T_1 = ~_csr_io_rw_cmd_T; // @[src/main/scala/rocket/CSR.scala 185:11]
  wire [31:0] _T_146 = 32'h1 << ll_waddr; // @[src/main/scala/rocket/RocketCore.scala 1183:58]
  wire [31:0] _T_147 = ll_wen ? _T_146 : 32'h0; // @[src/main/scala/rocket/RocketCore.scala 1183:49]
  wire [31:0] _T_148 = ~_T_147; // @[src/main/scala/rocket/RocketCore.scala 1175:64]
  wire [31:0] _T_149 = r & _T_148; // @[src/main/scala/rocket/RocketCore.scala 1175:62]
  wire  line_1236_clock;
  wire  line_1236_reset;
  wire  line_1236_valid;
  reg  line_1236_valid_reg;
  wire  _T_151 = wb_set_sboard & wb_wen; // @[src/main/scala/rocket/RocketCore.scala 856:28]
  wire [31:0] _T_152 = 32'h1 << wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 1183:58]
  wire [31:0] _T_153 = _T_151 ? _T_152 : 32'h0; // @[src/main/scala/rocket/RocketCore.scala 1183:49]
  wire [31:0] _T_154 = _T_149 | _T_153; // @[src/main/scala/rocket/RocketCore.scala 1174:60]
  wire  _T_155 = ll_wen | _T_151; // @[src/main/scala/rocket/RocketCore.scala 1186:17]
  wire  line_1237_clock;
  wire  line_1237_reset;
  wire  line_1237_valid;
  reg  line_1237_valid_reg;
  wire [39:0] _io_imem_req_bits_pc_T_1 = replay_wb ? wb_reg_pc : mem_npc; // @[src/main/scala/rocket/RocketCore.scala 916:8]
  wire  _io_imem_progress_T = ~replay_wb_common; // @[src/main/scala/rocket/RocketCore.scala 923:47]
  reg  io_imem_progress_REG; // @[src/main/scala/rocket/RocketCore.scala 923:30]
  wire [5:0] ex_dcache_tag = {ex_waddr,ex_ctrl_fp}; // @[src/main/scala/rocket/RocketCore.scala 970:26]
  wire [24:0] io_dmem_req_bits_addr_a = ex_rs_0[63:39]; // @[src/main/scala/rocket/RocketCore.scala 1167:23]
  wire  io_dmem_req_bits_addr_msb = $signed(io_dmem_req_bits_addr_a) == 25'sh0 | $signed(io_dmem_req_bits_addr_a) == -25'sh1
     ? alu_io_adder_out[39] : ~alu_io_adder_out[38]; // @[src/main/scala/rocket/RocketCore.scala 1168:18]
  wire  unpause = csr_io_time[4:0] == 5'h0 | io_dmem_perf_release | take_pc_mem_wb; // @[src/main/scala/rocket/RocketCore.scala 1002:118]
  wire  line_1238_clock;
  wire  line_1238_reset;
  wire  line_1238_valid;
  reg  line_1238_valid_reg;
  wire [39:0] _coreMonitorBundle_pc_T = csr_io_trace_0_iaddr; // @[src/main/scala/rocket/RocketCore.scala 1031:48]
  wire [23:0] _coreMonitorBundle_pc_T_2 = _coreMonitorBundle_pc_T[39] ? 24'hffffff : 24'h0; // @[src/main/scala/util/package.scala 124:20]
  wire  rf_delayed = _T_151 & wb_waddr != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 1103:46]
  wire [31:0] coreMonitorBundle_inst = csr_io_trace_0_insn; // @[src/main/scala/rocket/RocketCore.scala 1024:31 1040:26]
  wire  isWFI = coreMonitorBundle_inst == 32'h10500073; // @[src/main/scala/rocket/RocketCore.scala 1106:32]
  wire  _T_156 = rf_delayed | wb_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 1108:32]
  wire [1:0] _difftest_special_T = {isWFI,_T_156}; // @[difftest/src/main/scala/Bundles.scala 81:19]
  IBuf ibuf ( // @[src/main/scala/rocket/RocketCore.scala 284:20]
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_gf_inst(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw)
  );
  CSRFile csr ( // @[src/main/scala/rocket/RocketCore.scala 313:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_ungated_clock(csr_io_ungated_clock),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_0_inst(csr_io_decode_0_inst),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_rocc_illegal(csr_io_decode_0_rocc_illegal),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_rw_stall(csr_io_rw_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_cease(csr_io_status_cease),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_dv(csr_io_status_dv),
    .io_status_prv(csr_io_status_prv),
    .io_status_v(csr_io_status_v),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_mpv(csr_io_status_mpv),
    .io_status_gva(csr_io_status_gva),
    .io_status_mbe(csr_io_status_mbe),
    .io_status_sbe(csr_io_status_sbe),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_vs(csr_io_status_vs),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_ube(csr_io_status_ube),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_tval(csr_io_tval),
    .io_gva(csr_io_gva),
    .io_time(csr_io_time),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_csrr_counter(csr_io_csrr_counter),
    .io_inst_0(csr_io_inst_0),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_trace_0_interrupt(csr_io_trace_0_interrupt),
    .io_difftest_privilegeMode(csr_io_difftest_privilegeMode),
    .io_difftest_mstatus(csr_io_difftest_mstatus),
    .io_difftest_sstatus(csr_io_difftest_sstatus),
    .io_difftest_mepc(csr_io_difftest_mepc),
    .io_difftest_sepc(csr_io_difftest_sepc),
    .io_difftest_mtval(csr_io_difftest_mtval),
    .io_difftest_stval(csr_io_difftest_stval),
    .io_difftest_mtvec(csr_io_difftest_mtvec),
    .io_difftest_stvec(csr_io_difftest_stvec),
    .io_difftest_mcause(csr_io_difftest_mcause),
    .io_difftest_scause(csr_io_difftest_scause),
    .io_difftest_satp(csr_io_difftest_satp),
    .io_difftest_mip(csr_io_difftest_mip),
    .io_difftest_mie(csr_io_difftest_mie),
    .io_difftest_mscratch(csr_io_difftest_mscratch),
    .io_difftest_sscratch(csr_io_difftest_sscratch),
    .io_difftest_mideleg(csr_io_difftest_mideleg),
    .io_difftest_medeleg(csr_io_difftest_medeleg),
    .io_snapshot_minstret(csr_io_snapshot_minstret),
    .io_snapshot_mcycle(csr_io_snapshot_mcycle)
  );
  BreakpointUnit bpu ( // @[src/main/scala/rocket/RocketCore.scala 351:19]
    .clock(bpu_clock),
    .reset(bpu_reset)
  );
  ALU alu ( // @[src/main/scala/rocket/RocketCore.scala 416:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div ( // @[src/main/scala/rocket/RocketCore.scala 454:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  DummyDPICWrapper_4 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_value_1(difftest_module_io_bits_value_1),
    .io_bits_value_2(difftest_module_io_bits_value_2),
    .io_bits_value_3(difftest_module_io_bits_value_3),
    .io_bits_value_4(difftest_module_io_bits_value_4),
    .io_bits_value_5(difftest_module_io_bits_value_5),
    .io_bits_value_6(difftest_module_io_bits_value_6),
    .io_bits_value_7(difftest_module_io_bits_value_7),
    .io_bits_value_8(difftest_module_io_bits_value_8),
    .io_bits_value_9(difftest_module_io_bits_value_9),
    .io_bits_value_10(difftest_module_io_bits_value_10),
    .io_bits_value_11(difftest_module_io_bits_value_11),
    .io_bits_value_12(difftest_module_io_bits_value_12),
    .io_bits_value_13(difftest_module_io_bits_value_13),
    .io_bits_value_14(difftest_module_io_bits_value_14),
    .io_bits_value_15(difftest_module_io_bits_value_15),
    .io_bits_value_16(difftest_module_io_bits_value_16),
    .io_bits_value_17(difftest_module_io_bits_value_17),
    .io_bits_value_18(difftest_module_io_bits_value_18),
    .io_bits_value_19(difftest_module_io_bits_value_19),
    .io_bits_value_20(difftest_module_io_bits_value_20),
    .io_bits_value_21(difftest_module_io_bits_value_21),
    .io_bits_value_22(difftest_module_io_bits_value_22),
    .io_bits_value_23(difftest_module_io_bits_value_23),
    .io_bits_value_24(difftest_module_io_bits_value_24),
    .io_bits_value_25(difftest_module_io_bits_value_25),
    .io_bits_value_26(difftest_module_io_bits_value_26),
    .io_bits_value_27(difftest_module_io_bits_value_27),
    .io_bits_value_28(difftest_module_io_bits_value_28),
    .io_bits_value_29(difftest_module_io_bits_value_29),
    .io_bits_value_30(difftest_module_io_bits_value_30),
    .io_bits_value_31(difftest_module_io_bits_value_31)
  );
  DummyDPICWrapper_5 difftest_module_1 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_1_clock),
    .reset(difftest_module_1_reset),
    .io_valid(difftest_module_1_io_valid),
    .io_bits_valid(difftest_module_1_io_bits_valid),
    .io_bits_address(difftest_module_1_io_bits_address),
    .io_bits_data(difftest_module_1_io_bits_data)
  );
  DummyDPICWrapper_6 difftest_module_2 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_2_clock),
    .reset(difftest_module_2_reset),
    .io_bits_privilegeMode(difftest_module_2_io_bits_privilegeMode),
    .io_bits_mstatus(difftest_module_2_io_bits_mstatus),
    .io_bits_sstatus(difftest_module_2_io_bits_sstatus),
    .io_bits_mepc(difftest_module_2_io_bits_mepc),
    .io_bits_sepc(difftest_module_2_io_bits_sepc),
    .io_bits_mtval(difftest_module_2_io_bits_mtval),
    .io_bits_stval(difftest_module_2_io_bits_stval),
    .io_bits_mtvec(difftest_module_2_io_bits_mtvec),
    .io_bits_stvec(difftest_module_2_io_bits_stvec),
    .io_bits_mcause(difftest_module_2_io_bits_mcause),
    .io_bits_scause(difftest_module_2_io_bits_scause),
    .io_bits_satp(difftest_module_2_io_bits_satp),
    .io_bits_mip(difftest_module_2_io_bits_mip),
    .io_bits_mie(difftest_module_2_io_bits_mie),
    .io_bits_mscratch(difftest_module_2_io_bits_mscratch),
    .io_bits_sscratch(difftest_module_2_io_bits_sscratch),
    .io_bits_mideleg(difftest_module_2_io_bits_mideleg),
    .io_bits_medeleg(difftest_module_2_io_bits_medeleg)
  );
  DummyDPICWrapper_7 difftest_module_3 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_3_clock),
    .reset(difftest_module_3_reset),
    .io_bits_minstret(difftest_module_3_io_bits_minstret),
    .io_bits_mcycle(difftest_module_3_io_bits_mcycle)
  );
  DelayReg_3 difftest_delayer ( // @[difftest/src/main/scala/util/Delayer.scala 54:15]
    .clock(difftest_delayer_clock),
    .reset(difftest_delayer_reset),
    .i_valid(difftest_delayer_i_valid),
    .i_skip(difftest_delayer_i_skip),
    .i_rfwen(difftest_delayer_i_rfwen),
    .i_fpwen(difftest_delayer_i_fpwen),
    .i_wpdest(difftest_delayer_i_wpdest),
    .i_wdest(difftest_delayer_i_wdest),
    .i_pc(difftest_delayer_i_pc),
    .i_instr(difftest_delayer_i_instr),
    .i_special(difftest_delayer_i_special),
    .o_valid(difftest_delayer_o_valid),
    .o_skip(difftest_delayer_o_skip),
    .o_rfwen(difftest_delayer_o_rfwen),
    .o_fpwen(difftest_delayer_o_fpwen),
    .o_wpdest(difftest_delayer_o_wpdest),
    .o_wdest(difftest_delayer_o_wdest),
    .o_pc(difftest_delayer_o_pc),
    .o_instr(difftest_delayer_o_instr),
    .o_special(difftest_delayer_o_special)
  );
  DummyDPICWrapper_8 difftest_module_4 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_4_clock),
    .reset(difftest_module_4_reset),
    .io_valid(difftest_module_4_io_valid),
    .io_bits_valid(difftest_module_4_io_bits_valid),
    .io_bits_skip(difftest_module_4_io_bits_skip),
    .io_bits_rfwen(difftest_module_4_io_bits_rfwen),
    .io_bits_fpwen(difftest_module_4_io_bits_fpwen),
    .io_bits_wpdest(difftest_module_4_io_bits_wpdest),
    .io_bits_wdest(difftest_module_4_io_bits_wdest),
    .io_bits_pc(difftest_module_4_io_bits_pc),
    .io_bits_instr(difftest_module_4_io_bits_instr),
    .io_bits_special(difftest_module_4_io_bits_special)
  );
  DelayReg_4 difftest_delayer_1 ( // @[difftest/src/main/scala/util/Delayer.scala 54:15]
    .clock(difftest_delayer_1_clock),
    .reset(difftest_delayer_1_reset),
    .i_valid(difftest_delayer_1_i_valid),
    .i_address(difftest_delayer_1_i_address),
    .i_data(difftest_delayer_1_i_data),
    .i_nack(difftest_delayer_1_i_nack),
    .o_valid(difftest_delayer_1_o_valid),
    .o_address(difftest_delayer_1_o_address),
    .o_data(difftest_delayer_1_o_data),
    .o_nack(difftest_delayer_1_o_nack)
  );
  DummyDPICWrapper_9 difftest_module_5 ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_5_clock),
    .reset(difftest_module_5_reset),
    .io_valid(difftest_module_5_io_valid),
    .io_bits_valid(difftest_module_5_io_bits_valid),
    .io_bits_address(difftest_module_5_io_bits_address),
    .io_bits_data(difftest_module_5_io_bits_data),
    .io_bits_nack(difftest_module_5_io_bits_nack)
  );
  PlusArgTimeout PlusArgTimeout ( // @[src/main/scala/util/PlusArg.scala 89:11]
    .clock(PlusArgTimeout_clock),
    .reset(PlusArgTimeout_reset),
    .io_count(PlusArgTimeout_io_count)
  );
  GEN_w1_line #(.COVER_INDEX(1117)) line_1117 (
    .clock(line_1117_clock),
    .reset(line_1117_reset),
    .valid(line_1117_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1118)) line_1118 (
    .clock(line_1118_clock),
    .reset(line_1118_reset),
    .valid(line_1118_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1119)) line_1119 (
    .clock(line_1119_clock),
    .reset(line_1119_reset),
    .valid(line_1119_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1120)) line_1120 (
    .clock(line_1120_clock),
    .reset(line_1120_reset),
    .valid(line_1120_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1121)) line_1121 (
    .clock(line_1121_clock),
    .reset(line_1121_reset),
    .valid(line_1121_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1122)) line_1122 (
    .clock(line_1122_clock),
    .reset(line_1122_reset),
    .valid(line_1122_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1123)) line_1123 (
    .clock(line_1123_clock),
    .reset(line_1123_reset),
    .valid(line_1123_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1124)) line_1124 (
    .clock(line_1124_clock),
    .reset(line_1124_reset),
    .valid(line_1124_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1125)) line_1125 (
    .clock(line_1125_clock),
    .reset(line_1125_reset),
    .valid(line_1125_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1126)) line_1126 (
    .clock(line_1126_clock),
    .reset(line_1126_reset),
    .valid(line_1126_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1127)) line_1127 (
    .clock(line_1127_clock),
    .reset(line_1127_reset),
    .valid(line_1127_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1128)) line_1128 (
    .clock(line_1128_clock),
    .reset(line_1128_reset),
    .valid(line_1128_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1129)) line_1129 (
    .clock(line_1129_clock),
    .reset(line_1129_reset),
    .valid(line_1129_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1130)) line_1130 (
    .clock(line_1130_clock),
    .reset(line_1130_reset),
    .valid(line_1130_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1131)) line_1131 (
    .clock(line_1131_clock),
    .reset(line_1131_reset),
    .valid(line_1131_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1132)) line_1132 (
    .clock(line_1132_clock),
    .reset(line_1132_reset),
    .valid(line_1132_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1133)) line_1133 (
    .clock(line_1133_clock),
    .reset(line_1133_reset),
    .valid(line_1133_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1134)) line_1134 (
    .clock(line_1134_clock),
    .reset(line_1134_reset),
    .valid(line_1134_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1135)) line_1135 (
    .clock(line_1135_clock),
    .reset(line_1135_reset),
    .valid(line_1135_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1136)) line_1136 (
    .clock(line_1136_clock),
    .reset(line_1136_reset),
    .valid(line_1136_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1137)) line_1137 (
    .clock(line_1137_clock),
    .reset(line_1137_reset),
    .valid(line_1137_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1138)) line_1138 (
    .clock(line_1138_clock),
    .reset(line_1138_reset),
    .valid(line_1138_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1139)) line_1139 (
    .clock(line_1139_clock),
    .reset(line_1139_reset),
    .valid(line_1139_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1140)) line_1140 (
    .clock(line_1140_clock),
    .reset(line_1140_reset),
    .valid(line_1140_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1141)) line_1141 (
    .clock(line_1141_clock),
    .reset(line_1141_reset),
    .valid(line_1141_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1142)) line_1142 (
    .clock(line_1142_clock),
    .reset(line_1142_reset),
    .valid(line_1142_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1143)) line_1143 (
    .clock(line_1143_clock),
    .reset(line_1143_reset),
    .valid(line_1143_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1144)) line_1144 (
    .clock(line_1144_clock),
    .reset(line_1144_reset),
    .valid(line_1144_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1145)) line_1145 (
    .clock(line_1145_clock),
    .reset(line_1145_reset),
    .valid(line_1145_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1146)) line_1146 (
    .clock(line_1146_clock),
    .reset(line_1146_reset),
    .valid(line_1146_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1147)) line_1147 (
    .clock(line_1147_clock),
    .reset(line_1147_reset),
    .valid(line_1147_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1148)) line_1148 (
    .clock(line_1148_clock),
    .reset(line_1148_reset),
    .valid(line_1148_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1149)) line_1149 (
    .clock(line_1149_clock),
    .reset(line_1149_reset),
    .valid(line_1149_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1150)) line_1150 (
    .clock(line_1150_clock),
    .reset(line_1150_reset),
    .valid(line_1150_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1151)) line_1151 (
    .clock(line_1151_clock),
    .reset(line_1151_reset),
    .valid(line_1151_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1152)) line_1152 (
    .clock(line_1152_clock),
    .reset(line_1152_reset),
    .valid(line_1152_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1153)) line_1153 (
    .clock(line_1153_clock),
    .reset(line_1153_reset),
    .valid(line_1153_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1154)) line_1154 (
    .clock(line_1154_clock),
    .reset(line_1154_reset),
    .valid(line_1154_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1155)) line_1155 (
    .clock(line_1155_clock),
    .reset(line_1155_reset),
    .valid(line_1155_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1156)) line_1156 (
    .clock(line_1156_clock),
    .reset(line_1156_reset),
    .valid(line_1156_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1157)) line_1157 (
    .clock(line_1157_clock),
    .reset(line_1157_reset),
    .valid(line_1157_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1158)) line_1158 (
    .clock(line_1158_clock),
    .reset(line_1158_reset),
    .valid(line_1158_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1159)) line_1159 (
    .clock(line_1159_clock),
    .reset(line_1159_reset),
    .valid(line_1159_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1160)) line_1160 (
    .clock(line_1160_clock),
    .reset(line_1160_reset),
    .valid(line_1160_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1161)) line_1161 (
    .clock(line_1161_clock),
    .reset(line_1161_reset),
    .valid(line_1161_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1162)) line_1162 (
    .clock(line_1162_clock),
    .reset(line_1162_reset),
    .valid(line_1162_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1163)) line_1163 (
    .clock(line_1163_clock),
    .reset(line_1163_reset),
    .valid(line_1163_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1164)) line_1164 (
    .clock(line_1164_clock),
    .reset(line_1164_reset),
    .valid(line_1164_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1165)) line_1165 (
    .clock(line_1165_clock),
    .reset(line_1165_reset),
    .valid(line_1165_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1166)) line_1166 (
    .clock(line_1166_clock),
    .reset(line_1166_reset),
    .valid(line_1166_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1167)) line_1167 (
    .clock(line_1167_clock),
    .reset(line_1167_reset),
    .valid(line_1167_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1168)) line_1168 (
    .clock(line_1168_clock),
    .reset(line_1168_reset),
    .valid(line_1168_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1169)) line_1169 (
    .clock(line_1169_clock),
    .reset(line_1169_reset),
    .valid(line_1169_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1170)) line_1170 (
    .clock(line_1170_clock),
    .reset(line_1170_reset),
    .valid(line_1170_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1171)) line_1171 (
    .clock(line_1171_clock),
    .reset(line_1171_reset),
    .valid(line_1171_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1172)) line_1172 (
    .clock(line_1172_clock),
    .reset(line_1172_reset),
    .valid(line_1172_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1173)) line_1173 (
    .clock(line_1173_clock),
    .reset(line_1173_reset),
    .valid(line_1173_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1174)) line_1174 (
    .clock(line_1174_clock),
    .reset(line_1174_reset),
    .valid(line_1174_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1175)) line_1175 (
    .clock(line_1175_clock),
    .reset(line_1175_reset),
    .valid(line_1175_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1176)) line_1176 (
    .clock(line_1176_clock),
    .reset(line_1176_reset),
    .valid(line_1176_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1177)) line_1177 (
    .clock(line_1177_clock),
    .reset(line_1177_reset),
    .valid(line_1177_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1178)) line_1178 (
    .clock(line_1178_clock),
    .reset(line_1178_reset),
    .valid(line_1178_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1179)) line_1179 (
    .clock(line_1179_clock),
    .reset(line_1179_reset),
    .valid(line_1179_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1180)) line_1180 (
    .clock(line_1180_clock),
    .reset(line_1180_reset),
    .valid(line_1180_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1181)) line_1181 (
    .clock(line_1181_clock),
    .reset(line_1181_reset),
    .valid(line_1181_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1182)) line_1182 (
    .clock(line_1182_clock),
    .reset(line_1182_reset),
    .valid(line_1182_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1183)) line_1183 (
    .clock(line_1183_clock),
    .reset(line_1183_reset),
    .valid(line_1183_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1184)) line_1184 (
    .clock(line_1184_clock),
    .reset(line_1184_reset),
    .valid(line_1184_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1185)) line_1185 (
    .clock(line_1185_clock),
    .reset(line_1185_reset),
    .valid(line_1185_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1186)) line_1186 (
    .clock(line_1186_clock),
    .reset(line_1186_reset),
    .valid(line_1186_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1187)) line_1187 (
    .clock(line_1187_clock),
    .reset(line_1187_reset),
    .valid(line_1187_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1188)) line_1188 (
    .clock(line_1188_clock),
    .reset(line_1188_reset),
    .valid(line_1188_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1189)) line_1189 (
    .clock(line_1189_clock),
    .reset(line_1189_reset),
    .valid(line_1189_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1190)) line_1190 (
    .clock(line_1190_clock),
    .reset(line_1190_reset),
    .valid(line_1190_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1191)) line_1191 (
    .clock(line_1191_clock),
    .reset(line_1191_reset),
    .valid(line_1191_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1192)) line_1192 (
    .clock(line_1192_clock),
    .reset(line_1192_reset),
    .valid(line_1192_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1193)) line_1193 (
    .clock(line_1193_clock),
    .reset(line_1193_reset),
    .valid(line_1193_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1194)) line_1194 (
    .clock(line_1194_clock),
    .reset(line_1194_reset),
    .valid(line_1194_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1195)) line_1195 (
    .clock(line_1195_clock),
    .reset(line_1195_reset),
    .valid(line_1195_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1196)) line_1196 (
    .clock(line_1196_clock),
    .reset(line_1196_reset),
    .valid(line_1196_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1197)) line_1197 (
    .clock(line_1197_clock),
    .reset(line_1197_reset),
    .valid(line_1197_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1198)) line_1198 (
    .clock(line_1198_clock),
    .reset(line_1198_reset),
    .valid(line_1198_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1199)) line_1199 (
    .clock(line_1199_clock),
    .reset(line_1199_reset),
    .valid(line_1199_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1200)) line_1200 (
    .clock(line_1200_clock),
    .reset(line_1200_reset),
    .valid(line_1200_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1201)) line_1201 (
    .clock(line_1201_clock),
    .reset(line_1201_reset),
    .valid(line_1201_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1202)) line_1202 (
    .clock(line_1202_clock),
    .reset(line_1202_reset),
    .valid(line_1202_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1203)) line_1203 (
    .clock(line_1203_clock),
    .reset(line_1203_reset),
    .valid(line_1203_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1204)) line_1204 (
    .clock(line_1204_clock),
    .reset(line_1204_reset),
    .valid(line_1204_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1205)) line_1205 (
    .clock(line_1205_clock),
    .reset(line_1205_reset),
    .valid(line_1205_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1206)) line_1206 (
    .clock(line_1206_clock),
    .reset(line_1206_reset),
    .valid(line_1206_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1207)) line_1207 (
    .clock(line_1207_clock),
    .reset(line_1207_reset),
    .valid(line_1207_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1208)) line_1208 (
    .clock(line_1208_clock),
    .reset(line_1208_reset),
    .valid(line_1208_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1209)) line_1209 (
    .clock(line_1209_clock),
    .reset(line_1209_reset),
    .valid(line_1209_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1210)) line_1210 (
    .clock(line_1210_clock),
    .reset(line_1210_reset),
    .valid(line_1210_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1211)) line_1211 (
    .clock(line_1211_clock),
    .reset(line_1211_reset),
    .valid(line_1211_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1212)) line_1212 (
    .clock(line_1212_clock),
    .reset(line_1212_reset),
    .valid(line_1212_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1213)) line_1213 (
    .clock(line_1213_clock),
    .reset(line_1213_reset),
    .valid(line_1213_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1214)) line_1214 (
    .clock(line_1214_clock),
    .reset(line_1214_reset),
    .valid(line_1214_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1215)) line_1215 (
    .clock(line_1215_clock),
    .reset(line_1215_reset),
    .valid(line_1215_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1216)) line_1216 (
    .clock(line_1216_clock),
    .reset(line_1216_reset),
    .valid(line_1216_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1217)) line_1217 (
    .clock(line_1217_clock),
    .reset(line_1217_reset),
    .valid(line_1217_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1218)) line_1218 (
    .clock(line_1218_clock),
    .reset(line_1218_reset),
    .valid(line_1218_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1219)) line_1219 (
    .clock(line_1219_clock),
    .reset(line_1219_reset),
    .valid(line_1219_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1220)) line_1220 (
    .clock(line_1220_clock),
    .reset(line_1220_reset),
    .valid(line_1220_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1221)) line_1221 (
    .clock(line_1221_clock),
    .reset(line_1221_reset),
    .valid(line_1221_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1222)) line_1222 (
    .clock(line_1222_clock),
    .reset(line_1222_reset),
    .valid(line_1222_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1223)) line_1223 (
    .clock(line_1223_clock),
    .reset(line_1223_reset),
    .valid(line_1223_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1224)) line_1224 (
    .clock(line_1224_clock),
    .reset(line_1224_reset),
    .valid(line_1224_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1225)) line_1225 (
    .clock(line_1225_clock),
    .reset(line_1225_reset),
    .valid(line_1225_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1226)) line_1226 (
    .clock(line_1226_clock),
    .reset(line_1226_reset),
    .valid(line_1226_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1227)) line_1227 (
    .clock(line_1227_clock),
    .reset(line_1227_reset),
    .valid(line_1227_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1228)) line_1228 (
    .clock(line_1228_clock),
    .reset(line_1228_reset),
    .valid(line_1228_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1229)) line_1229 (
    .clock(line_1229_clock),
    .reset(line_1229_reset),
    .valid(line_1229_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1230)) line_1230 (
    .clock(line_1230_clock),
    .reset(line_1230_reset),
    .valid(line_1230_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1231)) line_1231 (
    .clock(line_1231_clock),
    .reset(line_1231_reset),
    .valid(line_1231_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1232)) line_1232 (
    .clock(line_1232_clock),
    .reset(line_1232_reset),
    .valid(line_1232_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1233)) line_1233 (
    .clock(line_1233_clock),
    .reset(line_1233_reset),
    .valid(line_1233_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1234)) line_1234 (
    .clock(line_1234_clock),
    .reset(line_1234_reset),
    .valid(line_1234_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1235)) line_1235 (
    .clock(line_1235_clock),
    .reset(line_1235_reset),
    .valid(line_1235_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1236)) line_1236 (
    .clock(line_1236_clock),
    .reset(line_1236_reset),
    .valid(line_1236_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1237)) line_1237 (
    .clock(line_1237_clock),
    .reset(line_1237_reset),
    .valid(line_1237_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1238)) line_1238 (
    .clock(line_1238_clock),
    .reset(line_1238_reset),
    .valid(line_1238_valid)
  );
  assign line_1117_clock = clock;
  assign line_1117_reset = reset;
  assign line_1117_valid = 5'h0 == _id_rs_T_3 ^ line_1117_valid_reg;
  assign line_1118_clock = clock;
  assign line_1118_reset = reset;
  assign line_1118_valid = 5'h1 == _id_rs_T_3 ^ line_1118_valid_reg;
  assign line_1119_clock = clock;
  assign line_1119_reset = reset;
  assign line_1119_valid = 5'h2 == _id_rs_T_3 ^ line_1119_valid_reg;
  assign line_1120_clock = clock;
  assign line_1120_reset = reset;
  assign line_1120_valid = 5'h3 == _id_rs_T_3 ^ line_1120_valid_reg;
  assign line_1121_clock = clock;
  assign line_1121_reset = reset;
  assign line_1121_valid = 5'h4 == _id_rs_T_3 ^ line_1121_valid_reg;
  assign line_1122_clock = clock;
  assign line_1122_reset = reset;
  assign line_1122_valid = 5'h5 == _id_rs_T_3 ^ line_1122_valid_reg;
  assign line_1123_clock = clock;
  assign line_1123_reset = reset;
  assign line_1123_valid = 5'h6 == _id_rs_T_3 ^ line_1123_valid_reg;
  assign line_1124_clock = clock;
  assign line_1124_reset = reset;
  assign line_1124_valid = 5'h7 == _id_rs_T_3 ^ line_1124_valid_reg;
  assign line_1125_clock = clock;
  assign line_1125_reset = reset;
  assign line_1125_valid = 5'h8 == _id_rs_T_3 ^ line_1125_valid_reg;
  assign line_1126_clock = clock;
  assign line_1126_reset = reset;
  assign line_1126_valid = 5'h9 == _id_rs_T_3 ^ line_1126_valid_reg;
  assign line_1127_clock = clock;
  assign line_1127_reset = reset;
  assign line_1127_valid = 5'ha == _id_rs_T_3 ^ line_1127_valid_reg;
  assign line_1128_clock = clock;
  assign line_1128_reset = reset;
  assign line_1128_valid = 5'hb == _id_rs_T_3 ^ line_1128_valid_reg;
  assign line_1129_clock = clock;
  assign line_1129_reset = reset;
  assign line_1129_valid = 5'hc == _id_rs_T_3 ^ line_1129_valid_reg;
  assign line_1130_clock = clock;
  assign line_1130_reset = reset;
  assign line_1130_valid = 5'hd == _id_rs_T_3 ^ line_1130_valid_reg;
  assign line_1131_clock = clock;
  assign line_1131_reset = reset;
  assign line_1131_valid = 5'he == _id_rs_T_3 ^ line_1131_valid_reg;
  assign line_1132_clock = clock;
  assign line_1132_reset = reset;
  assign line_1132_valid = 5'hf == _id_rs_T_3 ^ line_1132_valid_reg;
  assign line_1133_clock = clock;
  assign line_1133_reset = reset;
  assign line_1133_valid = 5'h10 == _id_rs_T_3 ^ line_1133_valid_reg;
  assign line_1134_clock = clock;
  assign line_1134_reset = reset;
  assign line_1134_valid = 5'h11 == _id_rs_T_3 ^ line_1134_valid_reg;
  assign line_1135_clock = clock;
  assign line_1135_reset = reset;
  assign line_1135_valid = 5'h12 == _id_rs_T_3 ^ line_1135_valid_reg;
  assign line_1136_clock = clock;
  assign line_1136_reset = reset;
  assign line_1136_valid = 5'h13 == _id_rs_T_3 ^ line_1136_valid_reg;
  assign line_1137_clock = clock;
  assign line_1137_reset = reset;
  assign line_1137_valid = 5'h14 == _id_rs_T_3 ^ line_1137_valid_reg;
  assign line_1138_clock = clock;
  assign line_1138_reset = reset;
  assign line_1138_valid = 5'h15 == _id_rs_T_3 ^ line_1138_valid_reg;
  assign line_1139_clock = clock;
  assign line_1139_reset = reset;
  assign line_1139_valid = 5'h16 == _id_rs_T_3 ^ line_1139_valid_reg;
  assign line_1140_clock = clock;
  assign line_1140_reset = reset;
  assign line_1140_valid = 5'h17 == _id_rs_T_3 ^ line_1140_valid_reg;
  assign line_1141_clock = clock;
  assign line_1141_reset = reset;
  assign line_1141_valid = 5'h18 == _id_rs_T_3 ^ line_1141_valid_reg;
  assign line_1142_clock = clock;
  assign line_1142_reset = reset;
  assign line_1142_valid = 5'h19 == _id_rs_T_3 ^ line_1142_valid_reg;
  assign line_1143_clock = clock;
  assign line_1143_reset = reset;
  assign line_1143_valid = 5'h1a == _id_rs_T_3 ^ line_1143_valid_reg;
  assign line_1144_clock = clock;
  assign line_1144_reset = reset;
  assign line_1144_valid = 5'h1b == _id_rs_T_3 ^ line_1144_valid_reg;
  assign line_1145_clock = clock;
  assign line_1145_reset = reset;
  assign line_1145_valid = 5'h1c == _id_rs_T_3 ^ line_1145_valid_reg;
  assign line_1146_clock = clock;
  assign line_1146_reset = reset;
  assign line_1146_valid = 5'h1d == _id_rs_T_3 ^ line_1146_valid_reg;
  assign line_1147_clock = clock;
  assign line_1147_reset = reset;
  assign line_1147_valid = 5'h1e == _id_rs_T_3 ^ line_1147_valid_reg;
  assign line_1148_clock = clock;
  assign line_1148_reset = reset;
  assign line_1148_valid = 5'h0 == _id_rs_T_8 ^ line_1148_valid_reg;
  assign line_1149_clock = clock;
  assign line_1149_reset = reset;
  assign line_1149_valid = 5'h1 == _id_rs_T_8 ^ line_1149_valid_reg;
  assign line_1150_clock = clock;
  assign line_1150_reset = reset;
  assign line_1150_valid = 5'h2 == _id_rs_T_8 ^ line_1150_valid_reg;
  assign line_1151_clock = clock;
  assign line_1151_reset = reset;
  assign line_1151_valid = 5'h3 == _id_rs_T_8 ^ line_1151_valid_reg;
  assign line_1152_clock = clock;
  assign line_1152_reset = reset;
  assign line_1152_valid = 5'h4 == _id_rs_T_8 ^ line_1152_valid_reg;
  assign line_1153_clock = clock;
  assign line_1153_reset = reset;
  assign line_1153_valid = 5'h5 == _id_rs_T_8 ^ line_1153_valid_reg;
  assign line_1154_clock = clock;
  assign line_1154_reset = reset;
  assign line_1154_valid = 5'h6 == _id_rs_T_8 ^ line_1154_valid_reg;
  assign line_1155_clock = clock;
  assign line_1155_reset = reset;
  assign line_1155_valid = 5'h7 == _id_rs_T_8 ^ line_1155_valid_reg;
  assign line_1156_clock = clock;
  assign line_1156_reset = reset;
  assign line_1156_valid = 5'h8 == _id_rs_T_8 ^ line_1156_valid_reg;
  assign line_1157_clock = clock;
  assign line_1157_reset = reset;
  assign line_1157_valid = 5'h9 == _id_rs_T_8 ^ line_1157_valid_reg;
  assign line_1158_clock = clock;
  assign line_1158_reset = reset;
  assign line_1158_valid = 5'ha == _id_rs_T_8 ^ line_1158_valid_reg;
  assign line_1159_clock = clock;
  assign line_1159_reset = reset;
  assign line_1159_valid = 5'hb == _id_rs_T_8 ^ line_1159_valid_reg;
  assign line_1160_clock = clock;
  assign line_1160_reset = reset;
  assign line_1160_valid = 5'hc == _id_rs_T_8 ^ line_1160_valid_reg;
  assign line_1161_clock = clock;
  assign line_1161_reset = reset;
  assign line_1161_valid = 5'hd == _id_rs_T_8 ^ line_1161_valid_reg;
  assign line_1162_clock = clock;
  assign line_1162_reset = reset;
  assign line_1162_valid = 5'he == _id_rs_T_8 ^ line_1162_valid_reg;
  assign line_1163_clock = clock;
  assign line_1163_reset = reset;
  assign line_1163_valid = 5'hf == _id_rs_T_8 ^ line_1163_valid_reg;
  assign line_1164_clock = clock;
  assign line_1164_reset = reset;
  assign line_1164_valid = 5'h10 == _id_rs_T_8 ^ line_1164_valid_reg;
  assign line_1165_clock = clock;
  assign line_1165_reset = reset;
  assign line_1165_valid = 5'h11 == _id_rs_T_8 ^ line_1165_valid_reg;
  assign line_1166_clock = clock;
  assign line_1166_reset = reset;
  assign line_1166_valid = 5'h12 == _id_rs_T_8 ^ line_1166_valid_reg;
  assign line_1167_clock = clock;
  assign line_1167_reset = reset;
  assign line_1167_valid = 5'h13 == _id_rs_T_8 ^ line_1167_valid_reg;
  assign line_1168_clock = clock;
  assign line_1168_reset = reset;
  assign line_1168_valid = 5'h14 == _id_rs_T_8 ^ line_1168_valid_reg;
  assign line_1169_clock = clock;
  assign line_1169_reset = reset;
  assign line_1169_valid = 5'h15 == _id_rs_T_8 ^ line_1169_valid_reg;
  assign line_1170_clock = clock;
  assign line_1170_reset = reset;
  assign line_1170_valid = 5'h16 == _id_rs_T_8 ^ line_1170_valid_reg;
  assign line_1171_clock = clock;
  assign line_1171_reset = reset;
  assign line_1171_valid = 5'h17 == _id_rs_T_8 ^ line_1171_valid_reg;
  assign line_1172_clock = clock;
  assign line_1172_reset = reset;
  assign line_1172_valid = 5'h18 == _id_rs_T_8 ^ line_1172_valid_reg;
  assign line_1173_clock = clock;
  assign line_1173_reset = reset;
  assign line_1173_valid = 5'h19 == _id_rs_T_8 ^ line_1173_valid_reg;
  assign line_1174_clock = clock;
  assign line_1174_reset = reset;
  assign line_1174_valid = 5'h1a == _id_rs_T_8 ^ line_1174_valid_reg;
  assign line_1175_clock = clock;
  assign line_1175_reset = reset;
  assign line_1175_valid = 5'h1b == _id_rs_T_8 ^ line_1175_valid_reg;
  assign line_1176_clock = clock;
  assign line_1176_reset = reset;
  assign line_1176_valid = 5'h1c == _id_rs_T_8 ^ line_1176_valid_reg;
  assign line_1177_clock = clock;
  assign line_1177_reset = reset;
  assign line_1177_valid = 5'h1d == _id_rs_T_8 ^ line_1177_valid_reg;
  assign line_1178_clock = clock;
  assign line_1178_reset = reset;
  assign line_1178_valid = 5'h1e == _id_rs_T_8 ^ line_1178_valid_reg;
  assign line_1179_clock = clock;
  assign line_1179_reset = reset;
  assign line_1179_valid = _T ^ line_1179_valid_reg;
  assign line_1180_clock = clock;
  assign line_1180_reset = reset;
  assign line_1180_valid = _ex_reg_valid_T ^ line_1180_valid_reg;
  assign line_1181_clock = clock;
  assign line_1181_reset = reset;
  assign line_1181_valid = _T_36 ^ line_1181_valid_reg;
  assign line_1182_clock = clock;
  assign line_1182_reset = reset;
  assign line_1182_valid = id_fence_next ^ line_1182_valid_reg;
  assign line_1183_clock = clock;
  assign line_1183_reset = reset;
  assign line_1183_valid = id_xcpt ^ line_1183_valid_reg;
  assign line_1184_clock = clock;
  assign line_1184_reset = reset;
  assign line_1184_valid = _T_38 ^ line_1184_valid_reg;
  assign line_1185_clock = clock;
  assign line_1185_reset = reset;
  assign line_1185_valid = _T_40 ^ line_1185_valid_reg;
  assign line_1186_clock = clock;
  assign line_1186_reset = reset;
  assign line_1186_valid = _T_48 ^ line_1186_valid_reg;
  assign line_1187_clock = clock;
  assign line_1187_reset = reset;
  assign line_1187_valid = _T_52 ^ line_1187_valid_reg;
  assign line_1188_clock = clock;
  assign line_1188_reset = reset;
  assign line_1188_valid = _T_54 ^ line_1188_valid_reg;
  assign line_1189_clock = clock;
  assign line_1189_reset = reset;
  assign line_1189_valid = id_illegal_insn ^ line_1189_valid_reg;
  assign line_1190_clock = clock;
  assign line_1190_reset = reset;
  assign line_1190_valid = _T_58 ^ line_1190_valid_reg;
  assign line_1191_clock = clock;
  assign line_1191_reset = reset;
  assign line_1191_valid = _T_69 ^ line_1191_valid_reg;
  assign line_1192_clock = clock;
  assign line_1192_reset = reset;
  assign line_1192_valid = _T_69 ^ line_1192_valid_reg;
  assign line_1193_clock = clock;
  assign line_1193_reset = reset;
  assign line_1193_valid = ex_pc_valid ^ line_1193_valid_reg;
  assign line_1194_clock = clock;
  assign line_1194_reset = reset;
  assign line_1194_valid = _T_72 ^ line_1194_valid_reg;
  assign line_1195_clock = clock;
  assign line_1195_reset = reset;
  assign line_1195_valid = _T_73 ^ line_1195_valid_reg;
  assign line_1196_clock = clock;
  assign line_1196_reset = reset;
  assign line_1196_valid = mem_pc_valid ^ line_1196_valid_reg;
  assign line_1197_clock = clock;
  assign line_1197_reset = reset;
  assign line_1197_valid = _T_91 ^ line_1197_valid_reg;
  assign line_1198_clock = clock;
  assign line_1198_reset = reset;
  assign line_1198_valid = _T_134 ^ line_1198_valid_reg;
  assign line_1199_clock = clock;
  assign line_1199_reset = reset;
  assign line_1199_valid = rf_wen ^ line_1199_valid_reg;
  assign line_1200_clock = clock;
  assign line_1200_reset = reset;
  assign line_1200_valid = _T_135 ^ line_1200_valid_reg;
  assign line_1201_clock = clock;
  assign line_1201_reset = reset;
  assign line_1201_valid = 5'h0 == _T_137 ^ line_1201_valid_reg;
  assign line_1202_clock = clock;
  assign line_1202_reset = reset;
  assign line_1202_valid = 5'h1 == _T_137 ^ line_1202_valid_reg;
  assign line_1203_clock = clock;
  assign line_1203_reset = reset;
  assign line_1203_valid = 5'h2 == _T_137 ^ line_1203_valid_reg;
  assign line_1204_clock = clock;
  assign line_1204_reset = reset;
  assign line_1204_valid = 5'h3 == _T_137 ^ line_1204_valid_reg;
  assign line_1205_clock = clock;
  assign line_1205_reset = reset;
  assign line_1205_valid = 5'h4 == _T_137 ^ line_1205_valid_reg;
  assign line_1206_clock = clock;
  assign line_1206_reset = reset;
  assign line_1206_valid = 5'h5 == _T_137 ^ line_1206_valid_reg;
  assign line_1207_clock = clock;
  assign line_1207_reset = reset;
  assign line_1207_valid = 5'h6 == _T_137 ^ line_1207_valid_reg;
  assign line_1208_clock = clock;
  assign line_1208_reset = reset;
  assign line_1208_valid = 5'h7 == _T_137 ^ line_1208_valid_reg;
  assign line_1209_clock = clock;
  assign line_1209_reset = reset;
  assign line_1209_valid = 5'h8 == _T_137 ^ line_1209_valid_reg;
  assign line_1210_clock = clock;
  assign line_1210_reset = reset;
  assign line_1210_valid = 5'h9 == _T_137 ^ line_1210_valid_reg;
  assign line_1211_clock = clock;
  assign line_1211_reset = reset;
  assign line_1211_valid = 5'ha == _T_137 ^ line_1211_valid_reg;
  assign line_1212_clock = clock;
  assign line_1212_reset = reset;
  assign line_1212_valid = 5'hb == _T_137 ^ line_1212_valid_reg;
  assign line_1213_clock = clock;
  assign line_1213_reset = reset;
  assign line_1213_valid = 5'hc == _T_137 ^ line_1213_valid_reg;
  assign line_1214_clock = clock;
  assign line_1214_reset = reset;
  assign line_1214_valid = 5'hd == _T_137 ^ line_1214_valid_reg;
  assign line_1215_clock = clock;
  assign line_1215_reset = reset;
  assign line_1215_valid = 5'he == _T_137 ^ line_1215_valid_reg;
  assign line_1216_clock = clock;
  assign line_1216_reset = reset;
  assign line_1216_valid = 5'hf == _T_137 ^ line_1216_valid_reg;
  assign line_1217_clock = clock;
  assign line_1217_reset = reset;
  assign line_1217_valid = 5'h10 == _T_137 ^ line_1217_valid_reg;
  assign line_1218_clock = clock;
  assign line_1218_reset = reset;
  assign line_1218_valid = 5'h11 == _T_137 ^ line_1218_valid_reg;
  assign line_1219_clock = clock;
  assign line_1219_reset = reset;
  assign line_1219_valid = 5'h12 == _T_137 ^ line_1219_valid_reg;
  assign line_1220_clock = clock;
  assign line_1220_reset = reset;
  assign line_1220_valid = 5'h13 == _T_137 ^ line_1220_valid_reg;
  assign line_1221_clock = clock;
  assign line_1221_reset = reset;
  assign line_1221_valid = 5'h14 == _T_137 ^ line_1221_valid_reg;
  assign line_1222_clock = clock;
  assign line_1222_reset = reset;
  assign line_1222_valid = 5'h15 == _T_137 ^ line_1222_valid_reg;
  assign line_1223_clock = clock;
  assign line_1223_reset = reset;
  assign line_1223_valid = 5'h16 == _T_137 ^ line_1223_valid_reg;
  assign line_1224_clock = clock;
  assign line_1224_reset = reset;
  assign line_1224_valid = 5'h17 == _T_137 ^ line_1224_valid_reg;
  assign line_1225_clock = clock;
  assign line_1225_reset = reset;
  assign line_1225_valid = 5'h18 == _T_137 ^ line_1225_valid_reg;
  assign line_1226_clock = clock;
  assign line_1226_reset = reset;
  assign line_1226_valid = 5'h19 == _T_137 ^ line_1226_valid_reg;
  assign line_1227_clock = clock;
  assign line_1227_reset = reset;
  assign line_1227_valid = 5'h1a == _T_137 ^ line_1227_valid_reg;
  assign line_1228_clock = clock;
  assign line_1228_reset = reset;
  assign line_1228_valid = 5'h1b == _T_137 ^ line_1228_valid_reg;
  assign line_1229_clock = clock;
  assign line_1229_reset = reset;
  assign line_1229_valid = 5'h1c == _T_137 ^ line_1229_valid_reg;
  assign line_1230_clock = clock;
  assign line_1230_reset = reset;
  assign line_1230_valid = 5'h1d == _T_137 ^ line_1230_valid_reg;
  assign line_1231_clock = clock;
  assign line_1231_reset = reset;
  assign line_1231_valid = 5'h1e == _T_137 ^ line_1231_valid_reg;
  assign line_1232_clock = clock;
  assign line_1232_reset = reset;
  assign line_1232_valid = _T_138 ^ line_1232_valid_reg;
  assign line_1233_clock = clock;
  assign line_1233_reset = reset;
  assign line_1233_valid = _T_139 ^ line_1233_valid_reg;
  assign line_1234_clock = clock;
  assign line_1234_reset = reset;
  assign line_1234_valid = _csr_io_htval_T_3 ^ line_1234_valid_reg;
  assign line_1235_clock = clock;
  assign line_1235_reset = reset;
  assign line_1235_valid = _csr_io_htval_T_4 ^ line_1235_valid_reg;
  assign line_1236_clock = clock;
  assign line_1236_reset = reset;
  assign line_1236_valid = ll_wen ^ line_1236_valid_reg;
  assign line_1237_clock = clock;
  assign line_1237_reset = reset;
  assign line_1237_valid = _T_155 ^ line_1237_valid_reg;
  assign line_1238_clock = clock;
  assign line_1238_reset = reset;
  assign line_1238_valid = unpause ^ line_1238_valid_reg;
  assign io_imem_might_request = imem_might_request_reg; // @[src/main/scala/rocket/RocketCore.scala 919:25]
  assign io_imem_req_valid = take_pc_wb | take_pc_mem; // @[src/main/scala/rocket/RocketCore.scala 280:35]
  assign io_imem_req_bits_pc = wb_xcpt | csr_io_eret ? csr_io_evec : _io_imem_req_bits_pc_T_1; // @[src/main/scala/rocket/RocketCore.scala 915:8]
  assign io_imem_req_bits_speculative = ~take_pc_wb; // @[src/main/scala/rocket/RocketCore.scala 913:35]
  assign io_imem_sfence_valid = wb_reg_valid & wb_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 924:40]
  assign io_imem_sfence_bits_rs1 = wb_reg_mem_size[0]; // @[src/main/scala/rocket/RocketCore.scala 925:45]
  assign io_imem_sfence_bits_rs2 = wb_reg_mem_size[1]; // @[src/main/scala/rocket/RocketCore.scala 926:45]
  assign io_imem_sfence_bits_addr = wb_reg_wdata[38:0]; // @[src/main/scala/rocket/RocketCore.scala 927:28]
  assign io_imem_resp_ready = ibuf_io_imem_ready; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign io_imem_btb_update_valid = mem_reg_valid & _wb_reg_replay_T & mem_wrong_npc & (~mem_cfi | mem_cfi_taken); // @[src/main/scala/rocket/RocketCore.scala 935:77]
  assign io_imem_bht_update_valid = mem_reg_valid & _wb_reg_replay_T; // @[src/main/scala/rocket/RocketCore.scala 948:45]
  assign io_imem_flush_icache = wb_reg_valid & wb_ctrl_fence_i & ~io_dmem_s2_nack; // @[src/main/scala/rocket/RocketCore.scala 918:59]
  assign io_imem_progress = io_imem_progress_REG; // @[src/main/scala/rocket/RocketCore.scala 923:20]
  assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 969:41]
  assign io_dmem_req_bits_addr = {io_dmem_req_bits_addr_msb,alu_io_adder_out[38:0]}; // @[src/main/scala/rocket/RocketCore.scala 1169:8]
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag}; // @[src/main/scala/rocket/RocketCore.scala 972:25]
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd; // @[src/main/scala/rocket/RocketCore.scala 973:25]
  assign io_dmem_req_bits_size = ex_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 974:25]
  assign io_dmem_req_bits_signed = ~ex_reg_inst[14]; // @[src/main/scala/rocket/RocketCore.scala 975:30]
  assign io_dmem_req_bits_dprv = csr_io_status_dprv; // @[src/main/scala/rocket/RocketCore.scala 979:31]
  assign io_dmem_req_bits_dv = 1'h0; // @[src/main/scala/rocket/RocketCore.scala 980:37]
  assign io_dmem_s1_kill = dcache_kill_mem | take_pc_wb | mem_reg_xcpt | ~mem_reg_valid; // @[src/main/scala/rocket/RocketCore.scala 640:68]
  assign io_dmem_s1_data_data = mem_reg_rs2; // @[src/main/scala/rocket/RocketCore.scala 986:24]
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode; // @[src/main/scala/rocket/RocketCore.scala 794:15]
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn; // @[src/main/scala/rocket/RocketCore.scala 794:15]
  assign io_ptw_sfence_valid = io_imem_sfence_valid; // @[src/main/scala/rocket/RocketCore.scala 931:17]
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1; // @[src/main/scala/rocket/RocketCore.scala 931:17]
  assign io_ptw_status_prv = csr_io_status_prv; // @[src/main/scala/rocket/RocketCore.scala 798:17]
  assign io_ptw_status_mxr = csr_io_status_mxr; // @[src/main/scala/rocket/RocketCore.scala 798:17]
  assign io_ptw_status_sum = csr_io_status_sum; // @[src/main/scala/rocket/RocketCore.scala 798:17]
  assign io_rocc_cmd_valid = replay_wb_rocc & _io_imem_progress_T; // @[src/main/scala/rocket/RocketCore.scala 994:53]
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 288:16]
  assign ibuf_io_kill = take_pc_wb | take_pc_mem; // @[src/main/scala/rocket/RocketCore.scala 280:35]
  assign ibuf_io_inst_0_ready = ~ctrl_stalld; // @[src/main/scala/rocket/RocketCore.scala 933:28]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_ungated_clock = clock; // @[src/main/scala/rocket/RocketCore.scala 763:24]
  assign csr_io_hartid = io_hartid; // @[src/main/scala/rocket/RocketCore.scala 770:17]
  assign csr_io_rw_addr = wb_reg_inst[31:20]; // @[src/main/scala/rocket/RocketCore.scala 802:32]
  assign csr_io_rw_cmd = wb_ctrl_csr & _csr_io_rw_cmd_T_1; // @[src/main/scala/rocket/CSR.scala 185:9]
  assign csr_io_rw_wdata = wb_reg_wdata; // @[src/main/scala/rocket/RocketCore.scala 804:19]
  assign csr_io_decode_0_inst = ibuf_io_inst_0_bits_inst_bits; // @[src/main/scala/rocket/RocketCore.scala 764:25]
  assign csr_io_exception = wb_reg_xcpt | _T_93 | _T_95 | _T_97 | _T_99 | _T_105 | _T_107; // @[src/main/scala/rocket/RocketCore.scala 1152:26]
  assign csr_io_retire = wb_reg_valid & ~replay_wb & ~wb_xcpt; // @[src/main/scala/rocket/RocketCore.scala 739:45]
  assign csr_io_cause = wb_reg_xcpt ? wb_reg_cause : {{59'd0}, _T_121}; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  assign csr_io_pc = wb_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 776:13]
  assign csr_io_tval = tval_valid ? _csr_io_tval_T_1 : 40'h0; // @[src/main/scala/rocket/RocketCore.scala 783:21]
  assign csr_io_gva = wb_xcpt & (tval_dmem_addr & wb_reg_hls_or_dv); // @[src/main/scala/rocket/RocketCore.scala 782:25]
  assign csr_io_inst_0 = {_csr_io_inst_0_T_3,wb_reg_raw_inst[15:0]}; // @[src/main/scala/rocket/RocketCore.scala 768:46]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw; // @[src/main/scala/rocket/RocketCore.scala 420:13]
  assign alu_io_fn = ex_ctrl_alu_fn; // @[src/main/scala/rocket/RocketCore.scala 421:13]
  assign alu_io_in2 = 2'h1 == ex_ctrl_sel_alu2 ? $signed({{60{_ex_op2_T_1[3]}},_ex_op2_T_1}) : $signed(_ex_op2_T_5); // @[src/main/scala/rocket/RocketCore.scala 422:24]
  assign alu_io_in1 = 2'h2 == ex_ctrl_sel_alu1 ? $signed({{24{_ex_op1_T_1[39]}},_ex_op1_T_1}) : $signed(_ex_op1_T_3); // @[src/main/scala/rocket/RocketCore.scala 423:24]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = ex_reg_valid & ex_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 455:36]
  assign div_io_req_bits_fn = ex_ctrl_alu_fn; // @[src/main/scala/rocket/RocketCore.scala 457:22]
  assign div_io_req_bits_dw = ex_ctrl_alu_dw; // @[src/main/scala/rocket/RocketCore.scala 456:22]
  assign div_io_req_bits_in1 = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[src/main/scala/rocket/RocketCore.scala 406:14]
  assign div_io_req_bits_in2 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[src/main/scala/rocket/RocketCore.scala 406:14]
  assign div_io_req_bits_tag = ex_reg_inst[11:7]; // @[src/main/scala/rocket/RocketCore.scala 390:29]
  assign div_io_kill = killm_common & div_io_kill_REG; // @[src/main/scala/rocket/RocketCore.scala 641:31]
  assign div_io_resp_ready = dmem_resp_replay & dmem_resp_xpu ? 1'h0 : _ctrl_stalld_T_17 | wb_waddr == 5'h0; // @[src/main/scala/rocket/RocketCore.scala 710:21 730:44 731:23]
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_value_1 = rf_30; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_2 = rf_29; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_3 = rf_28; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_4 = rf_27; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_5 = rf_26; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_6 = rf_25; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_7 = rf_24; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_8 = rf_23; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_9 = rf_22; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_10 = rf_21; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_11 = rf_20; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_12 = rf_19; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_13 = rf_18; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_14 = rf_17; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_15 = rf_16; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_16 = rf_15; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_17 = rf_14; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_18 = rf_13; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_19 = rf_12; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_20 = rf_11; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_21 = rf_10; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_22 = rf_9; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_23 = rf_8; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_24 = rf_7; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_25 = rf_6; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_26 = rf_5; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_27 = rf_4; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_28 = rf_3; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_29 = rf_2; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_30 = rf_1; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_io_bits_value_31 = rf_0; // @[src/main/scala/rocket/RocketCore.scala 1212:{34,34}]
  assign difftest_module_1_clock = clock;
  assign difftest_module_1_reset = reset;
  assign difftest_module_1_io_valid = wb_wen | ll_wen; // @[src/main/scala/rocket/RocketCore.scala 741:23]
  assign difftest_module_1_io_bits_valid = wb_wen | ll_wen; // @[src/main/scala/rocket/RocketCore.scala 741:23]
  assign difftest_module_1_io_bits_address = ll_wen ? ll_waddr : wb_waddr; // @[src/main/scala/rocket/RocketCore.scala 742:21]
  assign difftest_module_1_io_bits_data = dmem_resp_valid & dmem_resp_xpu & dmem_resp_waddr != 5'h0 ?
    io_dmem_resp_bits_data : _rf_wdata_T_7; // @[src/main/scala/rocket/RocketCore.scala 743:21]
  assign difftest_module_2_clock = clock;
  assign difftest_module_2_reset = reset;
  assign difftest_module_2_io_bits_privilegeMode = csr_io_difftest_privilegeMode; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mstatus = csr_io_difftest_mstatus; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_sstatus = csr_io_difftest_sstatus; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mepc = csr_io_difftest_mepc; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_sepc = csr_io_difftest_sepc; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mtval = csr_io_difftest_mtval; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_stval = csr_io_difftest_stval; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mtvec = csr_io_difftest_mtvec; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_stvec = csr_io_difftest_stvec; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mcause = csr_io_difftest_mcause; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_scause = csr_io_difftest_scause; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_satp = csr_io_difftest_satp; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mip = csr_io_difftest_mip; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mie = csr_io_difftest_mie; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mscratch = csr_io_difftest_mscratch; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_sscratch = csr_io_difftest_sscratch; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_mideleg = csr_io_difftest_mideleg; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_2_io_bits_medeleg = csr_io_difftest_medeleg; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 833:14]
  assign difftest_module_3_clock = clock;
  assign difftest_module_3_reset = reset;
  assign difftest_module_3_io_bits_minstret = csr_io_snapshot_minstret; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 837:14]
  assign difftest_module_3_io_bits_mcycle = csr_io_snapshot_mcycle; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 837:14]
  assign difftest_delayer_clock = clock;
  assign difftest_delayer_reset = reset;
  assign difftest_delayer_i_valid = csr_io_trace_0_valid & ~(csr_io_trace_0_exception | csr_io_trace_0_interrupt); // @[src/main/scala/rocket/CSR.scala 236:30]
  assign difftest_delayer_i_skip = _rf_wdata_T_4 & csr_io_csrr_counter; // @[src/main/scala/rocket/RocketCore.scala 1092:47]
  assign difftest_delayer_i_rfwen = wb_ctrl_wxd; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 1095:20]
  assign difftest_delayer_i_fpwen = wb_ctrl_wfd; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 1096:20]
  assign difftest_delayer_i_wpdest = wb_reg_inst[11:7]; // @[src/main/scala/rocket/RocketCore.scala 392:29]
  assign difftest_delayer_i_wdest = {{3'd0}, wb_waddr}; // @[difftest/src/main/scala/Difftest.scala 466:27 src/main/scala/rocket/RocketCore.scala 1098:20]
  assign difftest_delayer_i_pc = {_coreMonitorBundle_pc_T_2,_coreMonitorBundle_pc_T}; // @[src/main/scala/util/package.scala 124:15]
  assign difftest_delayer_i_instr = csr_io_trace_0_insn; // @[src/main/scala/rocket/RocketCore.scala 1024:31 1040:26]
  assign difftest_delayer_i_special = {{6'd0}, _difftest_special_T}; // @[difftest/src/main/scala/Difftest.scala 466:27 difftest/src/main/scala/Bundles.scala 81:13]
  assign difftest_module_4_clock = clock;
  assign difftest_module_4_reset = reset;
  assign difftest_module_4_io_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 158:15]
  assign difftest_module_4_io_bits_valid = difftest_delayer_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_skip = difftest_delayer_o_skip; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_rfwen = difftest_delayer_o_rfwen; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_fpwen = difftest_delayer_o_fpwen; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_wpdest = difftest_delayer_o_wpdest; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_wdest = difftest_delayer_o_wdest; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_pc = difftest_delayer_o_pc; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_instr = difftest_delayer_o_instr; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_4_io_bits_special = difftest_delayer_o_special; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_delayer_1_clock = clock;
  assign difftest_delayer_1_reset = reset;
  assign difftest_delayer_1_i_valid = ll_wen_try & ll_waddr != 5'h0; // @[src/main/scala/rocket/RocketCore.scala 1116:34]
  assign difftest_delayer_1_i_address = dmem_resp_replay & dmem_resp_xpu ? dmem_resp_waddr : div_io_resp_bits_tag; // @[src/main/scala/rocket/RocketCore.scala 730:44 734:14 712:29]
  assign difftest_delayer_1_i_data = dmem_resp_valid & dmem_resp_xpu & dmem_resp_waddr != 5'h0 ? io_dmem_resp_bits_data
     : _rf_wdata_T_7; // @[src/main/scala/rocket/RocketCore.scala 743:21]
  assign difftest_delayer_1_i_nack = ~ll_wen; // @[src/main/scala/rocket/RocketCore.scala 1119:22]
  assign difftest_module_5_clock = clock;
  assign difftest_module_5_reset = reset;
  assign difftest_module_5_io_valid = difftest_delayer_1_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 158:15]
  assign difftest_module_5_io_bits_valid = difftest_delayer_1_o_valid; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_5_io_bits_address = difftest_delayer_1_o_address; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_5_io_bits_data = difftest_delayer_1_o_data; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign difftest_module_5_io_bits_nack = difftest_delayer_1_o_nack; // @[difftest/src/main/scala/Difftest.scala 157:19 159:14]
  assign PlusArgTimeout_clock = clock;
  assign PlusArgTimeout_reset = reset;
  assign PlusArgTimeout_io_count = csr_io_time[31:0]; // @[src/main/scala/util/PlusArg.scala 89:82]
  always @(posedge clock) begin
    if (unpause) begin // @[src/main/scala/rocket/RocketCore.scala 1003:18]
      id_reg_pause <= 1'h0; // @[src/main/scala/rocket/RocketCore.scala 1003:33]
    end else if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      id_reg_pause <= _GEN_186;
    end
    imem_might_request_reg <= ex_pc_valid | mem_pc_valid; // @[src/main/scala/rocket/RocketCore.scala 920:43]
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_fp <= id_ctrl_decoder_1; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_rocc <= id_ctrl_decoder_2; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_branch <= id_ctrl_decoder_3; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_jal <= id_ctrl_decoder_4; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_jalr <= id_ctrl_decoder_5; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_rxs2 <= id_ctrl_decoder_6; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_zbk <= id_ctrl_decoder_8; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_zkn <= id_ctrl_decoder_9; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_zks <= id_ctrl_decoder_10; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_xcpt) begin // @[src/main/scala/rocket/RocketCore.scala 479:20]
        if (|_T_39) begin // @[src/main/scala/rocket/RocketCore.scala 489:52]
          ex_ctrl_sel_alu2 <= 2'h0; // @[src/main/scala/rocket/RocketCore.scala 491:26]
        end else if (|_T_37) begin // @[src/main/scala/rocket/RocketCore.scala 484:34]
          ex_ctrl_sel_alu2 <= 2'h1; // @[src/main/scala/rocket/RocketCore.scala 486:26]
        end else begin
          ex_ctrl_sel_alu2 <= 2'h0; // @[src/main/scala/rocket/RocketCore.scala 483:24]
        end
      end else begin
        ex_ctrl_sel_alu2 <= id_ctrl_decoder_11; // @[src/main/scala/rocket/RocketCore.scala 474:13]
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_xcpt) begin // @[src/main/scala/rocket/RocketCore.scala 479:20]
        if (|_T_39) begin // @[src/main/scala/rocket/RocketCore.scala 489:52]
          ex_ctrl_sel_alu1 <= 2'h2; // @[src/main/scala/rocket/RocketCore.scala 490:26]
        end else if (|_T_37) begin // @[src/main/scala/rocket/RocketCore.scala 484:34]
          ex_ctrl_sel_alu1 <= 2'h2; // @[src/main/scala/rocket/RocketCore.scala 485:26]
        end else begin
          ex_ctrl_sel_alu1 <= 2'h1; // @[src/main/scala/rocket/RocketCore.scala 482:24]
        end
      end else begin
        ex_ctrl_sel_alu1 <= id_ctrl_decoder_12; // @[src/main/scala/rocket/RocketCore.scala 474:13]
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_sel_imm <= id_ctrl_decoder_13; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_alu_dw <= _GEN_194;
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_xcpt) begin // @[src/main/scala/rocket/RocketCore.scala 479:20]
        ex_ctrl_alu_fn <= 4'h0; // @[src/main/scala/rocket/RocketCore.scala 480:22]
      end else begin
        ex_ctrl_alu_fn <= id_ctrl_decoder_15; // @[src/main/scala/rocket/RocketCore.scala 474:13]
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_mem <= id_ctrl_decoder_16; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_mem_cmd <= id_ctrl_decoder_17;
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_wfd <= id_ctrl_decoder_21; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_mul <= id_ctrl_decoder_22; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_div <= id_ctrl_decoder_23; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_wxd <= id_ctrl_decoder_24; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_system_insn & id_ctrl_decoder_16) begin // @[src/main/scala/rocket/RocketCore.scala 317:19]
        ex_ctrl_csr <= 3'h0;
      end else if (id_csr_ren) begin // @[src/main/scala/rocket/RocketCore.scala 317:61]
        ex_ctrl_csr <= 3'h2;
      end else begin
        ex_ctrl_csr <= id_ctrl_decoder_25;
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_ctrl_fence_i <= id_ctrl_decoder_26; // @[src/main/scala/rocket/RocketCore.scala 474:13]
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_fp <= ex_ctrl_fp; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_rocc <= ex_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_branch <= ex_ctrl_branch; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_jal <= ex_ctrl_jal; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_jalr <= ex_ctrl_jalr; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_mem <= ex_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_wfd <= ex_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_mul <= ex_ctrl_mul; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_div <= ex_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_wxd <= ex_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_csr <= ex_ctrl_csr; // @[src/main/scala/rocket/RocketCore.scala 582:14]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_ctrl_fence_i <= _GEN_263;
      end
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_rocc <= mem_ctrl_rocc; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_mem <= mem_ctrl_mem; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_wfd <= mem_ctrl_wfd; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_div <= mem_ctrl_div; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_wxd <= mem_ctrl_wxd; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_csr <= mem_ctrl_csr; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_ctrl_fence_i <= mem_ctrl_fence_i; // @[src/main/scala/rocket/RocketCore.scala 650:13]
    end
    ex_reg_xcpt_interrupt <= _ex_reg_replay_T_1 & csr_io_interrupt; // @[src/main/scala/rocket/RocketCore.scala 471:62]
    ex_reg_valid <= ~ctrl_killd; // @[src/main/scala/rocket/RocketCore.scala 468:19]
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_xcpt) begin // @[src/main/scala/rocket/RocketCore.scala 479:20]
        ex_reg_rvc <= _GEN_190;
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc; // @[src/main/scala/rocket/RocketCore.scala 475:16]
      end
    end
    ex_reg_xcpt <= _ex_reg_valid_T & id_xcpt; // @[src/main/scala/rocket/RocketCore.scala 470:30]
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_reg_flush_pipe <= id_ctrl_decoder_26 | id_csr_flush; // @[src/main/scala/rocket/RocketCore.scala 494:23]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_reg_load_use <= id_load_use; // @[src/main/scala/rocket/RocketCore.scala 495:21]
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin // @[src/main/scala/rocket/RocketCore.scala 527:73]
      if (csr_io_interrupt) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        ex_reg_cause <= csr_io_interrupt_cause;
      end else begin
        ex_reg_cause <= {{59'd0}, _T_16};
      end
    end
    ex_reg_replay <= ~take_pc_mem_wb & ibuf_io_inst_0_valid & ibuf_io_inst_0_bits_replay; // @[src/main/scala/rocket/RocketCore.scala 469:54]
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin // @[src/main/scala/rocket/RocketCore.scala 527:73]
      ex_reg_pc <= ibuf_io_pc; // @[src/main/scala/rocket/RocketCore.scala 531:15]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (_T_48) begin // @[src/main/scala/rocket/RocketCore.scala 498:81]
        ex_reg_mem_size <= _ex_reg_mem_size_T_6; // @[src/main/scala/rocket/RocketCore.scala 499:23]
      end else begin
        ex_reg_mem_size <= ibuf_io_inst_0_bits_inst_bits[13:12]; // @[src/main/scala/rocket/RocketCore.scala 497:21]
      end
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin // @[src/main/scala/rocket/RocketCore.scala 527:73]
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits; // @[src/main/scala/rocket/RocketCore.scala 529:17]
    end
    if (_ex_reg_valid_T | csr_io_interrupt | ibuf_io_inst_0_bits_replay) begin // @[src/main/scala/rocket/RocketCore.scala 527:73]
      ex_reg_raw_inst <= ibuf_io_inst_0_bits_raw; // @[src/main/scala/rocket/RocketCore.scala 530:21]
    end
    mem_reg_xcpt_interrupt <= _ex_reg_replay_T & ex_reg_xcpt_interrupt; // @[src/main/scala/rocket/RocketCore.scala 575:45]
    mem_reg_valid <= ~ctrl_killx; // @[src/main/scala/rocket/RocketCore.scala 572:20]
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_rvc <= ex_reg_rvc; // @[src/main/scala/rocket/RocketCore.scala 583:17]
      end
    end
    mem_reg_xcpt <= _mem_reg_valid_T & ex_xcpt; // @[src/main/scala/rocket/RocketCore.scala 574:31]
    mem_reg_replay <= _ex_reg_replay_T & replay_ex; // @[src/main/scala/rocket/RocketCore.scala 573:37]
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_flush_pipe <= _GEN_264;
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_cause <= ex_reg_cause; // @[src/main/scala/rocket/RocketCore.scala 592:19]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_slow_bypass <= ex_slow_bypass; // @[src/main/scala/rocket/RocketCore.scala 589:25]
      end
    end
    if (mem_reg_valid & mem_reg_flush_pipe) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      mem_reg_sfence <= 1'h0; // @[src/main/scala/rocket/RocketCore.scala 580:20]
    end else if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
      mem_reg_sfence <= ex_sfence; // @[src/main/scala/rocket/RocketCore.scala 586:20]
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_pc <= ex_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 597:16]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_inst <= ex_reg_inst; // @[src/main/scala/rocket/RocketCore.scala 593:18]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_mem_size <= ex_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 595:22]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_hls_or_dv <= io_dmem_req_bits_dv; // @[src/main/scala/rocket/RocketCore.scala 596:23]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_reg_raw_inst <= ex_reg_raw_inst; // @[src/main/scala/rocket/RocketCore.scala 594:22]
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        if (_mem_reg_wdata_T_4) begin // @[src/main/scala/chisel3/util/Mux.scala 30:73]
          mem_reg_wdata <= alu_io_out;
        end else begin
          mem_reg_wdata <= 64'h0;
        end
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        if (ex_ctrl_rxs2 & (ex_ctrl_mem | ex_ctrl_rocc | ex_sfence)) begin // @[src/main/scala/rocket/RocketCore.scala 608:71]
          if (size == 2'h0) begin // @[src/main/scala/rocket/AMOALU.scala 28:13]
            mem_reg_rs2 <= _mem_reg_rs2_T_4;
          end else begin
            mem_reg_rs2 <= _mem_reg_rs2_T_13;
          end
        end
      end
    end
    if (!(mem_reg_valid & mem_reg_flush_pipe)) begin // @[src/main/scala/rocket/RocketCore.scala 579:46]
      if (ex_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 581:28]
        mem_br_taken <= alu_io_cmp_out; // @[src/main/scala/rocket/RocketCore.scala 606:18]
      end
    end
    wb_reg_valid <= ~ctrl_killm; // @[src/main/scala/rocket/RocketCore.scala 645:19]
    wb_reg_xcpt <= mem_xcpt & _wb_reg_replay_T; // @[src/main/scala/rocket/RocketCore.scala 647:27]
    wb_reg_replay <= replay_mem & ~take_pc_wb; // @[src/main/scala/rocket/RocketCore.scala 646:31]
    wb_reg_flush_pipe <= _wb_reg_valid_T & mem_reg_flush_pipe; // @[src/main/scala/rocket/RocketCore.scala 648:36]
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      if (_T_74) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{60'd0}, _T_78};
      end
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_sfence <= mem_reg_sfence; // @[src/main/scala/rocket/RocketCore.scala 651:19]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_pc <= mem_reg_pc; // @[src/main/scala/rocket/RocketCore.scala 663:15]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_mem_size <= mem_reg_mem_size; // @[src/main/scala/rocket/RocketCore.scala 659:21]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_hls_or_dv <= mem_reg_hls_or_dv; // @[src/main/scala/rocket/RocketCore.scala 660:22]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_inst <= mem_reg_inst; // @[src/main/scala/rocket/RocketCore.scala 657:17]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      wb_reg_raw_inst <= mem_reg_raw_inst; // @[src/main/scala/rocket/RocketCore.scala 658:21]
    end
    if (mem_pc_valid) begin // @[src/main/scala/rocket/RocketCore.scala 649:23]
      if (_take_pc_mem_T & mem_ctrl_fp & mem_ctrl_wxd) begin // @[src/main/scala/rocket/RocketCore.scala 652:24]
        wb_reg_wdata <= 64'h0;
      end else begin
        wb_reg_wdata <= mem_int_wdata;
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 305:29]
      id_reg_fence <= 1'h0; // @[src/main/scala/rocket/RocketCore.scala 305:29]
    end else if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      id_reg_fence <= _GEN_187;
    end else if (~id_mem_busy) begin // @[src/main/scala/rocket/RocketCore.scala 344:23]
      id_reg_fence <= 1'h0; // @[src/main/scala/rocket/RocketCore.scala 344:38]
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_0 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h0 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_0 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_1 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_1 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_2 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h2 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_2 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_3 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h3 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_3 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_4 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h4 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_4 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_5 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h5 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_5 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_6 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h6 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_6 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_7 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h7 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_7 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_8 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h8 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_8 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_9 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h9 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_9 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_10 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'ha == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_10 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_11 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'hb == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_11 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_12 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'hc == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_12 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_13 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'hd == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_13 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_14 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'he == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_14 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_15 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'hf == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_15 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_16 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h10 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_16 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_17 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h11 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_17 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_18 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h12 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_18 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_19 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h13 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_19 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_20 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h14 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_20 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_21 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h15 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_21 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_22 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h16 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_22 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_23 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h17 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_23 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_24 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h18 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_24 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_25 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h19 == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_25 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_26 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1a == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_26 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_27 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1b == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_27 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_28 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1c == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_28 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_29 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1d == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_29 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1194:19]
      rf_30 <= 64'h0; // @[src/main/scala/rocket/RocketCore.scala 1194:19]
    end else if (rf_wen) begin // @[src/main/scala/rocket/RocketCore.scala 748:17]
      if (rf_waddr != 5'h0) begin // @[src/main/scala/rocket/RocketCore.scala 1206:25]
        if (5'h1e == _T_137) begin // @[src/main/scala/rocket/RocketCore.scala 1207:20]
          rf_30 <= rf_wdata; // @[src/main/scala/rocket/RocketCore.scala 1207:20]
        end
      end
    end
    line_1117_valid_reg <= 5'h0 == _id_rs_T_3;
    line_1118_valid_reg <= 5'h1 == _id_rs_T_3;
    line_1119_valid_reg <= 5'h2 == _id_rs_T_3;
    line_1120_valid_reg <= 5'h3 == _id_rs_T_3;
    line_1121_valid_reg <= 5'h4 == _id_rs_T_3;
    line_1122_valid_reg <= 5'h5 == _id_rs_T_3;
    line_1123_valid_reg <= 5'h6 == _id_rs_T_3;
    line_1124_valid_reg <= 5'h7 == _id_rs_T_3;
    line_1125_valid_reg <= 5'h8 == _id_rs_T_3;
    line_1126_valid_reg <= 5'h9 == _id_rs_T_3;
    line_1127_valid_reg <= 5'ha == _id_rs_T_3;
    line_1128_valid_reg <= 5'hb == _id_rs_T_3;
    line_1129_valid_reg <= 5'hc == _id_rs_T_3;
    line_1130_valid_reg <= 5'hd == _id_rs_T_3;
    line_1131_valid_reg <= 5'he == _id_rs_T_3;
    line_1132_valid_reg <= 5'hf == _id_rs_T_3;
    line_1133_valid_reg <= 5'h10 == _id_rs_T_3;
    line_1134_valid_reg <= 5'h11 == _id_rs_T_3;
    line_1135_valid_reg <= 5'h12 == _id_rs_T_3;
    line_1136_valid_reg <= 5'h13 == _id_rs_T_3;
    line_1137_valid_reg <= 5'h14 == _id_rs_T_3;
    line_1138_valid_reg <= 5'h15 == _id_rs_T_3;
    line_1139_valid_reg <= 5'h16 == _id_rs_T_3;
    line_1140_valid_reg <= 5'h17 == _id_rs_T_3;
    line_1141_valid_reg <= 5'h18 == _id_rs_T_3;
    line_1142_valid_reg <= 5'h19 == _id_rs_T_3;
    line_1143_valid_reg <= 5'h1a == _id_rs_T_3;
    line_1144_valid_reg <= 5'h1b == _id_rs_T_3;
    line_1145_valid_reg <= 5'h1c == _id_rs_T_3;
    line_1146_valid_reg <= 5'h1d == _id_rs_T_3;
    line_1147_valid_reg <= 5'h1e == _id_rs_T_3;
    line_1148_valid_reg <= 5'h0 == _id_rs_T_8;
    line_1149_valid_reg <= 5'h1 == _id_rs_T_8;
    line_1150_valid_reg <= 5'h2 == _id_rs_T_8;
    line_1151_valid_reg <= 5'h3 == _id_rs_T_8;
    line_1152_valid_reg <= 5'h4 == _id_rs_T_8;
    line_1153_valid_reg <= 5'h5 == _id_rs_T_8;
    line_1154_valid_reg <= 5'h6 == _id_rs_T_8;
    line_1155_valid_reg <= 5'h7 == _id_rs_T_8;
    line_1156_valid_reg <= 5'h8 == _id_rs_T_8;
    line_1157_valid_reg <= 5'h9 == _id_rs_T_8;
    line_1158_valid_reg <= 5'ha == _id_rs_T_8;
    line_1159_valid_reg <= 5'hb == _id_rs_T_8;
    line_1160_valid_reg <= 5'hc == _id_rs_T_8;
    line_1161_valid_reg <= 5'hd == _id_rs_T_8;
    line_1162_valid_reg <= 5'he == _id_rs_T_8;
    line_1163_valid_reg <= 5'hf == _id_rs_T_8;
    line_1164_valid_reg <= 5'h10 == _id_rs_T_8;
    line_1165_valid_reg <= 5'h11 == _id_rs_T_8;
    line_1166_valid_reg <= 5'h12 == _id_rs_T_8;
    line_1167_valid_reg <= 5'h13 == _id_rs_T_8;
    line_1168_valid_reg <= 5'h14 == _id_rs_T_8;
    line_1169_valid_reg <= 5'h15 == _id_rs_T_8;
    line_1170_valid_reg <= 5'h16 == _id_rs_T_8;
    line_1171_valid_reg <= 5'h17 == _id_rs_T_8;
    line_1172_valid_reg <= 5'h18 == _id_rs_T_8;
    line_1173_valid_reg <= 5'h19 == _id_rs_T_8;
    line_1174_valid_reg <= 5'h1a == _id_rs_T_8;
    line_1175_valid_reg <= 5'h1b == _id_rs_T_8;
    line_1176_valid_reg <= 5'h1c == _id_rs_T_8;
    line_1177_valid_reg <= 5'h1d == _id_rs_T_8;
    line_1178_valid_reg <= 5'h1e == _id_rs_T_8;
    line_1179_valid_reg <= _T;
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_illegal_insn) begin // @[src/main/scala/rocket/RocketCore.scala 520:47]
        ex_reg_rs_bypass_0 <= 1'h0; // @[src/main/scala/rocket/RocketCore.scala 522:27]
      end else begin
        ex_reg_rs_bypass_0 <= do_bypass; // @[src/main/scala/rocket/RocketCore.scala 513:27]
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      ex_reg_rs_bypass_1 <= do_bypass_1; // @[src/main/scala/rocket/RocketCore.scala 513:27]
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_illegal_insn) begin // @[src/main/scala/rocket/RocketCore.scala 520:47]
        ex_reg_rs_lsb_0 <= inst[1:0]; // @[src/main/scala/rocket/RocketCore.scala 523:24]
      end else if (id_ctrl_decoder_7 & ~do_bypass) begin // @[src/main/scala/rocket/RocketCore.scala 515:38]
        ex_reg_rs_lsb_0 <= id_rs_0[1:0]; // @[src/main/scala/rocket/RocketCore.scala 516:26]
      end else if (id_bypass_src_0_0) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        ex_reg_rs_lsb_0 <= 2'h0;
      end else begin
        ex_reg_rs_lsb_0 <= _bypass_src_T_1;
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_ctrl_decoder_6 & ~do_bypass_1) begin // @[src/main/scala/rocket/RocketCore.scala 515:38]
        ex_reg_rs_lsb_1 <= id_rs_1[1:0]; // @[src/main/scala/rocket/RocketCore.scala 516:26]
      end else if (id_bypass_src_1_0) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        ex_reg_rs_lsb_1 <= 2'h0;
      end else if (id_bypass_src_1_1) begin // @[src/main/scala/chisel3/util/Mux.scala 50:70]
        ex_reg_rs_lsb_1 <= 2'h1;
      end else begin
        ex_reg_rs_lsb_1 <= _bypass_src_T_2;
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_illegal_insn) begin // @[src/main/scala/rocket/RocketCore.scala 520:47]
        ex_reg_rs_msb_0 <= {{32'd0}, inst[31:2]}; // @[src/main/scala/rocket/RocketCore.scala 524:24]
      end else if (id_ctrl_decoder_7 & ~do_bypass) begin // @[src/main/scala/rocket/RocketCore.scala 515:38]
        ex_reg_rs_msb_0 <= id_rs_0[63:2]; // @[src/main/scala/rocket/RocketCore.scala 517:26]
      end
    end
    if (_ex_reg_valid_T) begin // @[src/main/scala/rocket/RocketCore.scala 473:22]
      if (id_ctrl_decoder_6 & ~do_bypass_1) begin // @[src/main/scala/rocket/RocketCore.scala 515:38]
        ex_reg_rs_msb_1 <= id_rs_1[63:2]; // @[src/main/scala/rocket/RocketCore.scala 517:26]
      end
    end
    if (reset) begin // @[src/main/scala/rocket/RocketCore.scala 1179:32]
      reg_r <= 32'h0; // @[src/main/scala/rocket/RocketCore.scala 1179:32]
    end else if (_T_155) begin // @[src/main/scala/rocket/RocketCore.scala 1187:18]
      reg_r <= _T_154; // @[src/main/scala/rocket/RocketCore.scala 1187:26]
    end else if (ll_wen) begin // @[src/main/scala/rocket/RocketCore.scala 1187:18]
      reg_r <= _T_149; // @[src/main/scala/rocket/RocketCore.scala 1187:26]
    end
    dcache_blocked_blocked <= _replay_ex_structural_T & _dcache_blocked_T & (dcache_blocked_blocked | io_dmem_req_valid
       | io_dmem_s2_nack); // @[src/main/scala/rocket/RocketCore.scala 891:83]
    rocc_blocked <= _wb_valid_T_2 & (io_rocc_cmd_valid | rocc_blocked); // @[src/main/scala/rocket/RocketCore.scala 895:50]
    line_1180_valid_reg <= _ex_reg_valid_T;
    line_1181_valid_reg <= _T_36;
    line_1182_valid_reg <= id_fence_next;
    line_1183_valid_reg <= id_xcpt;
    line_1184_valid_reg <= _T_38;
    line_1185_valid_reg <= _T_40;
    line_1186_valid_reg <= _T_48;
    line_1187_valid_reg <= _T_52;
    line_1188_valid_reg <= _T_54;
    line_1189_valid_reg <= id_illegal_insn;
    line_1190_valid_reg <= _T_58;
    line_1191_valid_reg <= _T_69;
    line_1192_valid_reg <= _T_69;
    line_1193_valid_reg <= ex_pc_valid;
    line_1194_valid_reg <= _T_72;
    line_1195_valid_reg <= _T_73;
    div_io_kill_REG <= div_io_req_ready & div_io_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    line_1196_valid_reg <= mem_pc_valid;
    line_1197_valid_reg <= _T_91;
    line_1198_valid_reg <= _T_134;
    line_1199_valid_reg <= rf_wen;
    line_1200_valid_reg <= _T_135;
    line_1201_valid_reg <= 5'h0 == _T_137;
    line_1202_valid_reg <= 5'h1 == _T_137;
    line_1203_valid_reg <= 5'h2 == _T_137;
    line_1204_valid_reg <= 5'h3 == _T_137;
    line_1205_valid_reg <= 5'h4 == _T_137;
    line_1206_valid_reg <= 5'h5 == _T_137;
    line_1207_valid_reg <= 5'h6 == _T_137;
    line_1208_valid_reg <= 5'h7 == _T_137;
    line_1209_valid_reg <= 5'h8 == _T_137;
    line_1210_valid_reg <= 5'h9 == _T_137;
    line_1211_valid_reg <= 5'ha == _T_137;
    line_1212_valid_reg <= 5'hb == _T_137;
    line_1213_valid_reg <= 5'hc == _T_137;
    line_1214_valid_reg <= 5'hd == _T_137;
    line_1215_valid_reg <= 5'he == _T_137;
    line_1216_valid_reg <= 5'hf == _T_137;
    line_1217_valid_reg <= 5'h10 == _T_137;
    line_1218_valid_reg <= 5'h11 == _T_137;
    line_1219_valid_reg <= 5'h12 == _T_137;
    line_1220_valid_reg <= 5'h13 == _T_137;
    line_1221_valid_reg <= 5'h14 == _T_137;
    line_1222_valid_reg <= 5'h15 == _T_137;
    line_1223_valid_reg <= 5'h16 == _T_137;
    line_1224_valid_reg <= 5'h17 == _T_137;
    line_1225_valid_reg <= 5'h18 == _T_137;
    line_1226_valid_reg <= 5'h19 == _T_137;
    line_1227_valid_reg <= 5'h1a == _T_137;
    line_1228_valid_reg <= 5'h1b == _T_137;
    line_1229_valid_reg <= 5'h1c == _T_137;
    line_1230_valid_reg <= 5'h1d == _T_137;
    line_1231_valid_reg <= 5'h1e == _T_137;
    line_1232_valid_reg <= _T_138;
    line_1233_valid_reg <= _T_139;
    line_1234_valid_reg <= _csr_io_htval_T_3;
    line_1235_valid_reg <= _csr_io_htval_T_4;
    line_1236_valid_reg <= ll_wen;
    line_1237_valid_reg <= _T_155;
    io_imem_progress_REG <= wb_reg_valid & ~replay_wb_common; // @[src/main/scala/rocket/RocketCore.scala 923:44]
    line_1238_valid_reg <= unpause;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~csr_io_htval_htval_valid_imem)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at RocketCore.scala:787 assert(!htval_valid_imem || io.imem.gpa.valid)\n"); // @[src/main/scala/rocket/RocketCore.scala 787:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  id_reg_pause = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  imem_might_request_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ex_ctrl_fp = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ex_ctrl_rocc = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_rxs2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_zbk = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_zkn = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_zks = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_alu_dw = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  ex_ctrl_wfd = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ex_ctrl_mul = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ex_ctrl_div = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ex_ctrl_csr = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  ex_ctrl_fence_i = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  mem_ctrl_fp = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_rocc = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_wfd = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_mul = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  mem_ctrl_csr = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  mem_ctrl_fence_i = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  wb_ctrl_rocc = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  wb_ctrl_wfd = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  wb_ctrl_div = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  wb_ctrl_csr = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  wb_ctrl_fence_i = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  ex_reg_xcpt_interrupt = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  ex_reg_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  ex_reg_rvc = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ex_reg_xcpt = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ex_reg_flush_pipe = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  ex_reg_load_use = _RAND_48[0:0];
  _RAND_49 = {2{`RANDOM}};
  ex_reg_cause = _RAND_49[63:0];
  _RAND_50 = {1{`RANDOM}};
  ex_reg_replay = _RAND_50[0:0];
  _RAND_51 = {2{`RANDOM}};
  ex_reg_pc = _RAND_51[39:0];
  _RAND_52 = {1{`RANDOM}};
  ex_reg_mem_size = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  ex_reg_inst = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  ex_reg_raw_inst = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  mem_reg_xcpt_interrupt = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  mem_reg_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  mem_reg_rvc = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  mem_reg_xcpt = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mem_reg_replay = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  mem_reg_flush_pipe = _RAND_60[0:0];
  _RAND_61 = {2{`RANDOM}};
  mem_reg_cause = _RAND_61[63:0];
  _RAND_62 = {1{`RANDOM}};
  mem_reg_slow_bypass = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  mem_reg_sfence = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  mem_reg_pc = _RAND_64[39:0];
  _RAND_65 = {1{`RANDOM}};
  mem_reg_inst = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mem_reg_mem_size = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  mem_reg_hls_or_dv = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  mem_reg_raw_inst = _RAND_68[31:0];
  _RAND_69 = {2{`RANDOM}};
  mem_reg_wdata = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  mem_reg_rs2 = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  mem_br_taken = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  wb_reg_valid = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  wb_reg_xcpt = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  wb_reg_replay = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  wb_reg_flush_pipe = _RAND_75[0:0];
  _RAND_76 = {2{`RANDOM}};
  wb_reg_cause = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  wb_reg_sfence = _RAND_77[0:0];
  _RAND_78 = {2{`RANDOM}};
  wb_reg_pc = _RAND_78[39:0];
  _RAND_79 = {1{`RANDOM}};
  wb_reg_mem_size = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  wb_reg_hls_or_dv = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  wb_reg_inst = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  wb_reg_raw_inst = _RAND_82[31:0];
  _RAND_83 = {2{`RANDOM}};
  wb_reg_wdata = _RAND_83[63:0];
  _RAND_84 = {1{`RANDOM}};
  id_reg_fence = _RAND_84[0:0];
  _RAND_85 = {2{`RANDOM}};
  rf_0 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  rf_1 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  rf_2 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  rf_3 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  rf_4 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  rf_5 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  rf_6 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  rf_7 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  rf_8 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  rf_9 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  rf_10 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  rf_11 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  rf_12 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  rf_13 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  rf_14 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  rf_15 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  rf_16 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  rf_17 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  rf_18 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  rf_19 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  rf_20 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  rf_21 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  rf_22 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  rf_23 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  rf_24 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  rf_25 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  rf_26 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  rf_27 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  rf_28 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  rf_29 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  rf_30 = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  line_1117_valid_reg = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  line_1118_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  line_1119_valid_reg = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  line_1120_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  line_1121_valid_reg = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  line_1122_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  line_1123_valid_reg = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  line_1124_valid_reg = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  line_1125_valid_reg = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  line_1126_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  line_1127_valid_reg = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  line_1128_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  line_1129_valid_reg = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  line_1130_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  line_1131_valid_reg = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  line_1132_valid_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  line_1133_valid_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  line_1134_valid_reg = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  line_1135_valid_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  line_1136_valid_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  line_1137_valid_reg = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  line_1138_valid_reg = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  line_1139_valid_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  line_1140_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  line_1141_valid_reg = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  line_1142_valid_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  line_1143_valid_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  line_1144_valid_reg = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  line_1145_valid_reg = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  line_1146_valid_reg = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  line_1147_valid_reg = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  line_1148_valid_reg = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  line_1149_valid_reg = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  line_1150_valid_reg = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  line_1151_valid_reg = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  line_1152_valid_reg = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  line_1153_valid_reg = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  line_1154_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  line_1155_valid_reg = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  line_1156_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  line_1157_valid_reg = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  line_1158_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  line_1159_valid_reg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  line_1160_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  line_1161_valid_reg = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  line_1162_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  line_1163_valid_reg = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  line_1164_valid_reg = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  line_1165_valid_reg = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  line_1166_valid_reg = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  line_1167_valid_reg = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  line_1168_valid_reg = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  line_1169_valid_reg = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  line_1170_valid_reg = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  line_1171_valid_reg = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  line_1172_valid_reg = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  line_1173_valid_reg = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  line_1174_valid_reg = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  line_1175_valid_reg = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  line_1176_valid_reg = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  line_1177_valid_reg = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  line_1178_valid_reg = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  line_1179_valid_reg = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ex_reg_rs_bypass_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ex_reg_rs_bypass_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ex_reg_rs_lsb_0 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  ex_reg_rs_lsb_1 = _RAND_182[1:0];
  _RAND_183 = {2{`RANDOM}};
  ex_reg_rs_msb_0 = _RAND_183[61:0];
  _RAND_184 = {2{`RANDOM}};
  ex_reg_rs_msb_1 = _RAND_184[61:0];
  _RAND_185 = {1{`RANDOM}};
  reg_r = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  dcache_blocked_blocked = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  rocc_blocked = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  line_1180_valid_reg = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  line_1181_valid_reg = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  line_1182_valid_reg = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  line_1183_valid_reg = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  line_1184_valid_reg = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  line_1185_valid_reg = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  line_1186_valid_reg = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  line_1187_valid_reg = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  line_1188_valid_reg = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  line_1189_valid_reg = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  line_1190_valid_reg = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  line_1191_valid_reg = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  line_1192_valid_reg = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  line_1193_valid_reg = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  line_1194_valid_reg = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  line_1195_valid_reg = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  div_io_kill_REG = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  line_1196_valid_reg = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  line_1197_valid_reg = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  line_1198_valid_reg = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  line_1199_valid_reg = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  line_1200_valid_reg = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  line_1201_valid_reg = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  line_1202_valid_reg = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  line_1203_valid_reg = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  line_1204_valid_reg = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  line_1205_valid_reg = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  line_1206_valid_reg = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  line_1207_valid_reg = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  line_1208_valid_reg = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  line_1209_valid_reg = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  line_1210_valid_reg = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  line_1211_valid_reg = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  line_1212_valid_reg = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  line_1213_valid_reg = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  line_1214_valid_reg = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  line_1215_valid_reg = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  line_1216_valid_reg = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  line_1217_valid_reg = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  line_1218_valid_reg = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  line_1219_valid_reg = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  line_1220_valid_reg = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  line_1221_valid_reg = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  line_1222_valid_reg = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  line_1223_valid_reg = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  line_1224_valid_reg = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  line_1225_valid_reg = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  line_1226_valid_reg = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  line_1227_valid_reg = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  line_1228_valid_reg = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  line_1229_valid_reg = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  line_1230_valid_reg = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  line_1231_valid_reg = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  line_1232_valid_reg = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  line_1233_valid_reg = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  line_1234_valid_reg = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  line_1235_valid_reg = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  line_1236_valid_reg = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  line_1237_valid_reg = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  io_imem_progress_REG = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  line_1238_valid_reg = _RAND_248[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~csr_io_htval_htval_valid_imem); // @[src/main/scala/rocket/RocketCore.scala 787:11]
    end
  end
endmodule
module RocketTile(
  input         clock,
  input         reset,
  input         auto_buffer_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_buffer_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_buffer_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_buffer_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_buffer_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_buffer_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_buffer_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_buffer_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_buffer_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_buffer_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_buffer_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_buffer_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_buffer_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_buffer_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_buffer_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_buffer_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_buffer_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_buffer_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_buffer_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_buffer_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_buffer_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_buffer_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_buffer_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_buffer_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_buffer_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_buffer_out_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_hartid_in // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  tlMasterXbar_clock; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_reset; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_1_a_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_1_a_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_in_1_a_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_1_d_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_in_1_d_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_1_d_bits_corrupt; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_a_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_a_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_a_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_in_0_a_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_in_0_a_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_b_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_b_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_b_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_b_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_in_0_b_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_c_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_c_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_c_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_in_0_c_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_in_0_c_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_d_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_d_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_d_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_d_bits_denied; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_in_0_d_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_e_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_in_0_e_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_a_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_a_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_a_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_out_a_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_out_a_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_b_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_b_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_out_b_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_c_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_c_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_c_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [31:0] tlMasterXbar_auto_out_c_bits_address; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_out_c_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_d_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_d_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_param; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_size; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_source; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_sink; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_d_bits_denied; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [63:0] tlMasterXbar_auto_out_d_bits_data; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_d_bits_corrupt; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_e_ready; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlMasterXbar_auto_out_e_valid; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire [1:0] tlMasterXbar_auto_out_e_bits_sink; // @[src/main/scala/tile/BaseTile.scala 224:42]
  wire  tlSlaveXbar_clock; // @[src/main/scala/tile/BaseTile.scala 225:41]
  wire  tlSlaveXbar_reset; // @[src/main/scala/tile/BaseTile.scala 225:41]
  wire  intXbar_clock; // @[src/main/scala/tile/BaseTile.scala 226:37]
  wire  intXbar_reset; // @[src/main/scala/tile/BaseTile.scala 226:37]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_auto_in; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_auto_out; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_1_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_1_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_2_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_2_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  nexus_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
  wire  nexus_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
  wire  broadcast_3_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_3_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  nexus_1_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
  wire  nexus_1_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
  wire  broadcast_4_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_4_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  widget_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_b_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_b_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_b_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_b_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_b_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_b_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_c_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_c_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_c_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_c_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_c_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_c_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_e_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_in_e_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_e_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_a_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [7:0] widget_auto_out_a_bits_mask; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_a_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_b_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_b_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_b_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_b_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_b_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_b_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_c_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_c_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_c_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_c_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_c_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_c_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_param; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_source; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_d_bits_denied; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_e_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_auto_out_e_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_e_bits_sink; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  dcache_clock; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_reset; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_a_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_a_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_a_bits_opcode; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_a_bits_param; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_a_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_a_bits_source; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [31:0] dcache_auto_out_a_bits_address; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [7:0] dcache_auto_out_a_bits_mask; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_auto_out_a_bits_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_b_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_b_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_auto_out_b_bits_param; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_b_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_b_bits_source; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [31:0] dcache_auto_out_b_bits_address; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_c_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_c_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_c_bits_param; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_c_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_c_bits_source; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [31:0] dcache_auto_out_c_bits_address; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_auto_out_c_bits_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_d_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_d_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_d_bits_opcode; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_auto_out_d_bits_param; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [2:0] dcache_auto_out_d_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_d_bits_source; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_auto_out_d_bits_sink; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_d_bits_denied; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_auto_out_d_bits_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_e_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_auto_out_e_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_auto_out_e_bits_sink; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_req_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_req_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [39:0] dcache_io_cpu_req_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [6:0] dcache_io_cpu_req_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [4:0] dcache_io_cpu_req_bits_cmd; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_io_cpu_req_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_req_bits_signed; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_io_cpu_req_bits_dprv; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_req_bits_phys; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s1_kill; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_io_cpu_s1_data_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [7:0] dcache_io_cpu_s1_data_mask; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_nack; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [39:0] dcache_io_cpu_resp_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [6:0] dcache_io_cpu_resp_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [4:0] dcache_io_cpu_resp_bits_cmd; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_io_cpu_resp_bits_size; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_resp_bits_signed; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_io_cpu_resp_bits_dprv; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_resp_bits_dv; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_io_cpu_resp_bits_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [7:0] dcache_io_cpu_resp_bits_mask; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_resp_bits_replay; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_resp_bits_has_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_io_cpu_resp_bits_data_word_bypass; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_io_cpu_resp_bits_data_raw; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [63:0] dcache_io_cpu_resp_bits_store_data; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_replay_next; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_ma_ld; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_ma_st; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_pf_ld; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_pf_st; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_gf_ld; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_gf_st; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_s2_xcpt_ae_st; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_ordered; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_perf_release; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_cpu_perf_grant; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_req_ready; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_req_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [26:0] dcache_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pf; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [43:0] dcache_io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [1:0] dcache_io_ptw_resp_bits_level; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire [3:0] dcache_io_ptw_ptbr_mode; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_status_mxr; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  dcache_io_ptw_status_sum; // @[src/main/scala/rocket/HellaCache.scala 269:43]
  wire  frontend_clock; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_reset; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_auto_icache_master_out_a_ready; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_auto_icache_master_out_a_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [31:0] frontend_auto_icache_master_out_a_bits_address; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_auto_icache_master_out_d_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_size; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [63:0] frontend_auto_icache_master_out_d_bits_data; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_auto_icache_master_out_d_bits_corrupt; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_might_request; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_req_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [39:0] frontend_io_cpu_req_bits_pc; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_req_bits_speculative; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_sfence_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_sfence_bits_rs1; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_sfence_bits_rs2; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [38:0] frontend_io_cpu_sfence_bits_addr; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_resp_ready; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_resp_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [39:0] frontend_io_cpu_resp_bits_pc; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [31:0] frontend_io_cpu_resp_bits_data; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_resp_bits_replay; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_btb_update_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_bht_update_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_flush_icache; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [39:0] frontend_io_cpu_npc; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_cpu_progress; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_req_ready; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_req_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_req_bits_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [26:0] frontend_io_ptw_req_bits_bits_addr; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_valid; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_ae_ptw; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_ae_final; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pf; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [43:0] frontend_io_ptw_resp_bits_pte_ppn; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_d; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_a; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_g; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_u; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_x; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_w; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_r; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_pte_v; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [1:0] frontend_io_ptw_resp_bits_level; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  frontend_io_ptw_resp_bits_homogeneous; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [3:0] frontend_io_ptw_ptbr_mode; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire [1:0] frontend_io_ptw_status_prv; // @[src/main/scala/rocket/Frontend.scala 386:28]
  wire  widget_1_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_in_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_in_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_1_auto_in_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_in_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_1_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_1_auto_in_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_1_auto_in_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_out_a_ready; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_out_a_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [31:0] widget_1_auto_out_a_bits_address; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_out_d_valid; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_1_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [2:0] widget_1_auto_out_d_bits_size; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire [63:0] widget_1_auto_out_d_bits_data; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_1_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  fragmenter_clock; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  fragmenter_reset; // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
  wire  widget_2_clock; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  widget_2_reset; // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_b_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_b_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_b_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_b_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_c_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_c_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_c_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_c_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_c_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_e_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_e_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_e_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_b_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_b_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_b_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_b_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_c_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_c_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_c_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_c_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_c_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_e_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_e_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_e_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  dcacheArb_clock; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_reset; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_req_ready; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_req_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [39:0] dcacheArb_io_requestor_0_req_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_s1_kill; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_s2_nack; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_requestor_0_resp_bits_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_req_ready; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_req_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [39:0] dcacheArb_io_requestor_1_req_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [1:0] dcacheArb_io_requestor_1_req_bits_size; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_req_bits_signed; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [1:0] dcacheArb_io_requestor_1_req_bits_dprv; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s1_kill; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_requestor_1_s1_data_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_nack; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_resp_bits_replay; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_resp_bits_has_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_replay_next; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_ordered; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_perf_release; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_requestor_1_perf_grant; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_req_ready; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_req_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [39:0] dcacheArb_io_mem_req_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [6:0] dcacheArb_io_mem_req_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [4:0] dcacheArb_io_mem_req_bits_cmd; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [1:0] dcacheArb_io_mem_req_bits_size; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_req_bits_signed; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [1:0] dcacheArb_io_mem_req_bits_dprv; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_req_bits_phys; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s1_kill; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_mem_s1_data_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_nack; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [6:0] dcacheArb_io_mem_resp_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_resp_bits_replay; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_resp_bits_has_data; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data_word_bypass; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_replay_next; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_st; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_ordered; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_perf_release; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  dcacheArb_io_mem_perf_grant; // @[src/main/scala/rocket/HellaCache.scala 286:25]
  wire  ptw_clock; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_reset; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_req_ready; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_req_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [26:0] ptw_io_requestor_0_req_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_req_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_ae_ptw; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_ae_final; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pf; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [43:0] ptw_io_requestor_0_resp_bits_pte_ppn; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_d; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_a; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_g; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_u; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_x; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_w; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_r; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_pte_v; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [1:0] ptw_io_requestor_0_resp_bits_level; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_resp_bits_homogeneous; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [3:0] ptw_io_requestor_0_ptbr_mode; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_status_mxr; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_0_status_sum; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_req_ready; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_req_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_req_bits_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [26:0] ptw_io_requestor_1_req_bits_bits_addr; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_req_bits_bits_need_gpa; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_ae_ptw; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_ae_final; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pf; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [43:0] ptw_io_requestor_1_resp_bits_pte_ppn; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_d; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_a; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_g; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_u; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_x; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_w; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_r; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_pte_v; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [1:0] ptw_io_requestor_1_resp_bits_level; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_requestor_1_resp_bits_homogeneous; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [3:0] ptw_io_requestor_1_ptbr_mode; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [1:0] ptw_io_requestor_1_status_prv; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_req_ready; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_req_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [39:0] ptw_io_mem_req_bits_addr; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_s1_kill; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_s2_nack; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_resp_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [63:0] ptw_io_mem_resp_bits_data; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_mem_s2_xcpt_ae_ld; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [3:0] ptw_io_dpath_ptbr_mode; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [43:0] ptw_io_dpath_ptbr_ppn; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_sfence_valid; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_sfence_bits_rs1; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire [1:0] ptw_io_dpath_status_prv; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_status_mxr; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_status_sum; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_perf_l2hit; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_perf_pte_miss; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  ptw_io_dpath_perf_pte_hit; // @[src/main/scala/rocket/PTW.scala 805:19]
  wire  core_clock; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_reset; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_hartid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_might_request; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_req_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [39:0] core_io_imem_req_bits_pc; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_req_bits_speculative; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_sfence_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_sfence_bits_rs1; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_sfence_bits_rs2; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [38:0] core_io_imem_sfence_bits_addr; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_resp_ready; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_resp_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [39:0] core_io_imem_resp_bits_pc; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [31:0] core_io_imem_resp_bits_data; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_resp_bits_xcpt_pf_inst; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_resp_bits_xcpt_ae_inst; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_resp_bits_replay; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_btb_update_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_bht_update_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_flush_icache; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_imem_progress; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_req_ready; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_req_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [39:0] core_io_dmem_req_bits_addr; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [6:0] core_io_dmem_req_bits_tag; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [4:0] core_io_dmem_req_bits_cmd; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [1:0] core_io_dmem_req_bits_size; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_req_bits_signed; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [1:0] core_io_dmem_req_bits_dprv; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_req_bits_dv; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s1_kill; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [63:0] core_io_dmem_s1_data_data; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_nack; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_resp_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [6:0] core_io_dmem_resp_bits_tag; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [63:0] core_io_dmem_resp_bits_data; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_resp_bits_replay; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_resp_bits_has_data; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_replay_next; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_ma_ld; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_ma_st; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_pf_ld; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_pf_st; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_ae_ld; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_s2_xcpt_ae_st; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_ordered; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_perf_release; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_dmem_perf_grant; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [3:0] core_io_ptw_ptbr_mode; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [43:0] core_io_ptw_ptbr_ppn; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_ptw_sfence_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_ptw_sfence_bits_rs1; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire [1:0] core_io_ptw_status_prv; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_ptw_status_mxr; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_ptw_status_sum; // @[src/main/scala/tile/RocketTile.scala 127:20]
  wire  core_io_rocc_cmd_valid; // @[src/main/scala/tile/RocketTile.scala 127:20]
  TLXbar_8 tlMasterXbar ( // @[src/main/scala/tile/BaseTile.scala 224:42]
    .clock(tlMasterXbar_clock),
    .reset(tlMasterXbar_reset),
    .auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
    .auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tlMasterXbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
    .auto_in_0_b_ready(tlMasterXbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(tlMasterXbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_param(tlMasterXbar_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tlMasterXbar_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tlMasterXbar_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tlMasterXbar_auto_in_0_b_bits_address),
    .auto_in_0_c_ready(tlMasterXbar_auto_in_0_c_ready),
    .auto_in_0_c_valid(tlMasterXbar_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tlMasterXbar_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tlMasterXbar_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tlMasterXbar_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tlMasterXbar_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tlMasterXbar_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tlMasterXbar_auto_in_0_c_bits_data),
    .auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tlMasterXbar_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tlMasterXbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tlMasterXbar_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
    .auto_in_0_e_ready(tlMasterXbar_auto_in_0_e_ready),
    .auto_in_0_e_valid(tlMasterXbar_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tlMasterXbar_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
    .auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
    .auto_out_b_ready(tlMasterXbar_auto_out_b_ready),
    .auto_out_b_valid(tlMasterXbar_auto_out_b_valid),
    .auto_out_b_bits_param(tlMasterXbar_auto_out_b_bits_param),
    .auto_out_b_bits_size(tlMasterXbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(tlMasterXbar_auto_out_b_bits_address),
    .auto_out_c_ready(tlMasterXbar_auto_out_c_ready),
    .auto_out_c_valid(tlMasterXbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(tlMasterXbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tlMasterXbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(tlMasterXbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(tlMasterXbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(tlMasterXbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(tlMasterXbar_auto_out_c_bits_data),
    .auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
    .auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt),
    .auto_out_e_ready(tlMasterXbar_auto_out_e_ready),
    .auto_out_e_valid(tlMasterXbar_auto_out_e_valid),
    .auto_out_e_bits_sink(tlMasterXbar_auto_out_e_bits_sink)
  );
  TLXbar_9 tlSlaveXbar ( // @[src/main/scala/tile/BaseTile.scala 225:41]
    .clock(tlSlaveXbar_clock),
    .reset(tlSlaveXbar_reset)
  );
  IntXbar_1 intXbar ( // @[src/main/scala/tile/BaseTile.scala 226:37]
    .clock(intXbar_clock),
    .reset(intXbar_reset)
  );
  BundleBridgeNexus_6 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset),
    .auto_in(broadcast_auto_in),
    .auto_out(broadcast_auto_out)
  );
  BundleBridgeNexus_7 broadcast_1 ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_1_clock),
    .reset(broadcast_1_reset)
  );
  BundleBridgeNexus_8 broadcast_2 ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_2_clock),
    .reset(broadcast_2_reset)
  );
  BundleBridgeNexus_9 nexus ( // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
    .clock(nexus_clock),
    .reset(nexus_reset)
  );
  BundleBridgeNexus_10 broadcast_3 ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_3_clock),
    .reset(broadcast_3_reset)
  );
  BundleBridgeNexus_11 nexus_1 ( // @[src/main/scala/diplomacy/BundleBridge.scala 184:27]
    .clock(nexus_1_clock),
    .reset(nexus_1_reset)
  );
  BundleBridgeNexus_12 broadcast_4 ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_4_clock),
    .reset(broadcast_4_reset)
  );
  TLWidthWidget_7 widget ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(widget_auto_in_a_bits_param),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_b_ready(widget_auto_in_b_ready),
    .auto_in_b_valid(widget_auto_in_b_valid),
    .auto_in_b_bits_param(widget_auto_in_b_bits_param),
    .auto_in_b_bits_size(widget_auto_in_b_bits_size),
    .auto_in_b_bits_source(widget_auto_in_b_bits_source),
    .auto_in_b_bits_address(widget_auto_in_b_bits_address),
    .auto_in_c_ready(widget_auto_in_c_ready),
    .auto_in_c_valid(widget_auto_in_c_valid),
    .auto_in_c_bits_opcode(widget_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(widget_auto_in_c_bits_param),
    .auto_in_c_bits_size(widget_auto_in_c_bits_size),
    .auto_in_c_bits_source(widget_auto_in_c_bits_source),
    .auto_in_c_bits_address(widget_auto_in_c_bits_address),
    .auto_in_c_bits_data(widget_auto_in_c_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(widget_auto_in_d_bits_param),
    .auto_in_d_bits_size(widget_auto_in_d_bits_size),
    .auto_in_d_bits_source(widget_auto_in_d_bits_source),
    .auto_in_d_bits_sink(widget_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(widget_auto_in_d_bits_denied),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_in_e_ready(widget_auto_in_e_ready),
    .auto_in_e_valid(widget_auto_in_e_valid),
    .auto_in_e_bits_sink(widget_auto_in_e_bits_sink),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(widget_auto_out_a_bits_param),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_b_ready(widget_auto_out_b_ready),
    .auto_out_b_valid(widget_auto_out_b_valid),
    .auto_out_b_bits_param(widget_auto_out_b_bits_param),
    .auto_out_b_bits_size(widget_auto_out_b_bits_size),
    .auto_out_b_bits_source(widget_auto_out_b_bits_source),
    .auto_out_b_bits_address(widget_auto_out_b_bits_address),
    .auto_out_c_ready(widget_auto_out_c_ready),
    .auto_out_c_valid(widget_auto_out_c_valid),
    .auto_out_c_bits_opcode(widget_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(widget_auto_out_c_bits_param),
    .auto_out_c_bits_size(widget_auto_out_c_bits_size),
    .auto_out_c_bits_source(widget_auto_out_c_bits_source),
    .auto_out_c_bits_address(widget_auto_out_c_bits_address),
    .auto_out_c_bits_data(widget_auto_out_c_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(widget_auto_out_d_bits_param),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_sink(widget_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(widget_auto_out_d_bits_denied),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data),
    .auto_out_e_ready(widget_auto_out_e_ready),
    .auto_out_e_valid(widget_auto_out_e_valid),
    .auto_out_e_bits_sink(widget_auto_out_e_bits_sink)
  );
  DCache dcache ( // @[src/main/scala/rocket/HellaCache.scala 269:43]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_size(dcache_io_cpu_req_bits_size),
    .io_cpu_req_bits_signed(dcache_io_cpu_req_bits_signed),
    .io_cpu_req_bits_dprv(dcache_io_cpu_req_bits_dprv),
    .io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s1_data_mask(dcache_io_cpu_s1_data_mask),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(dcache_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(dcache_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_size(dcache_io_cpu_resp_bits_size),
    .io_cpu_resp_bits_signed(dcache_io_cpu_resp_bits_signed),
    .io_cpu_resp_bits_dprv(dcache_io_cpu_resp_bits_dprv),
    .io_cpu_resp_bits_dv(dcache_io_cpu_resp_bits_dv),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_mask(dcache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_data_raw(dcache_io_cpu_resp_bits_data_raw),
    .io_cpu_resp_bits_store_data(dcache_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(dcache_io_cpu_replay_next),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_gf_ld(dcache_io_cpu_s2_xcpt_gf_ld),
    .io_cpu_s2_xcpt_gf_st(dcache_io_cpu_s2_xcpt_gf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_cpu_perf_release(dcache_io_cpu_perf_release),
    .io_cpu_perf_grant(dcache_io_cpu_perf_grant),
    .io_ptw_req_ready(dcache_io_ptw_req_ready),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(dcache_io_ptw_req_bits_bits_addr),
    .io_ptw_req_bits_bits_need_gpa(dcache_io_ptw_req_bits_bits_need_gpa),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_ptw(dcache_io_ptw_resp_bits_ae_ptw),
    .io_ptw_resp_bits_ae_final(dcache_io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pf(dcache_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum)
  );
  Frontend frontend ( // @[src/main/scala/rocket/Frontend.scala 386:28]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
    .io_cpu_might_request(frontend_io_cpu_might_request),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),
    .io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_cpu_progress(frontend_io_cpu_progress),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),
    .io_ptw_req_bits_bits_need_gpa(frontend_io_ptw_req_bits_bits_need_gpa),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_ptw(frontend_io_ptw_resp_bits_ae_ptw),
    .io_ptw_resp_bits_ae_final(frontend_io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pf(frontend_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_status_prv(frontend_io_ptw_status_prv)
  );
  TLWidthWidget_8 widget_1 ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_1_clock),
    .reset(widget_1_reset),
    .auto_in_a_ready(widget_1_auto_in_a_ready),
    .auto_in_a_valid(widget_1_auto_in_a_valid),
    .auto_in_a_bits_address(widget_1_auto_in_a_bits_address),
    .auto_in_d_valid(widget_1_auto_in_d_valid),
    .auto_in_d_bits_opcode(widget_1_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(widget_1_auto_in_d_bits_size),
    .auto_in_d_bits_data(widget_1_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(widget_1_auto_in_d_bits_corrupt),
    .auto_out_a_ready(widget_1_auto_out_a_ready),
    .auto_out_a_valid(widget_1_auto_out_a_valid),
    .auto_out_a_bits_address(widget_1_auto_out_a_bits_address),
    .auto_out_d_valid(widget_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(widget_1_auto_out_d_bits_size),
    .auto_out_d_bits_data(widget_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(widget_1_auto_out_d_bits_corrupt)
  );
  TLFragmenter_1 fragmenter ( // @[src/main/scala/tilelink/Fragmenter.scala 335:34]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset)
  );
  TLWidthWidget_9 widget_2 ( // @[src/main/scala/tilelink/WidthWidget.scala 220:28]
    .clock(widget_2_clock),
    .reset(widget_2_reset)
  );
  TLBuffer_6 buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_b_ready(buffer_auto_in_b_ready),
    .auto_in_b_valid(buffer_auto_in_b_valid),
    .auto_in_b_bits_param(buffer_auto_in_b_bits_param),
    .auto_in_b_bits_size(buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(buffer_auto_in_b_bits_address),
    .auto_in_c_ready(buffer_auto_in_c_ready),
    .auto_in_c_valid(buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(buffer_auto_in_c_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_in_e_ready(buffer_auto_in_e_ready),
    .auto_in_e_valid(buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_b_ready(buffer_auto_out_b_ready),
    .auto_out_b_valid(buffer_auto_out_b_valid),
    .auto_out_b_bits_param(buffer_auto_out_b_bits_param),
    .auto_out_b_bits_size(buffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(buffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(buffer_auto_out_b_bits_address),
    .auto_out_c_ready(buffer_auto_out_c_ready),
    .auto_out_c_valid(buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(buffer_auto_out_c_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .auto_out_e_ready(buffer_auto_out_e_ready),
    .auto_out_e_valid(buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(buffer_auto_out_e_bits_sink)
  );
  TLBuffer_7 buffer_1 ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset)
  );
  HellaCacheArbiter dcacheArb ( // @[src/main/scala/rocket/HellaCache.scala 286:25]
    .clock(dcacheArb_clock),
    .reset(dcacheArb_reset),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_size(dcacheArb_io_requestor_1_req_bits_size),
    .io_requestor_1_req_bits_signed(dcacheArb_io_requestor_1_req_bits_signed),
    .io_requestor_1_req_bits_dprv(dcacheArb_io_requestor_1_req_bits_dprv),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
    .io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_requestor_1_perf_release(dcacheArb_io_requestor_1_perf_release),
    .io_requestor_1_perf_grant(dcacheArb_io_requestor_1_perf_grant),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_size(dcacheArb_io_mem_req_bits_size),
    .io_mem_req_bits_signed(dcacheArb_io_mem_req_bits_signed),
    .io_mem_req_bits_dprv(dcacheArb_io_mem_req_bits_dprv),
    .io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_replay_next(dcacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(dcacheArb_io_mem_ordered),
    .io_mem_perf_release(dcacheArb_io_mem_perf_release),
    .io_mem_perf_grant(dcacheArb_io_mem_perf_grant)
  );
  PTW ptw ( // @[src/main/scala/rocket/PTW.scala 805:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),
    .io_requestor_0_req_bits_bits_need_gpa(ptw_io_requestor_0_req_bits_bits_need_gpa),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae_ptw(ptw_io_requestor_0_resp_bits_ae_ptw),
    .io_requestor_0_resp_bits_ae_final(ptw_io_requestor_0_resp_bits_ae_final),
    .io_requestor_0_resp_bits_pf(ptw_io_requestor_0_resp_bits_pf),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),
    .io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),
    .io_requestor_1_req_bits_bits_need_gpa(ptw_io_requestor_1_req_bits_bits_need_gpa),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae_ptw(ptw_io_requestor_1_resp_bits_ae_ptw),
    .io_requestor_1_resp_bits_ae_final(ptw_io_requestor_1_resp_bits_ae_final),
    .io_requestor_1_resp_bits_pf(ptw_io_requestor_1_resp_bits_pf),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_perf_l2hit(ptw_io_dpath_perf_l2hit),
    .io_dpath_perf_pte_miss(ptw_io_dpath_perf_pte_miss),
    .io_dpath_perf_pte_hit(ptw_io_dpath_perf_pte_hit)
  );
  Rocket core ( // @[src/main/scala/tile/RocketTile.scala 127:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_imem_might_request(core_io_imem_might_request),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),
    .io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_progress(core_io_imem_progress),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_size(core_io_dmem_req_bits_size),
    .io_dmem_req_bits_signed(core_io_dmem_req_bits_signed),
    .io_dmem_req_bits_dprv(core_io_dmem_req_bits_dprv),
    .io_dmem_req_bits_dv(core_io_dmem_req_bits_dv),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
    .io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_dmem_perf_release(core_io_dmem_perf_release),
    .io_dmem_perf_grant(core_io_dmem_perf_grant),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid)
  );
  assign auto_buffer_out_a_valid = buffer_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_param = buffer_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_size = buffer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_source = buffer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_address = buffer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_mask = buffer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_a_bits_data = buffer_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_b_ready = buffer_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_valid = buffer_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_opcode = buffer_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_param = buffer_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_size = buffer_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_source = buffer_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_address = buffer_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_c_bits_data = buffer_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_d_ready = buffer_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_e_valid = buffer_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_buffer_out_e_bits_sink = buffer_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tlMasterXbar_clock = clock;
  assign tlMasterXbar_reset = reset;
  assign tlMasterXbar_auto_in_1_a_valid = widget_1_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_1_a_bits_address = widget_1_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_valid = widget_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_param = widget_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_size = widget_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_source = widget_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_address = widget_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_mask = widget_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_a_bits_data = widget_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_b_ready = widget_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_valid = widget_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_opcode = widget_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_param = widget_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_size = widget_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_source = widget_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_address = widget_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_c_bits_data = widget_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_d_ready = widget_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_e_valid = widget_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_in_0_e_bits_sink = widget_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tlMasterXbar_auto_out_a_ready = buffer_auto_in_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_b_valid = buffer_auto_in_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_b_bits_param = buffer_auto_in_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_b_bits_size = buffer_auto_in_b_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_b_bits_source = buffer_auto_in_b_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_b_bits_address = buffer_auto_in_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_c_ready = buffer_auto_in_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_valid = buffer_auto_in_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlMasterXbar_auto_out_e_ready = buffer_auto_in_e_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tlSlaveXbar_clock = clock;
  assign tlSlaveXbar_reset = reset;
  assign intXbar_clock = clock;
  assign intXbar_reset = reset;
  assign broadcast_clock = clock;
  assign broadcast_reset = reset;
  assign broadcast_auto_in = auto_hartid_in; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign broadcast_1_clock = clock;
  assign broadcast_1_reset = reset;
  assign broadcast_2_clock = clock;
  assign broadcast_2_reset = reset;
  assign nexus_clock = clock;
  assign nexus_reset = reset;
  assign broadcast_3_clock = clock;
  assign broadcast_3_reset = reset;
  assign nexus_1_clock = clock;
  assign nexus_1_reset = reset;
  assign broadcast_4_clock = clock;
  assign broadcast_4_reset = reset;
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = dcache_auto_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_opcode = dcache_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_param = dcache_auto_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_size = dcache_auto_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_source = dcache_auto_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_address = dcache_auto_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_mask = dcache_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_a_bits_data = dcache_auto_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_b_ready = dcache_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_valid = dcache_auto_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_param = dcache_auto_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_size = dcache_auto_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_source = dcache_auto_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_address = dcache_auto_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_c_bits_data = dcache_auto_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_d_ready = dcache_auto_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_e_valid = dcache_auto_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_in_e_bits_sink = dcache_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = widget_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_b_valid = widget_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_b_bits_param = widget_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_b_bits_size = widget_auto_in_b_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_b_bits_source = widget_auto_in_b_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_b_bits_address = widget_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_c_ready = widget_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_valid = widget_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_param = widget_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_size = widget_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_source = widget_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_sink = widget_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_denied = widget_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_auto_out_e_ready = widget_auto_in_e_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_size = dcacheArb_io_mem_req_bits_size; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_signed = dcacheArb_io_mem_req_bits_signed; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_dprv = dcacheArb_io_mem_req_bits_dprv; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_req_bits_phys = dcacheArb_io_mem_req_bits_phys; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_cpu_s1_data_mask = 8'h0; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcache_io_ptw_req_ready = ptw_io_requestor_0_req_ready; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_ae_ptw = ptw_io_requestor_0_resp_bits_ae_ptw; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_ae_final = ptw_io_requestor_0_resp_bits_ae_final; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pf = ptw_io_requestor_0_resp_bits_pf; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = widget_1_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_auto_icache_master_out_d_valid = widget_1_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_auto_icache_master_out_d_bits_opcode = widget_1_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_auto_icache_master_out_d_bits_size = widget_1_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_auto_icache_master_out_d_bits_data = widget_1_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_auto_icache_master_out_d_bits_corrupt = widget_1_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign frontend_io_cpu_might_request = core_io_imem_might_request; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_sfence_valid = core_io_imem_sfence_valid; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_sfence_bits_addr = core_io_imem_sfence_bits_addr; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_btb_update_valid = core_io_imem_btb_update_valid; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_bht_update_valid = core_io_imem_bht_update_valid; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_cpu_progress = core_io_imem_progress; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_ae_ptw = ptw_io_requestor_1_resp_bits_ae_ptw; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_ae_final = ptw_io_requestor_1_resp_bits_ae_final; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pf = ptw_io_requestor_1_resp_bits_pf; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign widget_1_clock = clock;
  assign widget_1_reset = reset;
  assign widget_1_auto_in_a_valid = frontend_auto_icache_master_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign widget_1_auto_in_a_bits_address = frontend_auto_icache_master_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign widget_1_auto_out_a_ready = tlMasterXbar_auto_in_1_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_1_auto_out_d_valid = tlMasterXbar_auto_in_1_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_1_auto_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_1_auto_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_1_auto_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign widget_1_auto_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign fragmenter_clock = clock;
  assign fragmenter_reset = reset;
  assign widget_2_clock = clock;
  assign widget_2_reset = reset;
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_a_valid = tlMasterXbar_auto_out_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_b_ready = tlMasterXbar_auto_out_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_valid = tlMasterXbar_auto_out_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_param = tlMasterXbar_auto_out_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_size = tlMasterXbar_auto_out_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_source = tlMasterXbar_auto_out_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_address = tlMasterXbar_auto_out_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_c_bits_data = tlMasterXbar_auto_out_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_d_ready = tlMasterXbar_auto_out_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_e_valid = tlMasterXbar_auto_out_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_in_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign buffer_auto_out_a_ready = auto_buffer_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_valid = auto_buffer_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_param = auto_buffer_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_size = auto_buffer_out_b_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_source = auto_buffer_out_b_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_address = auto_buffer_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_c_ready = auto_buffer_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_valid = auto_buffer_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_opcode = auto_buffer_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_param = auto_buffer_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_size = auto_buffer_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_source = auto_buffer_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_sink = auto_buffer_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_denied = auto_buffer_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_data = auto_buffer_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_corrupt = auto_buffer_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_e_ready = auto_buffer_out_e_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign dcacheArb_clock = clock;
  assign dcacheArb_reset = reset;
  assign dcacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_size = core_io_dmem_req_bits_size; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_signed = core_io_dmem_req_bits_signed; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_req_bits_dprv = core_io_dmem_req_bits_dprv; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_perf_release = dcache_io_cpu_perf_release; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign dcacheArb_io_mem_perf_grant = dcache_io_cpu_perf_grant; // @[src/main/scala/rocket/HellaCache.scala 287:30]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_0_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_0_req_bits_bits_need_gpa = dcache_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_1_req_bits_valid = frontend_io_ptw_req_bits_valid; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_1_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_requestor_1_req_bits_bits_need_gpa = frontend_io_ptw_req_bits_bits_need_gpa; // @[src/main/scala/tile/RocketTile.scala 211:20]
  assign ptw_io_mem_req_ready = dcacheArb_io_requestor_0_req_ready; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign ptw_io_mem_s2_nack = dcacheArb_io_requestor_0_s2_nack; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign ptw_io_mem_resp_valid = dcacheArb_io_requestor_0_resp_valid; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign ptw_io_mem_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign ptw_io_mem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum; // @[src/main/scala/tile/RocketTile.scala 173:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = broadcast_auto_out; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay; // @[src/main/scala/tile/RocketTile.scala 163:32]
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_1_resp_bits_replay; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_replay_next = dcacheArb_io_requestor_1_replay_next; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_perf_release = dcacheArb_io_requestor_1_perf_release; // @[src/main/scala/tile/RocketTile.scala 210:26]
  assign core_io_dmem_perf_grant = dcacheArb_io_requestor_1_perf_grant; // @[src/main/scala/tile/RocketTile.scala 210:26]
endmodule
module TileResetDomain(
  input         auto_tile_buffer_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tile_buffer_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tile_buffer_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tile_buffer_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_tile_buffer_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tile_buffer_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tile_buffer_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tile_buffer_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tile_buffer_out_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tile_buffer_out_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tile_buffer_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tile_buffer_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tile_buffer_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tile_buffer_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tile_buffer_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tile_buffer_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tile_buffer_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tile_buffer_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tile_buffer_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tile_buffer_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tile_buffer_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tile_buffer_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tile_buffer_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_buffer_out_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tile_buffer_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tile_buffer_out_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tile_hartid_in, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_clock_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_clock_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  tile_clock; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_reset; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_a_ready; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_a_valid; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_a_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_a_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_a_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_a_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [31:0] tile_auto_buffer_out_a_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [7:0] tile_auto_buffer_out_a_bits_mask; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [63:0] tile_auto_buffer_out_a_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_b_ready; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_b_valid; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_b_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_b_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_b_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [31:0] tile_auto_buffer_out_b_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_c_ready; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_c_valid; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_c_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_c_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_c_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_c_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [31:0] tile_auto_buffer_out_c_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [63:0] tile_auto_buffer_out_c_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_d_ready; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_d_valid; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_d_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_d_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [2:0] tile_auto_buffer_out_d_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_d_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_d_bits_sink; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_d_bits_denied; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [63:0] tile_auto_buffer_out_d_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_d_bits_corrupt; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_e_ready; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_buffer_out_e_valid; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire [1:0] tile_auto_buffer_out_e_bits_sink; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  wire  tile_auto_hartid_in; // @[src/main/scala/subsystem/HasTiles.scala 251:53]
  RocketTile tile ( // @[src/main/scala/subsystem/HasTiles.scala 251:53]
    .clock(tile_clock),
    .reset(tile_reset),
    .auto_buffer_out_a_ready(tile_auto_buffer_out_a_ready),
    .auto_buffer_out_a_valid(tile_auto_buffer_out_a_valid),
    .auto_buffer_out_a_bits_opcode(tile_auto_buffer_out_a_bits_opcode),
    .auto_buffer_out_a_bits_param(tile_auto_buffer_out_a_bits_param),
    .auto_buffer_out_a_bits_size(tile_auto_buffer_out_a_bits_size),
    .auto_buffer_out_a_bits_source(tile_auto_buffer_out_a_bits_source),
    .auto_buffer_out_a_bits_address(tile_auto_buffer_out_a_bits_address),
    .auto_buffer_out_a_bits_mask(tile_auto_buffer_out_a_bits_mask),
    .auto_buffer_out_a_bits_data(tile_auto_buffer_out_a_bits_data),
    .auto_buffer_out_b_ready(tile_auto_buffer_out_b_ready),
    .auto_buffer_out_b_valid(tile_auto_buffer_out_b_valid),
    .auto_buffer_out_b_bits_param(tile_auto_buffer_out_b_bits_param),
    .auto_buffer_out_b_bits_size(tile_auto_buffer_out_b_bits_size),
    .auto_buffer_out_b_bits_source(tile_auto_buffer_out_b_bits_source),
    .auto_buffer_out_b_bits_address(tile_auto_buffer_out_b_bits_address),
    .auto_buffer_out_c_ready(tile_auto_buffer_out_c_ready),
    .auto_buffer_out_c_valid(tile_auto_buffer_out_c_valid),
    .auto_buffer_out_c_bits_opcode(tile_auto_buffer_out_c_bits_opcode),
    .auto_buffer_out_c_bits_param(tile_auto_buffer_out_c_bits_param),
    .auto_buffer_out_c_bits_size(tile_auto_buffer_out_c_bits_size),
    .auto_buffer_out_c_bits_source(tile_auto_buffer_out_c_bits_source),
    .auto_buffer_out_c_bits_address(tile_auto_buffer_out_c_bits_address),
    .auto_buffer_out_c_bits_data(tile_auto_buffer_out_c_bits_data),
    .auto_buffer_out_d_ready(tile_auto_buffer_out_d_ready),
    .auto_buffer_out_d_valid(tile_auto_buffer_out_d_valid),
    .auto_buffer_out_d_bits_opcode(tile_auto_buffer_out_d_bits_opcode),
    .auto_buffer_out_d_bits_param(tile_auto_buffer_out_d_bits_param),
    .auto_buffer_out_d_bits_size(tile_auto_buffer_out_d_bits_size),
    .auto_buffer_out_d_bits_source(tile_auto_buffer_out_d_bits_source),
    .auto_buffer_out_d_bits_sink(tile_auto_buffer_out_d_bits_sink),
    .auto_buffer_out_d_bits_denied(tile_auto_buffer_out_d_bits_denied),
    .auto_buffer_out_d_bits_data(tile_auto_buffer_out_d_bits_data),
    .auto_buffer_out_d_bits_corrupt(tile_auto_buffer_out_d_bits_corrupt),
    .auto_buffer_out_e_ready(tile_auto_buffer_out_e_ready),
    .auto_buffer_out_e_valid(tile_auto_buffer_out_e_valid),
    .auto_buffer_out_e_bits_sink(tile_auto_buffer_out_e_bits_sink),
    .auto_hartid_in(tile_auto_hartid_in)
  );
  assign auto_tile_buffer_out_a_valid = tile_auto_buffer_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_opcode = tile_auto_buffer_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_param = tile_auto_buffer_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_size = tile_auto_buffer_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_source = tile_auto_buffer_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_address = tile_auto_buffer_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_mask = tile_auto_buffer_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_a_bits_data = tile_auto_buffer_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_b_ready = tile_auto_buffer_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_valid = tile_auto_buffer_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_opcode = tile_auto_buffer_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_param = tile_auto_buffer_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_size = tile_auto_buffer_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_source = tile_auto_buffer_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_address = tile_auto_buffer_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_c_bits_data = tile_auto_buffer_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_d_ready = tile_auto_buffer_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_e_valid = tile_auto_buffer_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_tile_buffer_out_e_bits_sink = tile_auto_buffer_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tile_clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tile_reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tile_auto_buffer_out_a_ready = auto_tile_buffer_out_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_b_valid = auto_tile_buffer_out_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_b_bits_param = auto_tile_buffer_out_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_b_bits_size = auto_tile_buffer_out_b_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_b_bits_source = auto_tile_buffer_out_b_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_b_bits_address = auto_tile_buffer_out_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_c_ready = auto_tile_buffer_out_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_valid = auto_tile_buffer_out_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_opcode = auto_tile_buffer_out_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_param = auto_tile_buffer_out_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_size = auto_tile_buffer_out_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_source = auto_tile_buffer_out_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_sink = auto_tile_buffer_out_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_denied = auto_tile_buffer_out_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_data = auto_tile_buffer_out_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_d_bits_corrupt = auto_tile_buffer_out_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_buffer_out_e_ready = auto_tile_buffer_out_e_ready; // @[src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign tile_auto_hartid_in = auto_tile_hartid_in; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module FixedClockBroadcast_6(
  input   auto_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input   auto_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output  auto_out_reset // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  assign auto_out_clock = auto_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_reset = auto_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module Queue_40(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_mask, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_param [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_address [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_mask [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_mask_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1239_clock;
  wire  line_1239_reset;
  wire  line_1239_valid;
  reg  line_1239_valid_reg;
  wire  line_1240_clock;
  wire  line_1240_reset;
  wire  line_1240_valid;
  reg  line_1240_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1241_clock;
  wire  line_1241_reset;
  wire  line_1241_valid;
  reg  line_1241_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1239)) line_1239 (
    .clock(line_1239_clock),
    .reset(line_1239_reset),
    .valid(line_1239_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1240)) line_1240 (
    .clock(line_1240_clock),
    .reset(line_1240_reset),
    .valid(line_1240_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1241)) line_1241 (
    .clock(line_1241_clock),
    .reset(line_1241_reset),
    .valid(line_1241_valid)
  );
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = enq_ptr_value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_en = 1'h1;
  assign ram_mask_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = enq_ptr_value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1239_clock = clock;
  assign line_1239_reset = reset;
  assign line_1239_valid = do_enq ^ line_1239_valid_reg;
  assign line_1240_clock = clock;
  assign line_1240_reset = reset;
  assign line_1240_valid = do_deq ^ line_1240_valid_reg;
  assign line_1241_clock = clock;
  assign line_1241_reset = reset;
  assign line_1241_valid = _T ^ line_1241_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1239_valid_reg <= do_enq;
    line_1240_valid_reg <= do_deq;
    line_1241_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  deq_ptr_value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1239_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1240_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1241_valid_reg = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_41(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_sink, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_denied, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_corrupt, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_sink, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_denied, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_corrupt // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_param [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_sink [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_denied [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_denied_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_corrupt [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_corrupt_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1242_clock;
  wire  line_1242_reset;
  wire  line_1242_valid;
  reg  line_1242_valid_reg;
  wire  line_1243_clock;
  wire  line_1243_reset;
  wire  line_1243_valid;
  reg  line_1243_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1244_clock;
  wire  line_1244_reset;
  wire  line_1244_valid;
  reg  line_1244_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1242)) line_1242 (
    .clock(line_1242_clock),
    .reset(line_1242_reset),
    .valid(line_1242_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1243)) line_1243 (
    .clock(line_1243_clock),
    .reset(line_1243_reset),
    .valid(line_1243_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1244)) line_1244 (
    .clock(line_1244_clock),
    .reset(line_1244_reset),
    .valid(line_1244_valid)
  );
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = enq_ptr_value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sink_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = enq_ptr_value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_en = 1'h1;
  assign ram_denied_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = enq_ptr_value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_en = 1'h1;
  assign ram_corrupt_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = enq_ptr_value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1242_clock = clock;
  assign line_1242_reset = reset;
  assign line_1242_valid = do_enq ^ line_1242_valid_reg;
  assign line_1243_clock = clock;
  assign line_1243_reset = reset;
  assign line_1243_valid = do_deq ^ line_1243_valid_reg;
  assign line_1244_clock = clock;
  assign line_1244_reset = reset;
  assign line_1244_valid = _T ^ line_1244_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1242_valid_reg <= do_enq;
    line_1243_valid_reg <= do_deq;
    line_1244_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enq_ptr_value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  deq_ptr_value = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1242_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1243_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1244_valid_reg = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_42(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_address // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_param [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_address [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1245_clock;
  wire  line_1245_reset;
  wire  line_1245_valid;
  reg  line_1245_valid_reg;
  wire  line_1246_clock;
  wire  line_1246_reset;
  wire  line_1246_valid;
  reg  line_1246_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1247_clock;
  wire  line_1247_reset;
  wire  line_1247_valid;
  reg  line_1247_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1245)) line_1245 (
    .clock(line_1245_clock),
    .reset(line_1245_reset),
    .valid(line_1245_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1246)) line_1246 (
    .clock(line_1246_clock),
    .reset(line_1246_reset),
    .valid(line_1246_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1247)) line_1247 (
    .clock(line_1247_clock),
    .reset(line_1247_reset),
    .valid(line_1247_valid)
  );
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = enq_ptr_value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = 3'h5;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = 2'h0;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1245_clock = clock;
  assign line_1245_reset = reset;
  assign line_1245_valid = do_enq ^ line_1245_valid_reg;
  assign line_1246_clock = clock;
  assign line_1246_reset = reset;
  assign line_1246_valid = do_deq ^ line_1246_valid_reg;
  assign line_1247_clock = clock;
  assign line_1247_reset = reset;
  assign line_1247_valid = _T ^ line_1247_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1245_valid_reg <= do_enq;
    line_1246_valid_reg <= do_deq;
    line_1247_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1245_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1246_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1247_valid_reg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_43(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_opcode, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_param, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_source, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_address, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_opcode_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_param [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_param_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_source [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_source_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_address [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_address_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1248_clock;
  wire  line_1248_reset;
  wire  line_1248_valid;
  reg  line_1248_valid_reg;
  wire  line_1249_clock;
  wire  line_1249_reset;
  wire  line_1249_valid;
  reg  line_1249_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1250_clock;
  wire  line_1250_reset;
  wire  line_1250_valid;
  reg  line_1250_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1248)) line_1248 (
    .clock(line_1248_clock),
    .reset(line_1248_reset),
    .valid(line_1248_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1249)) line_1249 (
    .clock(line_1249_clock),
    .reset(line_1249_reset),
    .valid(line_1249_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1250)) line_1250 (
    .clock(line_1250_clock),
    .reset(line_1250_reset),
    .valid(line_1250_valid)
  );
  assign ram_opcode_io_deq_bits_MPORT_en = 1'h1;
  assign ram_opcode_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = enq_ptr_value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_en = 1'h1;
  assign ram_param_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = enq_ptr_value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = enq_ptr_value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_en = 1'h1;
  assign ram_source_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = enq_ptr_value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_en = 1'h1;
  assign ram_address_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = enq_ptr_value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1248_clock = clock;
  assign line_1248_reset = reset;
  assign line_1248_valid = do_enq ^ line_1248_valid_reg;
  assign line_1249_clock = clock;
  assign line_1249_reset = reset;
  assign line_1249_valid = do_deq ^ line_1249_valid_reg;
  assign line_1250_clock = clock;
  assign line_1250_reset = reset;
  assign line_1250_valid = _T ^ line_1250_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1248_valid_reg <= do_enq;
    line_1249_valid_reg <= do_deq;
    line_1250_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  deq_ptr_value = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  maybe_full = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1248_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1249_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1250_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_44(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0] io_enq_bits_sink, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0] io_deq_bits_sink // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram_sink [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_sink_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1251_clock;
  wire  line_1251_reset;
  wire  line_1251_valid;
  reg  line_1251_valid_reg;
  wire  line_1252_clock;
  wire  line_1252_reset;
  wire  line_1252_valid;
  reg  line_1252_valid_reg;
  wire  _T = do_enq != io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1253_clock;
  wire  line_1253_reset;
  wire  line_1253_valid;
  reg  line_1253_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1251)) line_1251 (
    .clock(line_1251_clock),
    .reset(line_1251_reset),
    .valid(line_1251_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1252)) line_1252 (
    .clock(line_1252_clock),
    .reset(line_1252_reset),
    .valid(line_1252_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1253)) line_1253 (
    .clock(line_1253_clock),
    .reset(line_1253_reset),
    .valid(line_1253_valid)
  );
  assign ram_sink_io_deq_bits_MPORT_en = 1'h1;
  assign ram_sink_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = enq_ptr_value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1251_clock = clock;
  assign line_1251_reset = reset;
  assign line_1251_valid = do_enq ^ line_1251_valid_reg;
  assign line_1252_clock = clock;
  assign line_1252_reset = reset;
  assign line_1252_valid = io_deq_valid ^ line_1252_valid_reg;
  assign line_1253_clock = clock;
  assign line_1253_reset = reset;
  assign line_1253_valid = _T ^ line_1253_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_deq_valid) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != io_deq_valid) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1251_valid_reg <= do_enq;
    line_1252_valid_reg <= io_deq_valid;
    line_1253_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1251_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1252_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1253_valid_reg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_8(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_b_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_in_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_e_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_e_bits_sink // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  nodeOut_a_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_enq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_enq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_a_q_io_enq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_a_q_io_enq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_a_q_io_enq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_a_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_a_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_deq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_deq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_a_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_a_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_a_q_io_deq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_a_q_io_deq_bits_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_a_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_enq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_enq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_enq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_enq_bits_sink; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_bits_denied; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_d_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_enq_bits_corrupt; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_deq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_deq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_d_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_d_q_io_deq_bits_sink; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_bits_denied; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_d_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_d_q_io_deq_bits_corrupt; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_b_q_io_enq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeIn_b_q_io_enq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_b_q_io_deq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeIn_b_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_b_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeIn_b_q_io_deq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_enq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_enq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_c_q_io_enq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_c_q_io_enq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_c_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_c_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_deq_bits_opcode; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_deq_bits_param; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] nodeOut_c_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_c_q_io_deq_bits_source; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_c_q_io_deq_bits_address; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_c_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_e_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_e_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_e_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_e_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_e_q_io_enq_bits_sink; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_e_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeOut_e_q_io_deq_bits_sink; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  Queue_40 nodeOut_a_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_a_q_clock),
    .reset(nodeOut_a_q_reset),
    .io_enq_ready(nodeOut_a_q_io_enq_ready),
    .io_enq_valid(nodeOut_a_q_io_enq_valid),
    .io_enq_bits_opcode(nodeOut_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(nodeOut_a_q_io_enq_bits_param),
    .io_enq_bits_size(nodeOut_a_q_io_enq_bits_size),
    .io_enq_bits_source(nodeOut_a_q_io_enq_bits_source),
    .io_enq_bits_address(nodeOut_a_q_io_enq_bits_address),
    .io_enq_bits_mask(nodeOut_a_q_io_enq_bits_mask),
    .io_enq_bits_data(nodeOut_a_q_io_enq_bits_data),
    .io_deq_ready(nodeOut_a_q_io_deq_ready),
    .io_deq_valid(nodeOut_a_q_io_deq_valid),
    .io_deq_bits_opcode(nodeOut_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(nodeOut_a_q_io_deq_bits_param),
    .io_deq_bits_size(nodeOut_a_q_io_deq_bits_size),
    .io_deq_bits_source(nodeOut_a_q_io_deq_bits_source),
    .io_deq_bits_address(nodeOut_a_q_io_deq_bits_address),
    .io_deq_bits_mask(nodeOut_a_q_io_deq_bits_mask),
    .io_deq_bits_data(nodeOut_a_q_io_deq_bits_data)
  );
  Queue_41 nodeIn_d_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeIn_d_q_clock),
    .reset(nodeIn_d_q_reset),
    .io_enq_ready(nodeIn_d_q_io_enq_ready),
    .io_enq_valid(nodeIn_d_q_io_enq_valid),
    .io_enq_bits_opcode(nodeIn_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(nodeIn_d_q_io_enq_bits_param),
    .io_enq_bits_size(nodeIn_d_q_io_enq_bits_size),
    .io_enq_bits_source(nodeIn_d_q_io_enq_bits_source),
    .io_enq_bits_sink(nodeIn_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(nodeIn_d_q_io_enq_bits_denied),
    .io_enq_bits_data(nodeIn_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(nodeIn_d_q_io_enq_bits_corrupt),
    .io_deq_ready(nodeIn_d_q_io_deq_ready),
    .io_deq_valid(nodeIn_d_q_io_deq_valid),
    .io_deq_bits_opcode(nodeIn_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(nodeIn_d_q_io_deq_bits_param),
    .io_deq_bits_size(nodeIn_d_q_io_deq_bits_size),
    .io_deq_bits_source(nodeIn_d_q_io_deq_bits_source),
    .io_deq_bits_sink(nodeIn_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(nodeIn_d_q_io_deq_bits_denied),
    .io_deq_bits_data(nodeIn_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(nodeIn_d_q_io_deq_bits_corrupt)
  );
  Queue_42 nodeIn_b_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeIn_b_q_clock),
    .reset(nodeIn_b_q_reset),
    .io_enq_ready(nodeIn_b_q_io_enq_ready),
    .io_enq_valid(nodeIn_b_q_io_enq_valid),
    .io_enq_bits_param(nodeIn_b_q_io_enq_bits_param),
    .io_enq_bits_address(nodeIn_b_q_io_enq_bits_address),
    .io_deq_ready(nodeIn_b_q_io_deq_ready),
    .io_deq_valid(nodeIn_b_q_io_deq_valid),
    .io_deq_bits_param(nodeIn_b_q_io_deq_bits_param),
    .io_deq_bits_size(nodeIn_b_q_io_deq_bits_size),
    .io_deq_bits_source(nodeIn_b_q_io_deq_bits_source),
    .io_deq_bits_address(nodeIn_b_q_io_deq_bits_address)
  );
  Queue_43 nodeOut_c_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_c_q_clock),
    .reset(nodeOut_c_q_reset),
    .io_enq_ready(nodeOut_c_q_io_enq_ready),
    .io_enq_valid(nodeOut_c_q_io_enq_valid),
    .io_enq_bits_opcode(nodeOut_c_q_io_enq_bits_opcode),
    .io_enq_bits_param(nodeOut_c_q_io_enq_bits_param),
    .io_enq_bits_size(nodeOut_c_q_io_enq_bits_size),
    .io_enq_bits_source(nodeOut_c_q_io_enq_bits_source),
    .io_enq_bits_address(nodeOut_c_q_io_enq_bits_address),
    .io_enq_bits_data(nodeOut_c_q_io_enq_bits_data),
    .io_deq_ready(nodeOut_c_q_io_deq_ready),
    .io_deq_valid(nodeOut_c_q_io_deq_valid),
    .io_deq_bits_opcode(nodeOut_c_q_io_deq_bits_opcode),
    .io_deq_bits_param(nodeOut_c_q_io_deq_bits_param),
    .io_deq_bits_size(nodeOut_c_q_io_deq_bits_size),
    .io_deq_bits_source(nodeOut_c_q_io_deq_bits_source),
    .io_deq_bits_address(nodeOut_c_q_io_deq_bits_address),
    .io_deq_bits_data(nodeOut_c_q_io_deq_bits_data)
  );
  Queue_44 nodeOut_e_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_e_q_clock),
    .reset(nodeOut_e_q_reset),
    .io_enq_ready(nodeOut_e_q_io_enq_ready),
    .io_enq_valid(nodeOut_e_q_io_enq_valid),
    .io_enq_bits_sink(nodeOut_e_q_io_enq_bits_sink),
    .io_deq_valid(nodeOut_e_q_io_deq_valid),
    .io_deq_bits_sink(nodeOut_e_q_io_deq_bits_sink)
  );
  assign auto_in_a_ready = nodeOut_a_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_b_valid = nodeIn_b_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 42:15]
  assign auto_in_b_bits_param = nodeIn_b_q_io_deq_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 42:15]
  assign auto_in_b_bits_size = nodeIn_b_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 42:15]
  assign auto_in_b_bits_source = nodeIn_b_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 42:15]
  assign auto_in_b_bits_address = nodeIn_b_q_io_deq_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 42:15]
  assign auto_in_c_ready = nodeOut_c_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_d_valid = nodeIn_d_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_opcode = nodeIn_d_q_io_deq_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_param = nodeIn_d_q_io_deq_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_size = nodeIn_d_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_source = nodeIn_d_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_sink = nodeIn_d_q_io_deq_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_denied = nodeIn_d_q_io_deq_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_data = nodeIn_d_q_io_deq_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_d_bits_corrupt = nodeIn_d_q_io_deq_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/tilelink/Buffer.scala 39:13]
  assign auto_in_e_ready = nodeOut_e_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_out_a_valid = nodeOut_a_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_opcode = nodeOut_a_q_io_deq_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_param = nodeOut_a_q_io_deq_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_size = nodeOut_a_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_source = nodeOut_a_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_address = nodeOut_a_q_io_deq_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_mask = nodeOut_a_q_io_deq_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_a_bits_data = nodeOut_a_q_io_deq_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 38:13]
  assign auto_out_b_ready = nodeIn_b_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_out_c_valid = nodeOut_c_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_opcode = nodeOut_c_q_io_deq_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_param = nodeOut_c_q_io_deq_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_size = nodeOut_c_q_io_deq_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_source = nodeOut_c_q_io_deq_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_address = nodeOut_c_q_io_deq_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_c_bits_data = nodeOut_c_q_io_deq_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 43:15]
  assign auto_out_d_ready = nodeIn_d_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_out_e_valid = nodeOut_e_q_io_deq_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 44:15]
  assign auto_out_e_bits_sink = nodeOut_e_q_io_deq_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/tilelink/Buffer.scala 44:15]
  assign nodeOut_a_q_clock = clock;
  assign nodeOut_a_q_reset = reset;
  assign nodeOut_a_q_io_enq_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_a_q_io_deq_ready = auto_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_clock = clock;
  assign nodeIn_d_q_reset = reset;
  assign nodeIn_d_q_io_enq_valid = auto_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_d_q_io_deq_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeIn_b_q_clock = clock;
  assign nodeIn_b_q_reset = reset;
  assign nodeIn_b_q_io_enq_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_q_io_enq_bits_param = auto_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_q_io_enq_bits_address = auto_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_q_io_deq_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_clock = clock;
  assign nodeOut_c_q_reset = reset;
  assign nodeOut_c_q_io_enq_valid = auto_in_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_opcode = auto_in_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_param = auto_in_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_size = auto_in_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_source = auto_in_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_address = auto_in_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_enq_bits_data = auto_in_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_c_q_io_deq_ready = auto_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeOut_e_q_clock = clock;
  assign nodeOut_e_q_reset = reset;
  assign nodeOut_e_q_io_enq_valid = auto_in_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_e_q_io_enq_bits_sink = auto_in_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module TLBuffer_9(
  input   clock,
  input   reset
);
endmodule
module NonSyncResetSynchronizerPrimitiveShiftReg_d3(
  input   clock,
  input   reset
);
endmodule
module SynchronizerShiftReg_w1_d3(
  input   clock,
  input   reset
);
  wire  output_chain_clock; // @[src/main/scala/util/ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[src/main/scala/util/ShiftReg.scala 45:23]
  NonSyncResetSynchronizerPrimitiveShiftReg_d3 output_chain ( // @[src/main/scala/util/ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset)
  );
  assign output_chain_clock = clock;
  assign output_chain_reset = reset;
endmodule
module IntSyncAsyncCrossingSink(
  input   clock,
  input   reset
);
  wire  chain_clock; // @[src/main/scala/util/ShiftReg.scala 45:23]
  wire  chain_reset; // @[src/main/scala/util/ShiftReg.scala 45:23]
  SynchronizerShiftReg_w1_d3 chain ( // @[src/main/scala/util/ShiftReg.scala 45:23]
    .clock(chain_clock),
    .reset(chain_reset)
  );
  assign chain_clock = clock;
  assign chain_reset = reset;
endmodule
module IntSyncSyncCrossingSink(
  input   clock,
  input   reset
);
endmodule
module IntSyncSyncCrossingSink_1(
  input   clock,
  input   reset
);
endmodule
module IntSyncSyncCrossingSink_2(
  input   clock,
  input   reset
);
endmodule
module AsyncResetRegVec_w1_i0(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module AsyncResetRegVec_w1_i0_1(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_1(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0_1 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module AsyncResetRegVec_w1_i0_2(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_2(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0_2 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module BundleBridgeNexus_13(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_14(
  input   clock,
  input   reset
);
endmodule
module TilePRCIDomain(
  input         auto_tile_reset_domain_tile_hartid_in, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_out_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_a_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_a_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_out_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_master_clock_xing_out_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_tl_master_clock_xing_out_a_bits_mask, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_master_clock_xing_out_a_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_out_b_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_tl_master_clock_xing_out_b_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_c_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_out_c_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_c_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_c_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_tl_master_clock_xing_out_c_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_out_c_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_tl_master_clock_xing_out_c_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_tl_master_clock_xing_out_c_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_out_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_out_d_bits_opcode, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_out_d_bits_param, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_tl_master_clock_xing_out_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_out_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_tl_master_clock_xing_out_d_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_d_bits_denied, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_tl_master_clock_xing_out_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tl_master_clock_xing_out_d_bits_corrupt, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_tl_master_clock_xing_out_e_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_tl_master_clock_xing_out_e_bits_sink, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tap_clock_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_tap_clock_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  tile_reset_domain_auto_tile_buffer_out_a_ready; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_a_valid; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_a_bits_opcode; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_a_bits_param; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_a_bits_size; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_a_bits_source; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [31:0] tile_reset_domain_auto_tile_buffer_out_a_bits_address; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [7:0] tile_reset_domain_auto_tile_buffer_out_a_bits_mask; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [63:0] tile_reset_domain_auto_tile_buffer_out_a_bits_data; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_b_ready; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_b_valid; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_b_bits_param; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_b_bits_size; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_b_bits_source; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [31:0] tile_reset_domain_auto_tile_buffer_out_b_bits_address; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_c_ready; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_c_valid; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_c_bits_opcode; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_c_bits_param; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_c_bits_size; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_c_bits_source; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [31:0] tile_reset_domain_auto_tile_buffer_out_c_bits_address; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [63:0] tile_reset_domain_auto_tile_buffer_out_c_bits_data; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_d_ready; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_d_valid; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_d_bits_opcode; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_d_bits_param; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [2:0] tile_reset_domain_auto_tile_buffer_out_d_bits_size; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_d_bits_source; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_d_bits_sink; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_d_bits_denied; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [63:0] tile_reset_domain_auto_tile_buffer_out_d_bits_data; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_d_bits_corrupt; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_e_ready; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_buffer_out_e_valid; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire [1:0] tile_reset_domain_auto_tile_buffer_out_e_bits_sink; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_tile_hartid_in; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_clock_in_clock; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_auto_clock_in_reset; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_clock; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  tile_reset_domain_reset; // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
  wire  clockNode_auto_in_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  clockNode_auto_in_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  clockNode_auto_out_clock; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  clockNode_auto_out_reset; // @[src/main/scala/prci/ClockGroup.scala 110:107]
  wire  buffer_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_b_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_b_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_b_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_b_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_b_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_c_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_c_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_c_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_c_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_in_c_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_c_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_in_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_in_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_e_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_in_e_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_in_e_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_a_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_a_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_a_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_a_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_a_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_b_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_b_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_b_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_b_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_c_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_c_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_c_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_c_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [31:0] buffer_auto_out_c_bits_address; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_c_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_ready; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_param; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [2:0] buffer_auto_out_d_bits_size; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_source; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_d_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_denied; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [63:0] buffer_auto_out_d_bits_data; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_d_bits_corrupt; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_auto_out_e_valid; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire [1:0] buffer_auto_out_e_bits_sink; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_clock; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  buffer_1_reset; // @[src/main/scala/tilelink/Buffer.scala 69:28]
  wire  intsink_clock; // @[src/main/scala/interrupts/Crossing.scala 78:29]
  wire  intsink_reset; // @[src/main/scala/interrupts/Crossing.scala 78:29]
  wire  intsink_1_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_1_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_2_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_2_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_3_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_3_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsource_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_1_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_1_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_2_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_2_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  trace_clock; // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
  wire  trace_reset; // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
  wire  tracecore_clock; // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
  wire  tracecore_reset; // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
  TileResetDomain tile_reset_domain ( // @[src/main/scala/tile/TilePRCIDomain.scala 45:37]
    .auto_tile_buffer_out_a_ready(tile_reset_domain_auto_tile_buffer_out_a_ready),
    .auto_tile_buffer_out_a_valid(tile_reset_domain_auto_tile_buffer_out_a_valid),
    .auto_tile_buffer_out_a_bits_opcode(tile_reset_domain_auto_tile_buffer_out_a_bits_opcode),
    .auto_tile_buffer_out_a_bits_param(tile_reset_domain_auto_tile_buffer_out_a_bits_param),
    .auto_tile_buffer_out_a_bits_size(tile_reset_domain_auto_tile_buffer_out_a_bits_size),
    .auto_tile_buffer_out_a_bits_source(tile_reset_domain_auto_tile_buffer_out_a_bits_source),
    .auto_tile_buffer_out_a_bits_address(tile_reset_domain_auto_tile_buffer_out_a_bits_address),
    .auto_tile_buffer_out_a_bits_mask(tile_reset_domain_auto_tile_buffer_out_a_bits_mask),
    .auto_tile_buffer_out_a_bits_data(tile_reset_domain_auto_tile_buffer_out_a_bits_data),
    .auto_tile_buffer_out_b_ready(tile_reset_domain_auto_tile_buffer_out_b_ready),
    .auto_tile_buffer_out_b_valid(tile_reset_domain_auto_tile_buffer_out_b_valid),
    .auto_tile_buffer_out_b_bits_param(tile_reset_domain_auto_tile_buffer_out_b_bits_param),
    .auto_tile_buffer_out_b_bits_size(tile_reset_domain_auto_tile_buffer_out_b_bits_size),
    .auto_tile_buffer_out_b_bits_source(tile_reset_domain_auto_tile_buffer_out_b_bits_source),
    .auto_tile_buffer_out_b_bits_address(tile_reset_domain_auto_tile_buffer_out_b_bits_address),
    .auto_tile_buffer_out_c_ready(tile_reset_domain_auto_tile_buffer_out_c_ready),
    .auto_tile_buffer_out_c_valid(tile_reset_domain_auto_tile_buffer_out_c_valid),
    .auto_tile_buffer_out_c_bits_opcode(tile_reset_domain_auto_tile_buffer_out_c_bits_opcode),
    .auto_tile_buffer_out_c_bits_param(tile_reset_domain_auto_tile_buffer_out_c_bits_param),
    .auto_tile_buffer_out_c_bits_size(tile_reset_domain_auto_tile_buffer_out_c_bits_size),
    .auto_tile_buffer_out_c_bits_source(tile_reset_domain_auto_tile_buffer_out_c_bits_source),
    .auto_tile_buffer_out_c_bits_address(tile_reset_domain_auto_tile_buffer_out_c_bits_address),
    .auto_tile_buffer_out_c_bits_data(tile_reset_domain_auto_tile_buffer_out_c_bits_data),
    .auto_tile_buffer_out_d_ready(tile_reset_domain_auto_tile_buffer_out_d_ready),
    .auto_tile_buffer_out_d_valid(tile_reset_domain_auto_tile_buffer_out_d_valid),
    .auto_tile_buffer_out_d_bits_opcode(tile_reset_domain_auto_tile_buffer_out_d_bits_opcode),
    .auto_tile_buffer_out_d_bits_param(tile_reset_domain_auto_tile_buffer_out_d_bits_param),
    .auto_tile_buffer_out_d_bits_size(tile_reset_domain_auto_tile_buffer_out_d_bits_size),
    .auto_tile_buffer_out_d_bits_source(tile_reset_domain_auto_tile_buffer_out_d_bits_source),
    .auto_tile_buffer_out_d_bits_sink(tile_reset_domain_auto_tile_buffer_out_d_bits_sink),
    .auto_tile_buffer_out_d_bits_denied(tile_reset_domain_auto_tile_buffer_out_d_bits_denied),
    .auto_tile_buffer_out_d_bits_data(tile_reset_domain_auto_tile_buffer_out_d_bits_data),
    .auto_tile_buffer_out_d_bits_corrupt(tile_reset_domain_auto_tile_buffer_out_d_bits_corrupt),
    .auto_tile_buffer_out_e_ready(tile_reset_domain_auto_tile_buffer_out_e_ready),
    .auto_tile_buffer_out_e_valid(tile_reset_domain_auto_tile_buffer_out_e_valid),
    .auto_tile_buffer_out_e_bits_sink(tile_reset_domain_auto_tile_buffer_out_e_bits_sink),
    .auto_tile_hartid_in(tile_reset_domain_auto_tile_hartid_in),
    .auto_clock_in_clock(tile_reset_domain_auto_clock_in_clock),
    .auto_clock_in_reset(tile_reset_domain_auto_clock_in_reset),
    .clock(tile_reset_domain_clock),
    .reset(tile_reset_domain_reset)
  );
  FixedClockBroadcast_6 clockNode ( // @[src/main/scala/prci/ClockGroup.scala 110:107]
    .auto_in_clock(clockNode_auto_in_clock),
    .auto_in_reset(clockNode_auto_in_reset),
    .auto_out_clock(clockNode_auto_out_clock),
    .auto_out_reset(clockNode_auto_out_reset)
  );
  TLBuffer_8 buffer ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_b_ready(buffer_auto_in_b_ready),
    .auto_in_b_valid(buffer_auto_in_b_valid),
    .auto_in_b_bits_param(buffer_auto_in_b_bits_param),
    .auto_in_b_bits_size(buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(buffer_auto_in_b_bits_address),
    .auto_in_c_ready(buffer_auto_in_c_ready),
    .auto_in_c_valid(buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(buffer_auto_in_c_bits_data),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_in_e_ready(buffer_auto_in_e_ready),
    .auto_in_e_valid(buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_b_ready(buffer_auto_out_b_ready),
    .auto_out_b_valid(buffer_auto_out_b_valid),
    .auto_out_b_bits_param(buffer_auto_out_b_bits_param),
    .auto_out_b_bits_address(buffer_auto_out_b_bits_address),
    .auto_out_c_ready(buffer_auto_out_c_ready),
    .auto_out_c_valid(buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(buffer_auto_out_c_bits_data),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_auto_out_d_bits_corrupt),
    .auto_out_e_valid(buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(buffer_auto_out_e_bits_sink)
  );
  TLBuffer_9 buffer_1 ( // @[src/main/scala/tilelink/Buffer.scala 69:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset)
  );
  IntSyncAsyncCrossingSink intsink ( // @[src/main/scala/interrupts/Crossing.scala 78:29]
    .clock(intsink_clock),
    .reset(intsink_reset)
  );
  IntSyncSyncCrossingSink intsink_1 ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_1_clock),
    .reset(intsink_1_reset)
  );
  IntSyncSyncCrossingSink_1 intsink_2 ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_2_clock),
    .reset(intsink_2_reset)
  );
  IntSyncSyncCrossingSink_2 intsink_3 ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_3_clock),
    .reset(intsink_3_reset)
  );
  IntSyncCrossingSource intsource ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_clock),
    .reset(intsource_reset)
  );
  IntSyncCrossingSource_1 intsource_1 ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_1_clock),
    .reset(intsource_1_reset)
  );
  IntSyncCrossingSource_2 intsource_2 ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_2_clock),
    .reset(intsource_2_reset)
  );
  BundleBridgeNexus_13 trace ( // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
    .clock(trace_clock),
    .reset(trace_reset)
  );
  BundleBridgeNexus_14 tracecore ( // @[src/main/scala/prci/BundleBridgeBlockDuringReset.scala 20:27]
    .clock(tracecore_clock),
    .reset(tracecore_reset)
  );
  assign auto_tl_master_clock_xing_out_a_valid = buffer_auto_out_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_param = buffer_auto_out_a_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_size = buffer_auto_out_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_source = buffer_auto_out_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_address = buffer_auto_out_a_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_mask = buffer_auto_out_a_bits_mask; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_a_bits_data = buffer_auto_out_a_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_b_ready = buffer_auto_out_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_valid = buffer_auto_out_c_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_opcode = buffer_auto_out_c_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_param = buffer_auto_out_c_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_size = buffer_auto_out_c_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_source = buffer_auto_out_c_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_address = buffer_auto_out_c_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_c_bits_data = buffer_auto_out_c_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_d_ready = buffer_auto_out_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_e_valid = buffer_auto_out_e_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign auto_tl_master_clock_xing_out_e_bits_sink = buffer_auto_out_e_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tile_reset_domain_auto_tile_buffer_out_a_ready = buffer_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_b_valid = buffer_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_b_bits_param = buffer_auto_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_b_bits_size = buffer_auto_in_b_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_b_bits_source = buffer_auto_in_b_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_b_bits_address = buffer_auto_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_c_ready = buffer_auto_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_valid = buffer_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_param = buffer_auto_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_size = buffer_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_source = buffer_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_data = buffer_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_buffer_out_e_ready = buffer_auto_in_e_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_reset_domain_auto_tile_hartid_in = auto_tile_reset_domain_tile_hartid_in; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tile_reset_domain_auto_clock_in_clock = clockNode_auto_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_reset_domain_auto_clock_in_reset = clockNode_auto_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign clockNode_auto_in_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clockNode_auto_in_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_auto_in_a_valid = tile_reset_domain_auto_tile_buffer_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_opcode = tile_reset_domain_auto_tile_buffer_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_param = tile_reset_domain_auto_tile_buffer_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_size = tile_reset_domain_auto_tile_buffer_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_source = tile_reset_domain_auto_tile_buffer_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_address = tile_reset_domain_auto_tile_buffer_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_mask = tile_reset_domain_auto_tile_buffer_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_a_bits_data = tile_reset_domain_auto_tile_buffer_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_b_ready = tile_reset_domain_auto_tile_buffer_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_valid = tile_reset_domain_auto_tile_buffer_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_opcode = tile_reset_domain_auto_tile_buffer_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_param = tile_reset_domain_auto_tile_buffer_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_size = tile_reset_domain_auto_tile_buffer_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_source = tile_reset_domain_auto_tile_buffer_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_address = tile_reset_domain_auto_tile_buffer_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_c_bits_data = tile_reset_domain_auto_tile_buffer_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_d_ready = tile_reset_domain_auto_tile_buffer_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_e_valid = tile_reset_domain_auto_tile_buffer_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_in_e_bits_sink = tile_reset_domain_auto_tile_buffer_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign buffer_auto_out_a_ready = auto_tl_master_clock_xing_out_a_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_valid = auto_tl_master_clock_xing_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_param = auto_tl_master_clock_xing_out_b_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_b_bits_address = auto_tl_master_clock_xing_out_b_bits_address; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_c_ready = auto_tl_master_clock_xing_out_c_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_valid = auto_tl_master_clock_xing_out_d_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_opcode = auto_tl_master_clock_xing_out_d_bits_opcode; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_param = auto_tl_master_clock_xing_out_d_bits_param; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_size = auto_tl_master_clock_xing_out_d_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_source = auto_tl_master_clock_xing_out_d_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_sink = auto_tl_master_clock_xing_out_d_bits_sink; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_denied = auto_tl_master_clock_xing_out_d_bits_denied; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_data = auto_tl_master_clock_xing_out_d_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_auto_out_d_bits_corrupt = auto_tl_master_clock_xing_out_d_bits_corrupt; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign buffer_1_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign buffer_1_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_1_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_1_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_2_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_2_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_3_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsink_3_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_1_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_1_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_2_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign intsource_2_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign trace_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign trace_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tracecore_clock = auto_tap_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign tracecore_reset = auto_tap_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module IntXbar_2(
  input   clock,
  input   reset
);
endmodule
module IntXbar_3(
  input   clock,
  input   reset
);
endmodule
module IntXbar_4(
  input   clock,
  input   reset
);
endmodule
module BundleBridgeNexus_15(
  input   clock,
  input   reset,
  output  auto_out // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  outputs_0 = 1'h0; // @[src/main/scala/subsystem/HasTiles.scala 159:32]
  assign auto_out = outputs_0; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/BundleBridge.scala 152:67]
endmodule
module BundleBridgeNexus_16(
  input   clock,
  input   reset
);
endmodule
module IntSyncXbar(
  input   clock,
  input   reset
);
endmodule
module AsyncResetRegVec_w1_i0_3(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_3(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0_3 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module NullIntSource(
  input   clock,
  input   reset
);
endmodule
module AsyncResetRegVec_w2_i0(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_4(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w2_i0 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module NullIntSource_1(
  input   clock,
  input   reset
);
endmodule
module AsyncResetRegVec_w1_i0_4(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_5(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0_4 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module AsyncResetRegVec_w1_i0_5(
  input   clock,
  input   reset
);
endmodule
module IntSyncCrossingSource_6(
  input   clock,
  input   reset
);
  wire  reg__clock; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  wire  reg__reset; // @[src/main/scala/util/AsyncResetReg.scala 86:21]
  AsyncResetRegVec_w1_i0_5 reg_ ( // @[src/main/scala/util/AsyncResetReg.scala 86:21]
    .clock(reg__clock),
    .reset(reg__reset)
  );
  assign reg__clock = clock;
  assign reg__reset = reset;
endmodule
module IntSyncSyncCrossingSink_3(
  input   clock,
  input   reset
);
endmodule
module IntSyncSyncCrossingSink_4(
  input   clock,
  input   reset
);
endmodule
module IntSyncSyncCrossingSink_5(
  input   clock,
  input   reset
);
endmodule
module TLROM(
  input         clock,
  input         reset,
  output        auto_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [4:0]  auto_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [4:0]  auto_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_d_bits_data // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  index = auto_in_a_bits_address[3]; // @[src/main/scala/devices/tilelink/BootROM.scala 53:34]
  wire [11:0] high = auto_in_a_bits_address[15:4]; // @[src/main/scala/devices/tilelink/BootROM.scala 54:64]
  wire  line_1254_clock;
  wire  line_1254_reset;
  wire  line_1254_valid;
  reg  line_1254_valid_reg;
  wire  line_1255_clock;
  wire  line_1255_reset;
  wire  line_1255_valid;
  reg  line_1255_valid_reg;
  wire [63:0] _GEN_3 = index ? 64'h28067 : 64'h1f292930010029b; // @[src/main/scala/devices/tilelink/BootROM.scala 55:{47,47}]
  GEN_w1_line #(.COVER_INDEX(1254)) line_1254 (
    .clock(line_1254_clock),
    .reset(line_1254_reset),
    .valid(line_1254_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1255)) line_1255 (
    .clock(line_1255_clock),
    .reset(line_1255_reset),
    .valid(line_1255_valid)
  );
  assign line_1254_clock = clock;
  assign line_1254_reset = reset;
  assign line_1254_valid = ~index ^ line_1254_valid_reg;
  assign line_1255_clock = clock;
  assign line_1255_reset = reset;
  assign line_1255_valid = index ^ line_1255_valid_reg;
  assign auto_in_a_ready = auto_in_d_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_in_d_valid = auto_in_a_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_in_d_bits_data = |high ? 64'h0 : _GEN_3; // @[src/main/scala/devices/tilelink/BootROM.scala 55:47]
  always @(posedge clock) begin
    line_1254_valid_reg <= ~index;
    line_1255_valid_reg <= index;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1254_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1255_valid_reg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockSinkDomain(
  output        auto_bootrom_in_a_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bootrom_in_a_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_bootrom_in_a_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [4:0]  auto_bootrom_in_a_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [28:0] auto_bootrom_in_a_bits_address, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_bootrom_in_d_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_bootrom_in_d_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_bootrom_in_d_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [4:0]  auto_bootrom_in_d_bits_source, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_bootrom_in_d_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_clock_in_clock, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_clock_in_reset, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        clock, // @[src/main/scala/prci/ClockDomain.scala 17:19]
  output        reset // @[src/main/scala/prci/ClockDomain.scala 18:19]
);
  wire  bootrom_clock; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire  bootrom_reset; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire  bootrom_auto_in_a_ready; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire  bootrom_auto_in_a_valid; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [1:0] bootrom_auto_in_a_bits_size; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [4:0] bootrom_auto_in_a_bits_source; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [28:0] bootrom_auto_in_a_bits_address; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire  bootrom_auto_in_d_ready; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire  bootrom_auto_in_d_valid; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [1:0] bootrom_auto_in_d_bits_size; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [4:0] bootrom_auto_in_d_bits_source; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  wire [63:0] bootrom_auto_in_d_bits_data; // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
  TLROM bootrom ( // @[src/main/scala/devices/tilelink/BootROM.scala 86:17]
    .clock(bootrom_clock),
    .reset(bootrom_reset),
    .auto_in_a_ready(bootrom_auto_in_a_ready),
    .auto_in_a_valid(bootrom_auto_in_a_valid),
    .auto_in_a_bits_size(bootrom_auto_in_a_bits_size),
    .auto_in_a_bits_source(bootrom_auto_in_a_bits_source),
    .auto_in_a_bits_address(bootrom_auto_in_a_bits_address),
    .auto_in_d_ready(bootrom_auto_in_d_ready),
    .auto_in_d_valid(bootrom_auto_in_d_valid),
    .auto_in_d_bits_size(bootrom_auto_in_d_bits_size),
    .auto_in_d_bits_source(bootrom_auto_in_d_bits_source),
    .auto_in_d_bits_data(bootrom_auto_in_d_bits_data)
  );
  assign auto_bootrom_in_a_ready = bootrom_auto_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bootrom_in_d_valid = bootrom_auto_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bootrom_in_d_bits_size = bootrom_auto_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bootrom_in_d_bits_source = bootrom_auto_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_bootrom_in_d_bits_data = bootrom_auto_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_clock = auto_clock_in_clock; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_reset = auto_clock_in_reset; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_auto_in_a_valid = auto_bootrom_in_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_auto_in_a_bits_size = auto_bootrom_in_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_auto_in_a_bits_source = auto_bootrom_in_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_auto_in_a_bits_address = auto_bootrom_in_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign bootrom_auto_in_d_ready = auto_bootrom_in_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module ExampleFuzzSystem(
  input         clock,
  input         reset,
  input         mem_axi4_0_aw_ready, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_aw_valid, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [3:0]  mem_axi4_0_aw_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [31:0] mem_axi4_0_aw_bits_addr, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [7:0]  mem_axi4_0_aw_bits_len, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [2:0]  mem_axi4_0_aw_bits_size, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [1:0]  mem_axi4_0_aw_bits_burst, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input         mem_axi4_0_w_ready, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_w_valid, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [63:0] mem_axi4_0_w_bits_data, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [7:0]  mem_axi4_0_w_bits_strb, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_w_bits_last, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_b_ready, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input         mem_axi4_0_b_valid, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input  [3:0]  mem_axi4_0_b_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input  [1:0]  mem_axi4_0_b_bits_resp, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input         mem_axi4_0_ar_ready, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_ar_valid, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [3:0]  mem_axi4_0_ar_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [31:0] mem_axi4_0_ar_bits_addr, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [7:0]  mem_axi4_0_ar_bits_len, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [2:0]  mem_axi4_0_ar_bits_size, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output [1:0]  mem_axi4_0_ar_bits_burst, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  output        mem_axi4_0_r_ready, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input         mem_axi4_0_r_valid, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input  [3:0]  mem_axi4_0_r_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input  [63:0] mem_axi4_0_r_bits_data, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input  [1:0]  mem_axi4_0_r_bits_resp, // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
  input         mem_axi4_0_r_bits_last // @[src/main/scala/diplomacy/Nodes.scala 1713:17]
);
  wire  ibus_auto_clock_in_clock; // @[src/main/scala/subsystem/BaseSubsystem.scala 49:24]
  wire  ibus_auto_clock_in_reset; // @[src/main/scala/subsystem/BaseSubsystem.scala 49:24]
  wire  ibus_clock; // @[src/main/scala/subsystem/BaseSubsystem.scala 49:24]
  wire  ibus_reset; // @[src/main/scala/subsystem/BaseSubsystem.scala 49:24]
  wire  dummyClockGroupSourceNode_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset; // @[src/main/scala/prci/ClockGroup.scala 82:81]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [31:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [28:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [7:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [2:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [1:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire [63:0] subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_1_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_1_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_0_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_fixedClockNode_out_0_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_clock; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_sbus_reset; // @[src/main/scala/subsystem/SystemBus.scala 24:26]
  wire  subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_pbus_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_pbus_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock; // @[src/main/scala/subsystem/FrontBus.scala 22:26]
  wire  subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset; // @[src/main/scala/subsystem/FrontBus.scala 22:26]
  wire  subsystem_fbus_clock; // @[src/main/scala/subsystem/FrontBus.scala 22:26]
  wire  subsystem_fbus_reset; // @[src/main/scala/subsystem/FrontBus.scala 22:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [4:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [28:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [4:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_fixedClockNode_out_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_fixedClockNode_out_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_a_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_a_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_a_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_bus_xing_in_a_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [28:0] subsystem_cbus_auto_bus_xing_in_a_bits_address; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [7:0] subsystem_cbus_auto_bus_xing_in_a_bits_mask; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_ready; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_valid; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_d_bits_opcode; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_bus_xing_in_d_bits_param; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [2:0] subsystem_cbus_auto_bus_xing_in_d_bits_size; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [1:0] subsystem_cbus_auto_bus_xing_in_d_bits_source; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_bits_sink; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_bits_denied; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire [63:0] subsystem_cbus_auto_bus_xing_in_d_bits_data; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_auto_bus_xing_in_d_bits_corrupt; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_clock; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_cbus_reset; // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [1:0] subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_a_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_a_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_a_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_bus_xing_in_a_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [31:0] subsystem_mbus_auto_bus_xing_in_a_bits_address; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [7:0] subsystem_mbus_auto_bus_xing_in_a_bits_mask; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_bus_xing_in_a_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_ready; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_valid; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_d_bits_opcode; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [2:0] subsystem_mbus_auto_bus_xing_in_d_bits_size; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [3:0] subsystem_mbus_auto_bus_xing_in_d_bits_source; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_bits_denied; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire [63:0] subsystem_mbus_auto_bus_xing_in_d_bits_data; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_auto_bus_xing_in_d_bits_corrupt; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_clock; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_mbus_reset; // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [3:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [31:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [7:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [63:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [3:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [63:0] subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [31:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [7:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [63:0] subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_b_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [31:0] subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_c_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [31:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_address; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [63:0] subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [2:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [63:0] subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_coherent_jbar_in_e_valid; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire [1:0] subsystem_l2_wrapper_auto_coherent_jbar_in_e_bits_sink; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_clock; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  subsystem_l2_wrapper_reset; // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
  wire  tile_prci_domain_auto_tile_reset_domain_tile_hartid_in; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_ready; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_a_valid; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [7:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [63:0] tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_b_ready; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_b_valid; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_c_ready; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_c_valid; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [31:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [63:0] tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_ready; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_valid; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [2:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [63:0] tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tl_master_clock_xing_out_e_valid; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire [1:0] tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tap_clock_in_clock; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_auto_tap_clock_in_reset; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_clock; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  tile_prci_domain_reset; // @[src/main/scala/subsystem/HasTiles.scala 250:38]
  wire  xbar_clock; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  xbar_reset; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  xbar_1_clock; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  xbar_1_reset; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  xbar_2_clock; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  xbar_2_reset; // @[src/main/scala/interrupts/Xbar.scala 50:26]
  wire  tileHartIdNexusNode_clock; // @[src/main/scala/subsystem/HasTiles.scala 156:39]
  wire  tileHartIdNexusNode_reset; // @[src/main/scala/subsystem/HasTiles.scala 156:39]
  wire  tileHartIdNexusNode_auto_out; // @[src/main/scala/subsystem/HasTiles.scala 156:39]
  wire  broadcast_clock; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  broadcast_reset; // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
  wire  xbar_3_clock; // @[src/main/scala/interrupts/Xbar.scala 57:26]
  wire  xbar_3_reset; // @[src/main/scala/interrupts/Xbar.scala 57:26]
  wire  intsource_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  null_int_source_clock; // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
  wire  null_int_source_reset; // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
  wire  intsource_1_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_1_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  null_int_source_1_clock; // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
  wire  null_int_source_1_reset; // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
  wire  intsource_2_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_2_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_3_clock; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsource_3_reset; // @[src/main/scala/interrupts/Crossing.scala 28:31]
  wire  intsink_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_1_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_1_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_2_clock; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  intsink_2_reset; // @[src/main/scala/interrupts/Crossing.scala 99:29]
  wire  bootROMDomainWrapper_auto_bootrom_in_a_ready; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_a_valid; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [1:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_size; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [4:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_source; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [28:0] bootROMDomainWrapper_auto_bootrom_in_a_bits_address; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_d_ready; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_auto_bootrom_in_d_valid; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [1:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_size; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [4:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_source; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire [63:0] bootROMDomainWrapper_auto_bootrom_in_d_bits_data; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_auto_clock_in_clock; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_auto_clock_in_reset; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_clock; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  wire  bootROMDomainWrapper_reset; // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
  InterruptBusWrapper ibus ( // @[src/main/scala/subsystem/BaseSubsystem.scala 49:24]
    .auto_clock_in_clock(ibus_auto_clock_in_clock),
    .auto_clock_in_reset(ibus_auto_clock_in_reset),
    .clock(ibus_clock),
    .reset(ibus_reset)
  );
  SimpleClockGroupSource dummyClockGroupSourceNode ( // @[src/main/scala/prci/ClockGroup.scala 82:81]
    .clock(dummyClockGroupSourceNode_clock),
    .reset(dummyClockGroupSourceNode_reset),
    .auto_out_member_subsystem_sbus_5_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock),
    .auto_out_member_subsystem_sbus_5_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset),
    .auto_out_member_subsystem_sbus_4_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock),
    .auto_out_member_subsystem_sbus_4_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset),
    .auto_out_member_subsystem_sbus_3_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock),
    .auto_out_member_subsystem_sbus_3_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset),
    .auto_out_member_subsystem_sbus_2_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock),
    .auto_out_member_subsystem_sbus_2_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset),
    .auto_out_member_subsystem_sbus_1_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock),
    .auto_out_member_subsystem_sbus_1_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset),
    .auto_out_member_subsystem_sbus_0_clock(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock),
    .auto_out_member_subsystem_sbus_0_reset(dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset)
  );
  SystemBus subsystem_sbus ( // @[src/main/scala/subsystem/SystemBus.scala 24:26]
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_ready(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_valid(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask),
    .auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data),
    .auto_coupler_from_tile_tl_master_clock_xing_in_b_ready(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_ready),
    .auto_coupler_from_tile_tl_master_clock_xing_in_b_valid(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid),
    .auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param),
    .auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_ready(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_valid(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_valid),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address),
    .auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_ready(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_valid(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data),
    .auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt),
    .auto_coupler_from_tile_tl_master_clock_xing_in_e_valid(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_valid),
    .auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink(
      subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid),
    .auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt(
      subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt),
    .auto_fixedClockNode_out_1_clock(subsystem_sbus_auto_fixedClockNode_out_1_clock),
    .auto_fixedClockNode_out_1_reset(subsystem_sbus_auto_fixedClockNode_out_1_reset),
    .auto_fixedClockNode_out_0_clock(subsystem_sbus_auto_fixedClockNode_out_0_clock),
    .auto_fixedClockNode_out_0_reset(subsystem_sbus_auto_fixedClockNode_out_0_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock),
    .auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock),
    .auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset),
    .auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock),
    .auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock),
    .auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset(
      subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset),
    .clock(subsystem_sbus_clock),
    .reset(subsystem_sbus_reset)
  );
  PeripheryBus subsystem_pbus ( // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
    .auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock(
      subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock),
    .auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset(
      subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset),
    .clock(subsystem_pbus_clock),
    .reset(subsystem_pbus_reset)
  );
  FrontBus subsystem_fbus ( // @[src/main/scala/subsystem/FrontBus.scala 22:26]
    .auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock(
      subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock),
    .auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset(
      subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset),
    .clock(subsystem_fbus_clock),
    .reset(subsystem_fbus_reset)
  );
  PeripheryBus_1 subsystem_cbus ( // @[src/main/scala/subsystem/PeripheryBus.scala 31:26]
    .auto_coupler_to_bootrom_fragmenter_out_a_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready),
    .auto_coupler_to_bootrom_fragmenter_out_a_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_size(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_source(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source),
    .auto_coupler_to_bootrom_fragmenter_out_a_bits_address(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address),
    .auto_coupler_to_bootrom_fragmenter_out_d_ready(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready),
    .auto_coupler_to_bootrom_fragmenter_out_d_valid(subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_size(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_source(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source),
    .auto_coupler_to_bootrom_fragmenter_out_d_bits_data(
      subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data),
    .auto_fixedClockNode_out_clock(subsystem_cbus_auto_fixedClockNode_out_clock),
    .auto_fixedClockNode_out_reset(subsystem_cbus_auto_fixedClockNode_out_reset),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock),
    .auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset),
    .auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock),
    .auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset(
      subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset),
    .auto_bus_xing_in_a_ready(subsystem_cbus_auto_bus_xing_in_a_ready),
    .auto_bus_xing_in_a_valid(subsystem_cbus_auto_bus_xing_in_a_valid),
    .auto_bus_xing_in_a_bits_size(subsystem_cbus_auto_bus_xing_in_a_bits_size),
    .auto_bus_xing_in_a_bits_source(subsystem_cbus_auto_bus_xing_in_a_bits_source),
    .auto_bus_xing_in_a_bits_address(subsystem_cbus_auto_bus_xing_in_a_bits_address),
    .auto_bus_xing_in_a_bits_mask(subsystem_cbus_auto_bus_xing_in_a_bits_mask),
    .auto_bus_xing_in_d_ready(subsystem_cbus_auto_bus_xing_in_d_ready),
    .auto_bus_xing_in_d_valid(subsystem_cbus_auto_bus_xing_in_d_valid),
    .auto_bus_xing_in_d_bits_opcode(subsystem_cbus_auto_bus_xing_in_d_bits_opcode),
    .auto_bus_xing_in_d_bits_param(subsystem_cbus_auto_bus_xing_in_d_bits_param),
    .auto_bus_xing_in_d_bits_size(subsystem_cbus_auto_bus_xing_in_d_bits_size),
    .auto_bus_xing_in_d_bits_source(subsystem_cbus_auto_bus_xing_in_d_bits_source),
    .auto_bus_xing_in_d_bits_sink(subsystem_cbus_auto_bus_xing_in_d_bits_sink),
    .auto_bus_xing_in_d_bits_denied(subsystem_cbus_auto_bus_xing_in_d_bits_denied),
    .auto_bus_xing_in_d_bits_data(subsystem_cbus_auto_bus_xing_in_d_bits_data),
    .auto_bus_xing_in_d_bits_corrupt(subsystem_cbus_auto_bus_xing_in_d_bits_corrupt),
    .clock(subsystem_cbus_clock),
    .reset(subsystem_cbus_reset)
  );
  MemoryBus subsystem_mbus ( // @[src/main/scala/subsystem/MemoryBus.scala 25:26]
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp),
    .auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last(
      subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last),
    .auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock(
      subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),
    .auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset(
      subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),
    .auto_bus_xing_in_a_ready(subsystem_mbus_auto_bus_xing_in_a_ready),
    .auto_bus_xing_in_a_valid(subsystem_mbus_auto_bus_xing_in_a_valid),
    .auto_bus_xing_in_a_bits_opcode(subsystem_mbus_auto_bus_xing_in_a_bits_opcode),
    .auto_bus_xing_in_a_bits_size(subsystem_mbus_auto_bus_xing_in_a_bits_size),
    .auto_bus_xing_in_a_bits_source(subsystem_mbus_auto_bus_xing_in_a_bits_source),
    .auto_bus_xing_in_a_bits_address(subsystem_mbus_auto_bus_xing_in_a_bits_address),
    .auto_bus_xing_in_a_bits_mask(subsystem_mbus_auto_bus_xing_in_a_bits_mask),
    .auto_bus_xing_in_a_bits_data(subsystem_mbus_auto_bus_xing_in_a_bits_data),
    .auto_bus_xing_in_d_ready(subsystem_mbus_auto_bus_xing_in_d_ready),
    .auto_bus_xing_in_d_valid(subsystem_mbus_auto_bus_xing_in_d_valid),
    .auto_bus_xing_in_d_bits_opcode(subsystem_mbus_auto_bus_xing_in_d_bits_opcode),
    .auto_bus_xing_in_d_bits_size(subsystem_mbus_auto_bus_xing_in_d_bits_size),
    .auto_bus_xing_in_d_bits_source(subsystem_mbus_auto_bus_xing_in_d_bits_source),
    .auto_bus_xing_in_d_bits_denied(subsystem_mbus_auto_bus_xing_in_d_bits_denied),
    .auto_bus_xing_in_d_bits_data(subsystem_mbus_auto_bus_xing_in_d_bits_data),
    .auto_bus_xing_in_d_bits_corrupt(subsystem_mbus_auto_bus_xing_in_d_bits_corrupt),
    .clock(subsystem_mbus_clock),
    .reset(subsystem_mbus_reset)
  );
  CoherenceManagerWrapper subsystem_l2_wrapper ( // @[src/main/scala/subsystem/BankedL2Params.scala 48:31]
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data),
    .auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt(
      subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt),
    .auto_coherent_jbar_in_a_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready),
    .auto_coherent_jbar_in_a_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid),
    .auto_coherent_jbar_in_a_bits_opcode(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode),
    .auto_coherent_jbar_in_a_bits_param(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_param),
    .auto_coherent_jbar_in_a_bits_size(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size),
    .auto_coherent_jbar_in_a_bits_source(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source),
    .auto_coherent_jbar_in_a_bits_address(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address),
    .auto_coherent_jbar_in_a_bits_mask(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask),
    .auto_coherent_jbar_in_a_bits_data(subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data),
    .auto_coherent_jbar_in_b_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_b_ready),
    .auto_coherent_jbar_in_b_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid),
    .auto_coherent_jbar_in_b_bits_param(subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param),
    .auto_coherent_jbar_in_b_bits_address(subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address),
    .auto_coherent_jbar_in_c_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready),
    .auto_coherent_jbar_in_c_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_c_valid),
    .auto_coherent_jbar_in_c_bits_opcode(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_opcode),
    .auto_coherent_jbar_in_c_bits_param(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_param),
    .auto_coherent_jbar_in_c_bits_size(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_size),
    .auto_coherent_jbar_in_c_bits_source(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_source),
    .auto_coherent_jbar_in_c_bits_address(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_address),
    .auto_coherent_jbar_in_c_bits_data(subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_data),
    .auto_coherent_jbar_in_d_ready(subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready),
    .auto_coherent_jbar_in_d_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid),
    .auto_coherent_jbar_in_d_bits_opcode(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode),
    .auto_coherent_jbar_in_d_bits_param(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param),
    .auto_coherent_jbar_in_d_bits_size(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size),
    .auto_coherent_jbar_in_d_bits_source(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source),
    .auto_coherent_jbar_in_d_bits_sink(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink),
    .auto_coherent_jbar_in_d_bits_denied(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied),
    .auto_coherent_jbar_in_d_bits_data(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data),
    .auto_coherent_jbar_in_d_bits_corrupt(subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt),
    .auto_coherent_jbar_in_e_valid(subsystem_l2_wrapper_auto_coherent_jbar_in_e_valid),
    .auto_coherent_jbar_in_e_bits_sink(subsystem_l2_wrapper_auto_coherent_jbar_in_e_bits_sink),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock),
    .auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset),
    .auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock),
    .auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset(
      subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset),
    .clock(subsystem_l2_wrapper_clock),
    .reset(subsystem_l2_wrapper_reset)
  );
  TilePRCIDomain tile_prci_domain ( // @[src/main/scala/subsystem/HasTiles.scala 250:38]
    .auto_tile_reset_domain_tile_hartid_in(tile_prci_domain_auto_tile_reset_domain_tile_hartid_in),
    .auto_tl_master_clock_xing_out_a_ready(tile_prci_domain_auto_tl_master_clock_xing_out_a_ready),
    .auto_tl_master_clock_xing_out_a_valid(tile_prci_domain_auto_tl_master_clock_xing_out_a_valid),
    .auto_tl_master_clock_xing_out_a_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode),
    .auto_tl_master_clock_xing_out_a_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param),
    .auto_tl_master_clock_xing_out_a_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size),
    .auto_tl_master_clock_xing_out_a_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source),
    .auto_tl_master_clock_xing_out_a_bits_address(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address),
    .auto_tl_master_clock_xing_out_a_bits_mask(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask),
    .auto_tl_master_clock_xing_out_a_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data),
    .auto_tl_master_clock_xing_out_b_ready(tile_prci_domain_auto_tl_master_clock_xing_out_b_ready),
    .auto_tl_master_clock_xing_out_b_valid(tile_prci_domain_auto_tl_master_clock_xing_out_b_valid),
    .auto_tl_master_clock_xing_out_b_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_param),
    .auto_tl_master_clock_xing_out_b_bits_address(tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_address),
    .auto_tl_master_clock_xing_out_c_ready(tile_prci_domain_auto_tl_master_clock_xing_out_c_ready),
    .auto_tl_master_clock_xing_out_c_valid(tile_prci_domain_auto_tl_master_clock_xing_out_c_valid),
    .auto_tl_master_clock_xing_out_c_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode),
    .auto_tl_master_clock_xing_out_c_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param),
    .auto_tl_master_clock_xing_out_c_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size),
    .auto_tl_master_clock_xing_out_c_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source),
    .auto_tl_master_clock_xing_out_c_bits_address(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address),
    .auto_tl_master_clock_xing_out_c_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data),
    .auto_tl_master_clock_xing_out_d_ready(tile_prci_domain_auto_tl_master_clock_xing_out_d_ready),
    .auto_tl_master_clock_xing_out_d_valid(tile_prci_domain_auto_tl_master_clock_xing_out_d_valid),
    .auto_tl_master_clock_xing_out_d_bits_opcode(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode),
    .auto_tl_master_clock_xing_out_d_bits_param(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param),
    .auto_tl_master_clock_xing_out_d_bits_size(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size),
    .auto_tl_master_clock_xing_out_d_bits_source(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source),
    .auto_tl_master_clock_xing_out_d_bits_sink(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink),
    .auto_tl_master_clock_xing_out_d_bits_denied(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied),
    .auto_tl_master_clock_xing_out_d_bits_data(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data),
    .auto_tl_master_clock_xing_out_d_bits_corrupt(tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt),
    .auto_tl_master_clock_xing_out_e_valid(tile_prci_domain_auto_tl_master_clock_xing_out_e_valid),
    .auto_tl_master_clock_xing_out_e_bits_sink(tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink),
    .auto_tap_clock_in_clock(tile_prci_domain_auto_tap_clock_in_clock),
    .auto_tap_clock_in_reset(tile_prci_domain_auto_tap_clock_in_reset),
    .clock(tile_prci_domain_clock),
    .reset(tile_prci_domain_reset)
  );
  IntXbar_2 xbar ( // @[src/main/scala/interrupts/Xbar.scala 50:26]
    .clock(xbar_clock),
    .reset(xbar_reset)
  );
  IntXbar_3 xbar_1 ( // @[src/main/scala/interrupts/Xbar.scala 50:26]
    .clock(xbar_1_clock),
    .reset(xbar_1_reset)
  );
  IntXbar_4 xbar_2 ( // @[src/main/scala/interrupts/Xbar.scala 50:26]
    .clock(xbar_2_clock),
    .reset(xbar_2_reset)
  );
  BundleBridgeNexus_15 tileHartIdNexusNode ( // @[src/main/scala/subsystem/HasTiles.scala 156:39]
    .clock(tileHartIdNexusNode_clock),
    .reset(tileHartIdNexusNode_reset),
    .auto_out(tileHartIdNexusNode_auto_out)
  );
  BundleBridgeNexus_16 broadcast ( // @[src/main/scala/diplomacy/BundleBridge.scala 197:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset)
  );
  IntSyncXbar xbar_3 ( // @[src/main/scala/interrupts/Xbar.scala 57:26]
    .clock(xbar_3_clock),
    .reset(xbar_3_reset)
  );
  IntSyncCrossingSource_3 intsource ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_clock),
    .reset(intsource_reset)
  );
  NullIntSource null_int_source ( // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
    .clock(null_int_source_clock),
    .reset(null_int_source_reset)
  );
  IntSyncCrossingSource_4 intsource_1 ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_1_clock),
    .reset(intsource_1_reset)
  );
  NullIntSource_1 null_int_source_1 ( // @[src/main/scala/interrupts/NullIntSource.scala 22:37]
    .clock(null_int_source_1_clock),
    .reset(null_int_source_1_reset)
  );
  IntSyncCrossingSource_5 intsource_2 ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_2_clock),
    .reset(intsource_2_reset)
  );
  IntSyncCrossingSource_6 intsource_3 ( // @[src/main/scala/interrupts/Crossing.scala 28:31]
    .clock(intsource_3_clock),
    .reset(intsource_3_reset)
  );
  IntSyncSyncCrossingSink_3 intsink ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_clock),
    .reset(intsink_reset)
  );
  IntSyncSyncCrossingSink_4 intsink_1 ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_1_clock),
    .reset(intsink_1_reset)
  );
  IntSyncSyncCrossingSink_5 intsink_2 ( // @[src/main/scala/interrupts/Crossing.scala 99:29]
    .clock(intsink_2_clock),
    .reset(intsink_2_reset)
  );
  ClockSinkDomain bootROMDomainWrapper ( // @[src/main/scala/devices/tilelink/BootROM.scala 74:42]
    .auto_bootrom_in_a_ready(bootROMDomainWrapper_auto_bootrom_in_a_ready),
    .auto_bootrom_in_a_valid(bootROMDomainWrapper_auto_bootrom_in_a_valid),
    .auto_bootrom_in_a_bits_size(bootROMDomainWrapper_auto_bootrom_in_a_bits_size),
    .auto_bootrom_in_a_bits_source(bootROMDomainWrapper_auto_bootrom_in_a_bits_source),
    .auto_bootrom_in_a_bits_address(bootROMDomainWrapper_auto_bootrom_in_a_bits_address),
    .auto_bootrom_in_d_ready(bootROMDomainWrapper_auto_bootrom_in_d_ready),
    .auto_bootrom_in_d_valid(bootROMDomainWrapper_auto_bootrom_in_d_valid),
    .auto_bootrom_in_d_bits_size(bootROMDomainWrapper_auto_bootrom_in_d_bits_size),
    .auto_bootrom_in_d_bits_source(bootROMDomainWrapper_auto_bootrom_in_d_bits_source),
    .auto_bootrom_in_d_bits_data(bootROMDomainWrapper_auto_bootrom_in_d_bits_data),
    .auto_clock_in_clock(bootROMDomainWrapper_auto_clock_in_clock),
    .auto_clock_in_reset(bootROMDomainWrapper_auto_clock_in_reset),
    .clock(bootROMDomainWrapper_clock),
    .reset(bootROMDomainWrapper_reset)
  );
  assign mem_axi4_0_aw_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_aw_bits_id =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_aw_bits_addr =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_aw_bits_len =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_aw_bits_size =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_aw_bits_burst =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_w_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_w_bits_data =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_w_bits_strb =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_w_bits_last =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_b_ready = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_valid = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_bits_id =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_bits_addr =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_bits_len =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_bits_size =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_ar_bits_burst =
    subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign mem_axi4_0_r_ready = subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign ibus_auto_clock_in_clock = subsystem_sbus_auto_fixedClockNode_out_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign ibus_auto_clock_in_reset = subsystem_sbus_auto_fixedClockNode_out_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign dummyClockGroupSourceNode_clock = clock;
  assign dummyClockGroupSourceNode_reset = reset;
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_valid =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data =
    tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_ready =
    tile_prci_domain_auto_tl_master_clock_xing_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_valid =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data =
    tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_ready =
    tile_prci_domain_auto_tl_master_clock_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_valid =
    tile_prci_domain_auto_tl_master_clock_xing_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink =
    tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready =
    subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid =
    subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param =
    subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address =
    subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready =
    subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt =
    subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready =
    subsystem_cbus_auto_bus_xing_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid =
    subsystem_cbus_auto_bus_xing_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode =
    subsystem_cbus_auto_bus_xing_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param =
    subsystem_cbus_auto_bus_xing_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size =
    subsystem_cbus_auto_bus_xing_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source =
    subsystem_cbus_auto_bus_xing_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink =
    subsystem_cbus_auto_bus_xing_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied =
    subsystem_cbus_auto_bus_xing_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data =
    subsystem_cbus_auto_bus_xing_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt =
    subsystem_cbus_auto_bus_xing_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_sbus_auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset =
    dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock =
    subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_pbus_auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset =
    subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_fbus_auto_subsystem_fbus_clock_groups_in_member_subsystem_fbus_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_ready = bootROMDomainWrapper_auto_bootrom_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_valid = bootROMDomainWrapper_auto_bootrom_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_size =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_source =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_bits_data =
    bootROMDomainWrapper_auto_bootrom_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_a_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_size =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_source =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_address =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_a_bits_mask =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_cbus_auto_bus_xing_in_d_ready =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready = mem_axi4_0_aw_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready = mem_axi4_0_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid = mem_axi4_0_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id = mem_axi4_0_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp =
    mem_axi4_0_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready = mem_axi4_0_ar_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid = mem_axi4_0_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id = mem_axi4_0_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data =
    mem_axi4_0_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp =
    mem_axi4_0_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last =
    mem_axi4_0_r_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 1715:56]
  assign subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock =
    subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset =
    subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_valid =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_opcode =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_size =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_source =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_address =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_mask =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_a_bits_data =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_mbus_auto_bus_xing_in_d_ready =
    subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready =
    subsystem_mbus_auto_bus_xing_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid =
    subsystem_mbus_auto_bus_xing_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode =
    subsystem_mbus_auto_bus_xing_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size =
    subsystem_mbus_auto_bus_xing_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source =
    subsystem_mbus_auto_bus_xing_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied =
    subsystem_mbus_auto_bus_xing_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data =
    subsystem_mbus_auto_bus_xing_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt =
    subsystem_mbus_auto_bus_xing_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_opcode =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_param =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_size =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_source =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_address =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_mask =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_a_bits_data =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_b_ready =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_opcode =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_param =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_size =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_source =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_address =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_c_bits_data =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_d_ready =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_e_valid =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_coherent_jbar_in_e_bits_sink =
    subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset =
    subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_prci_domain_auto_tile_reset_domain_tile_hartid_in = tileHartIdNexusNode_auto_out; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_a_ready =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_b_valid =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_param =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_b_bits_address =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_c_ready =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_valid =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_opcode =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_param =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_size =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_source =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_sink =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_denied =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_data =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tl_master_clock_xing_out_d_bits_corrupt =
    subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign tile_prci_domain_auto_tap_clock_in_clock = subsystem_sbus_auto_fixedClockNode_out_1_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign tile_prci_domain_auto_tap_clock_in_reset = subsystem_sbus_auto_fixedClockNode_out_1_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_1_clock = clock;
  assign xbar_1_reset = reset;
  assign xbar_2_clock = clock;
  assign xbar_2_reset = reset;
  assign tileHartIdNexusNode_clock = clock;
  assign tileHartIdNexusNode_reset = reset;
  assign broadcast_clock = clock;
  assign broadcast_reset = reset;
  assign xbar_3_clock = clock;
  assign xbar_3_reset = reset;
  assign intsource_clock = clock;
  assign intsource_reset = reset;
  assign null_int_source_clock = clock;
  assign null_int_source_reset = reset;
  assign intsource_1_clock = clock;
  assign intsource_1_reset = reset;
  assign null_int_source_1_clock = clock;
  assign null_int_source_1_reset = reset;
  assign intsource_2_clock = clock;
  assign intsource_2_reset = reset;
  assign intsource_3_clock = clock;
  assign intsource_3_reset = reset;
  assign intsink_clock = clock;
  assign intsink_reset = reset;
  assign intsink_1_clock = clock;
  assign intsink_1_reset = reset;
  assign intsink_2_clock = clock;
  assign intsink_2_reset = reset;
  assign bootROMDomainWrapper_auto_bootrom_in_a_valid = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_size =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_source =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_bootrom_in_a_bits_address =
    subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_bootrom_in_d_ready = subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_clock_in_clock = subsystem_cbus_auto_fixedClockNode_out_clock; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign bootROMDomainWrapper_auto_clock_in_reset = subsystem_cbus_auto_fixedClockNode_out_reset; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
endmodule
module DifftestMem2P(
  input         clock,
  input         reset,
  input         read_valid, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input  [63:0] read_index, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  output [63:0] read_data_0, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input         write_valid, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_index, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_data_0, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_mask_0 // @[difftest/src/main/scala/common/Mem.scala 204:17]
);
  wire  helper_0_r_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_w_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_mask; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_clock; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  _T_1 = ~reset; // @[difftest/src/main/scala/common/Mem.scala 214:16]
  wire [64:0] _T_3 = read_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 215:26]
  wire [65:0] _T_4 = {{1'd0}, _T_3}; // @[difftest/src/main/scala/common/Mem.scala 215:39]
  wire [64:0] _T_9 = write_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 223:27]
  wire [65:0] _T_10 = {{1'd0}, _T_9}; // @[difftest/src/main/scala/common/Mem.scala 223:40]
  MemRWHelper helper_0 ( // @[difftest/src/main/scala/common/Mem.scala 197:49]
    .r_enable(helper_0_r_enable),
    .r_index(helper_0_r_index),
    .r_data(helper_0_r_data),
    .w_enable(helper_0_w_enable),
    .w_index(helper_0_w_index),
    .w_data(helper_0_w_data),
    .w_mask(helper_0_w_mask),
    .clock(helper_0_clock)
  );
  assign read_data_0 = helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 211:13]
  assign helper_0_r_enable = ~reset & read_valid; // @[difftest/src/main/scala/common/Mem.scala 214:30]
  assign helper_0_r_index = _T_4[63:0]; // @[difftest/src/main/scala/common/Mem.scala 102:13]
  assign helper_0_w_enable = _T_1 & write_valid; // @[difftest/src/main/scala/common/Mem.scala 222:30]
  assign helper_0_w_index = _T_10[63:0]; // @[difftest/src/main/scala/common/Mem.scala 150:13]
  assign helper_0_w_data = write_data_0; // @[difftest/src/main/scala/common/Mem.scala 151:12]
  assign helper_0_w_mask = write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 152:12]
  assign helper_0_clock = clock; // @[difftest/src/main/scala/common/Mem.scala 220:13]
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_echo_real_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  mem_clock; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire  mem_reset; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire  mem_read_valid; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [63:0] mem_read_index; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [63:0] mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire  mem_write_valid; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [63:0] mem_write_index; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [63:0] mem_write_data_0; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [63:0] mem_write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 323:36]
  wire [6:0] r_addr_lo_lo = {auto_in_ar_bits_addr[9],auto_in_ar_bits_addr[8],auto_in_ar_bits_addr[7],
    auto_in_ar_bits_addr[6],auto_in_ar_bits_addr[5],auto_in_ar_bits_addr[4],auto_in_ar_bits_addr[3]}; // @[src/main/scala/amba/axi4/SRAM.scala 67:21]
  wire [13:0] r_addr_lo = {auto_in_ar_bits_addr[16],auto_in_ar_bits_addr[15],auto_in_ar_bits_addr[14],
    auto_in_ar_bits_addr[13],auto_in_ar_bits_addr[12],auto_in_ar_bits_addr[11],auto_in_ar_bits_addr[10],r_addr_lo_lo}; // @[src/main/scala/amba/axi4/SRAM.scala 67:21]
  wire [6:0] r_addr_hi_lo = {auto_in_ar_bits_addr[23],auto_in_ar_bits_addr[22],auto_in_ar_bits_addr[21],
    auto_in_ar_bits_addr[20],auto_in_ar_bits_addr[19],auto_in_ar_bits_addr[18],auto_in_ar_bits_addr[17]}; // @[src/main/scala/amba/axi4/SRAM.scala 67:21]
  wire [27:0] r_addr = {auto_in_ar_bits_addr[30],auto_in_ar_bits_addr[29],auto_in_ar_bits_addr[28],auto_in_ar_bits_addr[
    27],auto_in_ar_bits_addr[26],auto_in_ar_bits_addr[25],auto_in_ar_bits_addr[24],r_addr_hi_lo,r_addr_lo}; // @[src/main/scala/amba/axi4/SRAM.scala 67:21]
  wire [6:0] w_addr_lo_lo = {auto_in_aw_bits_addr[9],auto_in_aw_bits_addr[8],auto_in_aw_bits_addr[7],
    auto_in_aw_bits_addr[6],auto_in_aw_bits_addr[5],auto_in_aw_bits_addr[4],auto_in_aw_bits_addr[3]}; // @[src/main/scala/amba/axi4/SRAM.scala 68:21]
  wire [13:0] w_addr_lo = {auto_in_aw_bits_addr[16],auto_in_aw_bits_addr[15],auto_in_aw_bits_addr[14],
    auto_in_aw_bits_addr[13],auto_in_aw_bits_addr[12],auto_in_aw_bits_addr[11],auto_in_aw_bits_addr[10],w_addr_lo_lo}; // @[src/main/scala/amba/axi4/SRAM.scala 68:21]
  wire [6:0] w_addr_hi_lo = {auto_in_aw_bits_addr[23],auto_in_aw_bits_addr[22],auto_in_aw_bits_addr[21],
    auto_in_aw_bits_addr[20],auto_in_aw_bits_addr[19],auto_in_aw_bits_addr[18],auto_in_aw_bits_addr[17]}; // @[src/main/scala/amba/axi4/SRAM.scala 68:21]
  wire [27:0] w_addr = {auto_in_aw_bits_addr[30],auto_in_aw_bits_addr[29],auto_in_aw_bits_addr[28],auto_in_aw_bits_addr[
    27],auto_in_aw_bits_addr[26],auto_in_aw_bits_addr[25],auto_in_aw_bits_addr[24],w_addr_hi_lo,w_addr_lo}; // @[src/main/scala/amba/axi4/SRAM.scala 68:21]
  wire [31:0] _r_sel0_T = auto_in_ar_bits_addr ^ 32'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [32:0] _r_sel0_T_1 = {1'b0,$signed(_r_sel0_T)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [32:0] _r_sel0_T_3 = $signed(_r_sel0_T_1) & -33'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire [31:0] _w_sel0_T = auto_in_aw_bits_addr ^ 32'h80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:31]
  wire [32:0] _w_sel0_T_1 = {1'b0,$signed(_w_sel0_T)}; // @[src/main/scala/diplomacy/Parameters.scala 137:41]
  wire [32:0] _w_sel0_T_3 = $signed(_w_sel0_T_1) & -33'sh80000000; // @[src/main/scala/diplomacy/Parameters.scala 137:46]
  wire  w_sel0 = $signed(_w_sel0_T_3) == 33'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
  reg  w_full; // @[src/main/scala/amba/axi4/SRAM.scala 72:25]
  reg [3:0] w_id; // @[src/main/scala/amba/axi4/SRAM.scala 73:21]
  reg  w_echo_real_last; // @[src/main/scala/amba/axi4/SRAM.scala 74:21]
  reg  r_sel1; // @[src/main/scala/amba/axi4/SRAM.scala 75:25]
  reg  w_sel1; // @[src/main/scala/amba/axi4/SRAM.scala 76:25]
  wire  _T = auto_in_b_ready & w_full; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1256_clock;
  wire  line_1256_reset;
  wire  line_1256_valid;
  reg  line_1256_valid_reg;
  wire  _GEN_8 = _T ? 1'h0 : w_full; // @[src/main/scala/amba/axi4/SRAM.scala 78:23 72:25 78:32]
  wire  _nodeIn_aw_ready_T_1 = auto_in_b_ready | ~w_full; // @[src/main/scala/amba/axi4/SRAM.scala 94:47]
  wire  nodeIn_aw_ready = auto_in_w_valid & (auto_in_b_ready | ~w_full); // @[src/main/scala/amba/axi4/SRAM.scala 94:32]
  wire  _T_1 = nodeIn_aw_ready & auto_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1257_clock;
  wire  line_1257_reset;
  wire  line_1257_valid;
  reg  line_1257_valid_reg;
  wire  _GEN_9 = _T_1 | _GEN_8; // @[src/main/scala/amba/axi4/SRAM.scala 79:{23,32}]
  wire  line_1258_clock;
  wire  line_1258_reset;
  wire  line_1258_valid;
  reg  line_1258_valid_reg;
  wire [7:0] wdata_0 = auto_in_w_bits_data[7:0]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_1 = auto_in_w_bits_data[15:8]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_2 = auto_in_w_bits_data[23:16]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_3 = auto_in_w_bits_data[31:24]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_4 = auto_in_w_bits_data[39:32]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_5 = auto_in_w_bits_data[47:40]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_6 = auto_in_w_bits_data[55:48]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire [7:0] wdata_7 = auto_in_w_bits_data[63:56]; // @[src/main/scala/amba/axi4/SRAM.scala 87:66]
  wire  _T_4 = _T_1 & w_sel0; // @[src/main/scala/amba/axi4/SRAM.scala 88:22]
  wire  line_1259_clock;
  wire  line_1259_reset;
  wire  line_1259_valid;
  reg  line_1259_valid_reg;
  wire [31:0] lo = {wdata_3,wdata_2,wdata_1,wdata_0}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [31:0] hi = {wdata_7,wdata_6,wdata_5,wdata_4}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [7:0] _T_15 = auto_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_16 = auto_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_17 = auto_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_18 = auto_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_19 = auto_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_20 = auto_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_21 = auto_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _T_22 = auto_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [31:0] lo_1 = {_T_18,_T_17,_T_16,_T_15}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  wire [31:0] hi_1 = {_T_22,_T_21,_T_20,_T_19}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  reg  r_full; // @[src/main/scala/amba/axi4/SRAM.scala 101:25]
  reg [3:0] r_id; // @[src/main/scala/amba/axi4/SRAM.scala 102:21]
  reg  r_echo_real_last; // @[src/main/scala/amba/axi4/SRAM.scala 103:21]
  wire  _T_25 = auto_in_r_ready & r_full; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1260_clock;
  wire  line_1260_reset;
  wire  line_1260_valid;
  reg  line_1260_valid_reg;
  wire  _GEN_17 = _T_25 ? 1'h0 : r_full; // @[src/main/scala/amba/axi4/SRAM.scala 105:23 101:25 105:32]
  wire  nodeIn_ar_ready = auto_in_r_ready | ~r_full; // @[src/main/scala/amba/axi4/SRAM.scala 119:31]
  wire  _T_26 = nodeIn_ar_ready & auto_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1261_clock;
  wire  line_1261_reset;
  wire  line_1261_valid;
  reg  line_1261_valid_reg;
  wire  _GEN_18 = _T_26 | _GEN_17; // @[src/main/scala/amba/axi4/SRAM.scala 106:{23,32}]
  wire  line_1262_clock;
  wire  line_1262_reset;
  wire  line_1262_valid;
  reg  line_1262_valid_reg;
  reg  rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  reg  rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  reg [63:0] rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire  line_1263_clock;
  wire  line_1263_reset;
  wire  line_1263_valid;
  reg  line_1263_valid_reg;
  wire [63:0] _rdata_T_0 = rdata_REG ? mem_read_data_0 : rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:8]
  wire [7:0] rdata_0 = _rdata_T_0[7:0]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_1 = _rdata_T_0[15:8]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_2 = _rdata_T_0[23:16]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_3 = _rdata_T_0[31:24]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_4 = _rdata_T_0[39:32]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_5 = _rdata_T_0[47:40]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_6 = _rdata_T_0[55:48]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [7:0] rdata_7 = _rdata_T_0[63:56]; // @[difftest/src/main/scala/common/Mem.scala 238:76]
  wire [31:0] nodeIn_r_bits_data_lo = {rdata_3,rdata_2,rdata_1,rdata_0}; // @[src/main/scala/amba/axi4/SRAM.scala 123:26]
  wire [31:0] nodeIn_r_bits_data_hi = {rdata_7,rdata_6,rdata_5,rdata_4}; // @[src/main/scala/amba/axi4/SRAM.scala 123:26]
  DifftestMem2P mem ( // @[difftest/src/main/scala/common/Mem.scala 323:36]
    .clock(mem_clock),
    .reset(mem_reset),
    .read_valid(mem_read_valid),
    .read_index(mem_read_index),
    .read_data_0(mem_read_data_0),
    .write_valid(mem_write_valid),
    .write_index(mem_write_index),
    .write_data_0(mem_write_data_0),
    .write_mask_0(mem_write_mask_0)
  );
  GEN_w1_line #(.COVER_INDEX(1256)) line_1256 (
    .clock(line_1256_clock),
    .reset(line_1256_reset),
    .valid(line_1256_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1257)) line_1257 (
    .clock(line_1257_clock),
    .reset(line_1257_reset),
    .valid(line_1257_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1258)) line_1258 (
    .clock(line_1258_clock),
    .reset(line_1258_reset),
    .valid(line_1258_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1259)) line_1259 (
    .clock(line_1259_clock),
    .reset(line_1259_reset),
    .valid(line_1259_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1260)) line_1260 (
    .clock(line_1260_clock),
    .reset(line_1260_reset),
    .valid(line_1260_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1261)) line_1261 (
    .clock(line_1261_clock),
    .reset(line_1261_reset),
    .valid(line_1261_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1262)) line_1262 (
    .clock(line_1262_clock),
    .reset(line_1262_reset),
    .valid(line_1262_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1263)) line_1263 (
    .clock(line_1263_clock),
    .reset(line_1263_reset),
    .valid(line_1263_valid)
  );
  assign line_1256_clock = clock;
  assign line_1256_reset = reset;
  assign line_1256_valid = _T ^ line_1256_valid_reg;
  assign line_1257_clock = clock;
  assign line_1257_reset = reset;
  assign line_1257_valid = _T_1 ^ line_1257_valid_reg;
  assign line_1258_clock = clock;
  assign line_1258_reset = reset;
  assign line_1258_valid = _T_1 ^ line_1258_valid_reg;
  assign line_1259_clock = clock;
  assign line_1259_reset = reset;
  assign line_1259_valid = _T_4 ^ line_1259_valid_reg;
  assign line_1260_clock = clock;
  assign line_1260_reset = reset;
  assign line_1260_valid = _T_25 ^ line_1260_valid_reg;
  assign line_1261_clock = clock;
  assign line_1261_reset = reset;
  assign line_1261_valid = _T_26 ^ line_1261_valid_reg;
  assign line_1262_clock = clock;
  assign line_1262_reset = reset;
  assign line_1262_valid = _T_26 ^ line_1262_valid_reg;
  assign line_1263_clock = clock;
  assign line_1263_reset = reset;
  assign line_1263_valid = rdata_REG_1 ^ line_1263_valid_reg;
  assign auto_in_aw_ready = auto_in_w_valid & (auto_in_b_ready | ~w_full); // @[src/main/scala/amba/axi4/SRAM.scala 94:32]
  assign auto_in_w_ready = auto_in_aw_valid & _nodeIn_aw_ready_T_1; // @[src/main/scala/amba/axi4/SRAM.scala 95:32]
  assign auto_in_b_valid = w_full; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/amba/axi4/SRAM.scala 93:17]
  assign auto_in_b_bits_id = w_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/amba/axi4/SRAM.scala 97:20]
  assign auto_in_b_bits_resp = w_sel1 ? 2'h0 : 2'h3; // @[src/main/scala/amba/axi4/SRAM.scala 98:26]
  assign auto_in_b_bits_echo_real_last = w_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/amba/axi4/SRAM.scala 99:20]
  assign auto_in_ar_ready = auto_in_r_ready | ~r_full; // @[src/main/scala/amba/axi4/SRAM.scala 119:31]
  assign auto_in_r_valid = r_full; // @[src/main/scala/amba/axi4/SRAM.scala 118:17 src/main/scala/diplomacy/Nodes.scala 1214:17]
  assign auto_in_r_bits_id = r_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/amba/axi4/SRAM.scala 121:20]
  assign auto_in_r_bits_data = {nodeIn_r_bits_data_hi,nodeIn_r_bits_data_lo}; // @[src/main/scala/amba/axi4/SRAM.scala 123:26]
  assign auto_in_r_bits_resp = r_sel1 ? 2'h0 : 2'h3; // @[src/main/scala/amba/axi4/SRAM.scala 122:26]
  assign auto_in_r_bits_echo_real_last = r_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/amba/axi4/SRAM.scala 124:20]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_read_valid = nodeIn_ar_ready & auto_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  assign mem_read_index = {{36'd0}, r_addr}; // @[difftest/src/main/scala/common/Mem.scala 237:16]
  assign mem_write_valid = _T_1 & w_sel0; // @[src/main/scala/amba/axi4/SRAM.scala 88:22]
  assign mem_write_index = {{36'd0}, w_addr};
  assign mem_write_data_0 = {hi,lo}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  assign mem_write_mask_0 = {hi_1,lo_1}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/amba/axi4/SRAM.scala 72:25]
      w_full <= 1'h0; // @[src/main/scala/amba/axi4/SRAM.scala 72:25]
    end else begin
      w_full <= _GEN_9;
    end
    if (_T_1) begin // @[src/main/scala/amba/axi4/SRAM.scala 81:23]
      w_id <= auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/SRAM.scala 82:12]
    end
    if (_T_1) begin // @[src/main/scala/amba/axi4/SRAM.scala 81:23]
      w_echo_real_last <= auto_in_aw_bits_echo_real_last; // @[src/main/scala/amba/axi4/SRAM.scala 84:14]
    end
    r_sel1 <= $signed(_r_sel0_T_3) == 33'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
    w_sel1 <= $signed(_w_sel0_T_3) == 33'sh0; // @[src/main/scala/diplomacy/Parameters.scala 137:59]
    line_1256_valid_reg <= _T;
    line_1257_valid_reg <= _T_1;
    line_1258_valid_reg <= _T_1;
    line_1259_valid_reg <= _T_4;
    if (reset) begin // @[src/main/scala/amba/axi4/SRAM.scala 101:25]
      r_full <= 1'h0; // @[src/main/scala/amba/axi4/SRAM.scala 101:25]
    end else begin
      r_full <= _GEN_18;
    end
    if (_T_26) begin // @[src/main/scala/amba/axi4/SRAM.scala 108:23]
      r_id <= auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/SRAM.scala 109:12]
    end
    if (_T_26) begin // @[src/main/scala/amba/axi4/SRAM.scala 108:23]
      r_echo_real_last <= auto_in_ar_bits_echo_real_last; // @[src/main/scala/amba/axi4/SRAM.scala 111:14]
    end
    line_1260_valid_reg <= _T_25;
    line_1261_valid_reg <= _T_26;
    line_1262_valid_reg <= _T_26;
    rdata_REG <= nodeIn_ar_ready & auto_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    rdata_REG_1 <= nodeIn_ar_ready & auto_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    if (rdata_REG_1) begin // @[difftest/src/main/scala/common/Mem.scala 238:42]
      rdata_r_0 <= mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    line_1263_valid_reg <= rdata_REG_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  w_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  w_id = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  w_echo_real_last = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_sel1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  w_sel1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1256_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1257_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1258_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1259_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_full = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_id = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  r_echo_real_last = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1260_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1261_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1262_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  rdata_REG = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  rdata_REG_1 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  rdata_r_0 = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  line_1263_valid_reg = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_45(
  input   clock,
  input   reset
);
endmodule
module Queue_46(
  input   clock,
  input   reset
);
endmodule
module AXI4Xbar(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [2:0]  auto_out_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_out_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  awIn_0_clock; // @[src/main/scala/amba/axi4/Xbar.scala 70:47]
  wire  awIn_0_reset; // @[src/main/scala/amba/axi4/Xbar.scala 70:47]
  wire  awOut_0_clock; // @[src/main/scala/amba/axi4/Xbar.scala 71:47]
  wire  awOut_0_reset; // @[src/main/scala/amba/axi4/Xbar.scala 71:47]
  wire  _awOut_0_io_enq_bits_T_1 = ~auto_in_aw_valid; // @[src/main/scala/amba/axi4/Xbar.scala 275:60]
  wire  _awOut_0_io_enq_bits_T_4 = ~reset; // @[src/main/scala/amba/axi4/Xbar.scala 275:11]
  wire  line_1264_clock;
  wire  line_1264_reset;
  wire  line_1264_valid;
  reg  line_1264_valid_reg;
  wire  line_1265_clock;
  wire  line_1265_reset;
  wire  line_1265_valid;
  reg  line_1265_valid_reg;
  wire  _awOut_0_io_enq_bits_T_10 = ~(_awOut_0_io_enq_bits_T_1 | auto_in_aw_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
  wire  line_1266_clock;
  wire  line_1266_reset;
  wire  line_1266_valid;
  reg  line_1266_valid_reg;
  wire  line_1267_clock;
  wire  line_1267_reset;
  wire  line_1267_valid;
  reg  line_1267_valid_reg;
  wire  _awOut_0_io_enq_bits_T_11 = auto_out_aw_ready & auto_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1268_clock;
  wire  line_1268_reset;
  wire  line_1268_valid;
  reg  line_1268_valid_reg;
  wire  _T_1 = ~auto_in_ar_valid; // @[src/main/scala/amba/axi4/Xbar.scala 275:60]
  wire  line_1269_clock;
  wire  line_1269_reset;
  wire  line_1269_valid;
  reg  line_1269_valid_reg;
  wire  line_1270_clock;
  wire  line_1270_reset;
  wire  line_1270_valid;
  reg  line_1270_valid_reg;
  wire  _T_10 = ~(_T_1 | auto_in_ar_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
  wire  line_1271_clock;
  wire  line_1271_reset;
  wire  line_1271_valid;
  reg  line_1271_valid_reg;
  wire  line_1272_clock;
  wire  line_1272_reset;
  wire  line_1272_valid;
  reg  line_1272_valid_reg;
  wire  _T_11 = auto_out_ar_ready & auto_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1273_clock;
  wire  line_1273_reset;
  wire  line_1273_valid;
  reg  line_1273_valid_reg;
  wire  _T_13 = ~auto_out_r_valid; // @[src/main/scala/amba/axi4/Xbar.scala 275:60]
  wire  line_1274_clock;
  wire  line_1274_reset;
  wire  line_1274_valid;
  reg  line_1274_valid_reg;
  wire  line_1275_clock;
  wire  line_1275_reset;
  wire  line_1275_valid;
  reg  line_1275_valid_reg;
  wire  _T_22 = ~(_T_13 | auto_out_r_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
  wire  line_1276_clock;
  wire  line_1276_reset;
  wire  line_1276_valid;
  reg  line_1276_valid_reg;
  wire  line_1277_clock;
  wire  line_1277_reset;
  wire  line_1277_valid;
  reg  line_1277_valid_reg;
  wire  _T_23 = auto_in_r_ready & auto_out_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1278_clock;
  wire  line_1278_reset;
  wire  line_1278_valid;
  reg  line_1278_valid_reg;
  wire  _T_25 = ~auto_out_b_valid; // @[src/main/scala/amba/axi4/Xbar.scala 275:60]
  wire  line_1279_clock;
  wire  line_1279_reset;
  wire  line_1279_valid;
  reg  line_1279_valid_reg;
  wire  line_1280_clock;
  wire  line_1280_reset;
  wire  line_1280_valid;
  reg  line_1280_valid_reg;
  wire  _T_34 = ~(_T_25 | auto_out_b_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
  wire  line_1281_clock;
  wire  line_1281_reset;
  wire  line_1281_valid;
  reg  line_1281_valid_reg;
  wire  line_1282_clock;
  wire  line_1282_reset;
  wire  line_1282_valid;
  reg  line_1282_valid_reg;
  wire  _T_35 = auto_in_b_ready & auto_out_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1283_clock;
  wire  line_1283_reset;
  wire  line_1283_valid;
  reg  line_1283_valid_reg;
  Queue_45 awIn_0 ( // @[src/main/scala/amba/axi4/Xbar.scala 70:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset)
  );
  Queue_46 awOut_0 ( // @[src/main/scala/amba/axi4/Xbar.scala 71:47]
    .clock(awOut_0_clock),
    .reset(awOut_0_reset)
  );
  GEN_w1_line #(.COVER_INDEX(1264)) line_1264 (
    .clock(line_1264_clock),
    .reset(line_1264_reset),
    .valid(line_1264_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1265)) line_1265 (
    .clock(line_1265_clock),
    .reset(line_1265_reset),
    .valid(line_1265_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1266)) line_1266 (
    .clock(line_1266_clock),
    .reset(line_1266_reset),
    .valid(line_1266_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1267)) line_1267 (
    .clock(line_1267_clock),
    .reset(line_1267_reset),
    .valid(line_1267_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1268)) line_1268 (
    .clock(line_1268_clock),
    .reset(line_1268_reset),
    .valid(line_1268_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1269)) line_1269 (
    .clock(line_1269_clock),
    .reset(line_1269_reset),
    .valid(line_1269_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1270)) line_1270 (
    .clock(line_1270_clock),
    .reset(line_1270_reset),
    .valid(line_1270_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1271)) line_1271 (
    .clock(line_1271_clock),
    .reset(line_1271_reset),
    .valid(line_1271_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1272)) line_1272 (
    .clock(line_1272_clock),
    .reset(line_1272_reset),
    .valid(line_1272_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1273)) line_1273 (
    .clock(line_1273_clock),
    .reset(line_1273_reset),
    .valid(line_1273_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1274)) line_1274 (
    .clock(line_1274_clock),
    .reset(line_1274_reset),
    .valid(line_1274_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1275)) line_1275 (
    .clock(line_1275_clock),
    .reset(line_1275_reset),
    .valid(line_1275_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1276)) line_1276 (
    .clock(line_1276_clock),
    .reset(line_1276_reset),
    .valid(line_1276_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1277)) line_1277 (
    .clock(line_1277_clock),
    .reset(line_1277_reset),
    .valid(line_1277_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1278)) line_1278 (
    .clock(line_1278_clock),
    .reset(line_1278_reset),
    .valid(line_1278_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1279)) line_1279 (
    .clock(line_1279_clock),
    .reset(line_1279_reset),
    .valid(line_1279_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1280)) line_1280 (
    .clock(line_1280_clock),
    .reset(line_1280_reset),
    .valid(line_1280_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1281)) line_1281 (
    .clock(line_1281_clock),
    .reset(line_1281_reset),
    .valid(line_1281_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1282)) line_1282 (
    .clock(line_1282_clock),
    .reset(line_1282_reset),
    .valid(line_1282_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1283)) line_1283 (
    .clock(line_1283_clock),
    .reset(line_1283_reset),
    .valid(line_1283_valid)
  );
  assign line_1264_clock = clock;
  assign line_1264_reset = reset;
  assign line_1264_valid = _awOut_0_io_enq_bits_T_4 ^ line_1264_valid_reg;
  assign line_1265_clock = clock;
  assign line_1265_reset = reset;
  assign line_1265_valid = _awOut_0_io_enq_bits_T_4 ^ line_1265_valid_reg;
  assign line_1266_clock = clock;
  assign line_1266_reset = reset;
  assign line_1266_valid = _awOut_0_io_enq_bits_T_10 ^ line_1266_valid_reg;
  assign line_1267_clock = clock;
  assign line_1267_reset = reset;
  assign line_1267_valid = auto_in_aw_valid ^ line_1267_valid_reg;
  assign line_1268_clock = clock;
  assign line_1268_reset = reset;
  assign line_1268_valid = _awOut_0_io_enq_bits_T_11 ^ line_1268_valid_reg;
  assign line_1269_clock = clock;
  assign line_1269_reset = reset;
  assign line_1269_valid = _awOut_0_io_enq_bits_T_4 ^ line_1269_valid_reg;
  assign line_1270_clock = clock;
  assign line_1270_reset = reset;
  assign line_1270_valid = _awOut_0_io_enq_bits_T_4 ^ line_1270_valid_reg;
  assign line_1271_clock = clock;
  assign line_1271_reset = reset;
  assign line_1271_valid = _T_10 ^ line_1271_valid_reg;
  assign line_1272_clock = clock;
  assign line_1272_reset = reset;
  assign line_1272_valid = auto_in_ar_valid ^ line_1272_valid_reg;
  assign line_1273_clock = clock;
  assign line_1273_reset = reset;
  assign line_1273_valid = _T_11 ^ line_1273_valid_reg;
  assign line_1274_clock = clock;
  assign line_1274_reset = reset;
  assign line_1274_valid = _awOut_0_io_enq_bits_T_4 ^ line_1274_valid_reg;
  assign line_1275_clock = clock;
  assign line_1275_reset = reset;
  assign line_1275_valid = _awOut_0_io_enq_bits_T_4 ^ line_1275_valid_reg;
  assign line_1276_clock = clock;
  assign line_1276_reset = reset;
  assign line_1276_valid = _T_22 ^ line_1276_valid_reg;
  assign line_1277_clock = clock;
  assign line_1277_reset = reset;
  assign line_1277_valid = auto_out_r_valid ^ line_1277_valid_reg;
  assign line_1278_clock = clock;
  assign line_1278_reset = reset;
  assign line_1278_valid = _T_23 ^ line_1278_valid_reg;
  assign line_1279_clock = clock;
  assign line_1279_reset = reset;
  assign line_1279_valid = _awOut_0_io_enq_bits_T_4 ^ line_1279_valid_reg;
  assign line_1280_clock = clock;
  assign line_1280_reset = reset;
  assign line_1280_valid = _awOut_0_io_enq_bits_T_4 ^ line_1280_valid_reg;
  assign line_1281_clock = clock;
  assign line_1281_reset = reset;
  assign line_1281_valid = _T_34 ^ line_1281_valid_reg;
  assign line_1282_clock = clock;
  assign line_1282_reset = reset;
  assign line_1282_valid = auto_out_b_valid ^ line_1282_valid_reg;
  assign line_1283_clock = clock;
  assign line_1283_reset = reset;
  assign line_1283_valid = _T_35 ^ line_1283_valid_reg;
  assign auto_in_aw_ready = auto_out_aw_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_w_ready = auto_out_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_valid = auto_out_b_valid; // @[src/main/scala/amba/axi4/Xbar.scala 297:22]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 91:65]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_valid = auto_out_r_valid; // @[src/main/scala/amba/axi4/Xbar.scala 297:22]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 91:65]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[src/main/scala/amba/axi4/Xbar.scala 297:22]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 94:47]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_len = auto_in_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_valid = auto_in_w_valid; // @[src/main/scala/amba/axi4/Xbar.scala 241:40]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_b_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[src/main/scala/amba/axi4/Xbar.scala 297:22]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 95:47]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_len = auto_in_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign auto_out_r_ready = auto_in_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awOut_0_clock = clock;
  assign awOut_0_reset = reset;
  always @(posedge clock) begin
    line_1264_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1265_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1266_valid_reg <= _awOut_0_io_enq_bits_T_10;
    line_1267_valid_reg <= auto_in_aw_valid;
    line_1268_valid_reg <= _awOut_0_io_enq_bits_T_11;
    line_1269_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1270_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1271_valid_reg <= _T_10;
    line_1272_valid_reg <= auto_in_ar_valid;
    line_1273_valid_reg <= _T_11;
    line_1274_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1275_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1276_valid_reg <= _T_22;
    line_1277_valid_reg <= auto_out_r_valid;
    line_1278_valid_reg <= _T_23;
    line_1279_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1280_valid_reg <= _awOut_0_io_enq_bits_T_4;
    line_1281_valid_reg <= _T_34;
    line_1282_valid_reg <= auto_out_b_valid;
    line_1283_valid_reg <= _T_35;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_awOut_0_io_enq_bits_T_1 | auto_in_aw_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:277 assert (!anyValid || winner.reduce(_||_))\n"); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_1 | auto_in_ar_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:277 assert (!anyValid || winner.reduce(_||_))\n"); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_13 | auto_out_r_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:277 assert (!anyValid || winner.reduce(_||_))\n"); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_awOut_0_io_enq_bits_T_4 & ~(_T_25 | auto_out_b_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:277 assert (!anyValid || winner.reduce(_||_))\n"); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_1264_valid_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  line_1265_valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  line_1266_valid_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  line_1267_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1268_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1269_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1270_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1271_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1272_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1273_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1274_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  line_1275_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  line_1276_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1277_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1278_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1279_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1280_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1281_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1282_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1283_valid_reg = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/amba/axi4/Xbar.scala 275:11]
    end
    //
    if (_awOut_0_io_enq_bits_T_4) begin
      assert(_awOut_0_io_enq_bits_T_1 | auto_in_aw_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/amba/axi4/Xbar.scala 275:11]
    end
    //
    if (_awOut_0_io_enq_bits_T_4) begin
      assert(_T_1 | auto_in_ar_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/amba/axi4/Xbar.scala 275:11]
    end
    //
    if (_awOut_0_io_enq_bits_T_4) begin
      assert(_T_13 | auto_out_r_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/amba/axi4/Xbar.scala 275:11]
    end
    //
    if (_awOut_0_io_enq_bits_T_4) begin
      assert(_T_25 | auto_out_b_valid); // @[src/main/scala/amba/axi4/Xbar.scala 277:12]
    end
  end
endmodule
module Queue_47(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_echo_real_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_echo_real_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_addr [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_echo_real_last [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1284_clock;
  wire  line_1284_reset;
  wire  line_1284_valid;
  reg  line_1284_valid_reg;
  wire  line_1285_clock;
  wire  line_1285_reset;
  wire  line_1285_valid;
  reg  line_1285_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1286_clock;
  wire  line_1286_reset;
  wire  line_1286_valid;
  reg  line_1286_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1284)) line_1284 (
    .clock(line_1284_clock),
    .reset(line_1284_reset),
    .valid(line_1284_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1285)) line_1285 (
    .clock(line_1285_clock),
    .reset(line_1285_reset),
    .valid(line_1285_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1286)) line_1286 (
    .clock(line_1286_clock),
    .reset(line_1286_reset),
    .valid(line_1286_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_real_last_io_deq_bits_MPORT_data = ram_echo_real_last[ram_echo_real_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_real_last_MPORT_data = io_enq_bits_echo_real_last;
  assign ram_echo_real_last_MPORT_addr = enq_ptr_value;
  assign ram_echo_real_last_MPORT_mask = 1'h1;
  assign ram_echo_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1284_clock = clock;
  assign line_1284_reset = reset;
  assign line_1284_valid = do_enq ^ line_1284_valid_reg;
  assign line_1285_clock = clock;
  assign line_1285_reset = reset;
  assign line_1285_valid = do_deq ^ line_1285_valid_reg;
  assign line_1286_clock = clock;
  assign line_1286_reset = reset;
  assign line_1286_valid = _T ^ line_1286_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_echo_real_last = ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_real_last_MPORT_en & ram_echo_real_last_MPORT_mask) begin
      ram_echo_real_last[ram_echo_real_last_MPORT_addr] <= ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1284_valid_reg <= do_enq;
    line_1285_valid_reg <= do_deq;
    line_1286_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_echo_real_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1284_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1285_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1286_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_48(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_strb // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_strb [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1287_clock;
  wire  line_1287_reset;
  wire  line_1287_valid;
  reg  line_1287_valid_reg;
  wire  line_1288_clock;
  wire  line_1288_reset;
  wire  line_1288_valid;
  reg  line_1288_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1289_clock;
  wire  line_1289_reset;
  wire  line_1289_valid;
  reg  line_1289_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1287)) line_1287 (
    .clock(line_1287_clock),
    .reset(line_1287_reset),
    .valid(line_1287_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1288)) line_1288 (
    .clock(line_1288_clock),
    .reset(line_1288_reset),
    .valid(line_1288_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1289)) line_1289 (
    .clock(line_1289_clock),
    .reset(line_1289_reset),
    .valid(line_1289_valid)
  );
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = enq_ptr_value;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1287_clock = clock;
  assign line_1287_reset = reset;
  assign line_1287_valid = do_enq ^ line_1287_valid_reg;
  assign line_1288_clock = clock;
  assign line_1288_reset = reset;
  assign line_1288_valid = do_deq ^ line_1288_valid_reg;
  assign line_1289_clock = clock;
  assign line_1289_reset = reset;
  assign line_1289_valid = _T ^ line_1289_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_strb = ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1287_valid_reg <= do_enq;
    line_1288_valid_reg <= do_deq;
    line_1289_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1287_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1288_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1289_valid_reg = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_49(
  input        clock,
  input        reset,
  output       io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0] io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0] io_enq_bits_resp, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_enq_bits_echo_real_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input        io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0] io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0] io_deq_bits_resp, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output       io_deq_bits_echo_real_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_resp [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_resp_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_echo_real_last [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1290_clock;
  wire  line_1290_reset;
  wire  line_1290_valid;
  reg  line_1290_valid_reg;
  wire  line_1291_clock;
  wire  line_1291_reset;
  wire  line_1291_valid;
  reg  line_1291_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1292_clock;
  wire  line_1292_reset;
  wire  line_1292_valid;
  reg  line_1292_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1290)) line_1290 (
    .clock(line_1290_clock),
    .reset(line_1290_reset),
    .valid(line_1290_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1291)) line_1291 (
    .clock(line_1291_clock),
    .reset(line_1291_reset),
    .valid(line_1291_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1292)) line_1292 (
    .clock(line_1292_clock),
    .reset(line_1292_reset),
    .valid(line_1292_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_real_last_io_deq_bits_MPORT_data = ram_echo_real_last[ram_echo_real_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_real_last_MPORT_data = io_enq_bits_echo_real_last;
  assign ram_echo_real_last_MPORT_addr = enq_ptr_value;
  assign ram_echo_real_last_MPORT_mask = 1'h1;
  assign ram_echo_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1290_clock = clock;
  assign line_1290_reset = reset;
  assign line_1290_valid = do_enq ^ line_1290_valid_reg;
  assign line_1291_clock = clock;
  assign line_1291_reset = reset;
  assign line_1291_valid = do_deq ^ line_1291_valid_reg;
  assign line_1292_clock = clock;
  assign line_1292_reset = reset;
  assign line_1292_valid = _T ^ line_1292_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_echo_real_last = ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_real_last_MPORT_en & ram_echo_real_last_MPORT_mask) begin
      ram_echo_real_last[ram_echo_real_last_MPORT_addr] <= ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1290_valid_reg <= do_enq;
    line_1291_valid_reg <= do_deq;
    line_1292_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_echo_real_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1290_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1291_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1292_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_50(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_echo_real_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_echo_real_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_addr [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_echo_real_last [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1293_clock;
  wire  line_1293_reset;
  wire  line_1293_valid;
  reg  line_1293_valid_reg;
  wire  line_1294_clock;
  wire  line_1294_reset;
  wire  line_1294_valid;
  reg  line_1294_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1295_clock;
  wire  line_1295_reset;
  wire  line_1295_valid;
  reg  line_1295_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1293)) line_1293 (
    .clock(line_1293_clock),
    .reset(line_1293_reset),
    .valid(line_1293_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1294)) line_1294 (
    .clock(line_1294_clock),
    .reset(line_1294_reset),
    .valid(line_1294_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1295)) line_1295 (
    .clock(line_1295_clock),
    .reset(line_1295_reset),
    .valid(line_1295_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_real_last_io_deq_bits_MPORT_data = ram_echo_real_last[ram_echo_real_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_real_last_MPORT_data = io_enq_bits_echo_real_last;
  assign ram_echo_real_last_MPORT_addr = enq_ptr_value;
  assign ram_echo_real_last_MPORT_mask = 1'h1;
  assign ram_echo_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1293_clock = clock;
  assign line_1293_reset = reset;
  assign line_1293_valid = do_enq ^ line_1293_valid_reg;
  assign line_1294_clock = clock;
  assign line_1294_reset = reset;
  assign line_1294_valid = do_deq ^ line_1294_valid_reg;
  assign line_1295_clock = clock;
  assign line_1295_reset = reset;
  assign line_1295_valid = _T ^ line_1295_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_echo_real_last = ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_real_last_MPORT_en & ram_echo_real_last_MPORT_mask) begin
      ram_echo_real_last[ram_echo_real_last_MPORT_addr] <= ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1293_valid_reg <= do_enq;
    line_1294_valid_reg <= do_deq;
    line_1295_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_echo_real_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enq_ptr_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  deq_ptr_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1293_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1294_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1295_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_51(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_resp, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_echo_real_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_resp, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_echo_real_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [63:0] ram_data [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_resp [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_resp_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_resp_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_resp_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_echo_real_last [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_echo_real_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_last [0:1]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/chisel3/util/Decoupled.scala 283:33]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:25]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 285:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1296_clock;
  wire  line_1296_reset;
  wire  line_1296_valid;
  reg  line_1296_valid_reg;
  wire  line_1297_clock;
  wire  line_1297_reset;
  wire  line_1297_valid;
  reg  line_1297_valid_reg;
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1298_clock;
  wire  line_1298_reset;
  wire  line_1298_valid;
  reg  line_1298_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1296)) line_1296 (
    .clock(line_1296_clock),
    .reset(line_1296_reset),
    .valid(line_1296_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1297)) line_1297 (
    .clock(line_1297_clock),
    .reset(line_1297_reset),
    .valid(line_1297_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1298)) line_1298 (
    .clock(line_1298_clock),
    .reset(line_1298_reset),
    .valid(line_1298_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_resp_io_deq_bits_MPORT_en = 1'h1;
  assign ram_resp_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_resp_io_deq_bits_MPORT_data = ram_resp[ram_resp_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_resp_MPORT_data = io_enq_bits_resp;
  assign ram_resp_MPORT_addr = enq_ptr_value;
  assign ram_resp_MPORT_mask = 1'h1;
  assign ram_resp_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_echo_real_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_echo_real_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_echo_real_last_io_deq_bits_MPORT_data = ram_echo_real_last[ram_echo_real_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_echo_real_last_MPORT_data = io_enq_bits_echo_real_last;
  assign ram_echo_real_last_MPORT_addr = enq_ptr_value;
  assign ram_echo_real_last_MPORT_mask = 1'h1;
  assign ram_echo_real_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_last_MPORT_data = 1'h1;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign line_1296_clock = clock;
  assign line_1296_reset = reset;
  assign line_1296_valid = do_enq ^ line_1296_valid_reg;
  assign line_1297_clock = clock;
  assign line_1297_reset = reset;
  assign line_1297_valid = do_deq ^ line_1297_valid_reg;
  assign line_1298_clock = clock;
  assign line_1298_reset = reset;
  assign line_1298_valid = _T ^ line_1298_valid_reg;
  assign io_enq_ready = ~full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_resp = ram_resp_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_echo_real_last = ram_echo_real_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_resp_MPORT_en & ram_resp_MPORT_mask) begin
      ram_resp[ram_resp_MPORT_addr] <= ram_resp_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_echo_real_last_MPORT_en & ram_echo_real_last_MPORT_mask) begin
      ram_echo_real_last[ram_echo_real_last_MPORT_addr] <= ram_echo_real_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_enq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 292:16]
      enq_ptr_value <= enq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 1'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 296:16]
      deq_ptr_value <= deq_ptr_value + 1'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      maybe_full <= do_enq; // @[src/main/scala/chisel3/util/Decoupled.scala 300:16]
    end
    line_1296_valid_reg <= do_enq;
    line_1297_valid_reg <= do_deq;
    line_1298_valid_reg <= _T;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_echo_real_last[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_4[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1296_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1297_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1298_valid_reg = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_echo_real_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
  wire  nodeOut_aw_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeOut_aw_deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_aw_deq_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_enq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeOut_aw_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_aw_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_aw_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_w_deq_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_w_deq_q_io_enq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeOut_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] nodeOut_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeIn_b_deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_b_deq_q_io_enq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_enq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeIn_b_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_b_deq_q_io_deq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_b_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeOut_ar_deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_ar_deq_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_enq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeOut_ar_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] nodeOut_ar_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeOut_ar_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeIn_r_deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_r_deq_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_r_deq_q_io_enq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_enq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] nodeIn_r_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] nodeIn_r_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] nodeIn_r_deq_q_io_deq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  nodeIn_r_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  Queue_47 nodeOut_aw_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_aw_deq_q_clock),
    .reset(nodeOut_aw_deq_q_reset),
    .io_enq_ready(nodeOut_aw_deq_q_io_enq_ready),
    .io_enq_valid(nodeOut_aw_deq_q_io_enq_valid),
    .io_enq_bits_id(nodeOut_aw_deq_q_io_enq_bits_id),
    .io_enq_bits_addr(nodeOut_aw_deq_q_io_enq_bits_addr),
    .io_enq_bits_echo_real_last(nodeOut_aw_deq_q_io_enq_bits_echo_real_last),
    .io_deq_ready(nodeOut_aw_deq_q_io_deq_ready),
    .io_deq_valid(nodeOut_aw_deq_q_io_deq_valid),
    .io_deq_bits_id(nodeOut_aw_deq_q_io_deq_bits_id),
    .io_deq_bits_addr(nodeOut_aw_deq_q_io_deq_bits_addr),
    .io_deq_bits_echo_real_last(nodeOut_aw_deq_q_io_deq_bits_echo_real_last)
  );
  Queue_48 nodeOut_w_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_w_deq_q_clock),
    .reset(nodeOut_w_deq_q_reset),
    .io_enq_ready(nodeOut_w_deq_q_io_enq_ready),
    .io_enq_valid(nodeOut_w_deq_q_io_enq_valid),
    .io_enq_bits_data(nodeOut_w_deq_q_io_enq_bits_data),
    .io_enq_bits_strb(nodeOut_w_deq_q_io_enq_bits_strb),
    .io_deq_ready(nodeOut_w_deq_q_io_deq_ready),
    .io_deq_valid(nodeOut_w_deq_q_io_deq_valid),
    .io_deq_bits_data(nodeOut_w_deq_q_io_deq_bits_data),
    .io_deq_bits_strb(nodeOut_w_deq_q_io_deq_bits_strb)
  );
  Queue_49 nodeIn_b_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeIn_b_deq_q_clock),
    .reset(nodeIn_b_deq_q_reset),
    .io_enq_ready(nodeIn_b_deq_q_io_enq_ready),
    .io_enq_valid(nodeIn_b_deq_q_io_enq_valid),
    .io_enq_bits_id(nodeIn_b_deq_q_io_enq_bits_id),
    .io_enq_bits_resp(nodeIn_b_deq_q_io_enq_bits_resp),
    .io_enq_bits_echo_real_last(nodeIn_b_deq_q_io_enq_bits_echo_real_last),
    .io_deq_ready(nodeIn_b_deq_q_io_deq_ready),
    .io_deq_valid(nodeIn_b_deq_q_io_deq_valid),
    .io_deq_bits_id(nodeIn_b_deq_q_io_deq_bits_id),
    .io_deq_bits_resp(nodeIn_b_deq_q_io_deq_bits_resp),
    .io_deq_bits_echo_real_last(nodeIn_b_deq_q_io_deq_bits_echo_real_last)
  );
  Queue_50 nodeOut_ar_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeOut_ar_deq_q_clock),
    .reset(nodeOut_ar_deq_q_reset),
    .io_enq_ready(nodeOut_ar_deq_q_io_enq_ready),
    .io_enq_valid(nodeOut_ar_deq_q_io_enq_valid),
    .io_enq_bits_id(nodeOut_ar_deq_q_io_enq_bits_id),
    .io_enq_bits_addr(nodeOut_ar_deq_q_io_enq_bits_addr),
    .io_enq_bits_echo_real_last(nodeOut_ar_deq_q_io_enq_bits_echo_real_last),
    .io_deq_ready(nodeOut_ar_deq_q_io_deq_ready),
    .io_deq_valid(nodeOut_ar_deq_q_io_deq_valid),
    .io_deq_bits_id(nodeOut_ar_deq_q_io_deq_bits_id),
    .io_deq_bits_addr(nodeOut_ar_deq_q_io_deq_bits_addr),
    .io_deq_bits_echo_real_last(nodeOut_ar_deq_q_io_deq_bits_echo_real_last)
  );
  Queue_51 nodeIn_r_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(nodeIn_r_deq_q_clock),
    .reset(nodeIn_r_deq_q_reset),
    .io_enq_ready(nodeIn_r_deq_q_io_enq_ready),
    .io_enq_valid(nodeIn_r_deq_q_io_enq_valid),
    .io_enq_bits_id(nodeIn_r_deq_q_io_enq_bits_id),
    .io_enq_bits_data(nodeIn_r_deq_q_io_enq_bits_data),
    .io_enq_bits_resp(nodeIn_r_deq_q_io_enq_bits_resp),
    .io_enq_bits_echo_real_last(nodeIn_r_deq_q_io_enq_bits_echo_real_last),
    .io_deq_ready(nodeIn_r_deq_q_io_deq_ready),
    .io_deq_valid(nodeIn_r_deq_q_io_deq_valid),
    .io_deq_bits_id(nodeIn_r_deq_q_io_deq_bits_id),
    .io_deq_bits_data(nodeIn_r_deq_q_io_deq_bits_data),
    .io_deq_bits_resp(nodeIn_r_deq_q_io_deq_bits_resp),
    .io_deq_bits_echo_real_last(nodeIn_r_deq_q_io_deq_bits_echo_real_last),
    .io_deq_bits_last(nodeIn_r_deq_q_io_deq_bits_last)
  );
  assign auto_in_aw_ready = nodeOut_aw_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_w_ready = nodeOut_w_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_b_valid = nodeIn_b_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_in_b_bits_id = nodeIn_b_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_b_bits_resp = nodeIn_b_deq_q_io_deq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_b_bits_echo_real_last = nodeIn_b_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_ar_ready = nodeOut_ar_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_r_valid = nodeIn_r_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_in_r_bits_id = nodeIn_r_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_r_bits_data = nodeIn_r_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_r_bits_resp = nodeIn_r_deq_q_io_deq_bits_resp; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_r_bits_echo_real_last = nodeIn_r_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_in_r_bits_last = nodeIn_r_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_valid = nodeOut_aw_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_out_aw_bits_id = nodeOut_aw_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_addr = nodeOut_aw_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_echo_real_last = nodeOut_aw_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_valid = nodeOut_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_out_w_bits_data = nodeOut_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_bits_strb = nodeOut_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_b_ready = nodeIn_b_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_out_ar_valid = nodeOut_ar_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_out_ar_bits_id = nodeOut_ar_deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_addr = nodeOut_ar_deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_echo_real_last = nodeOut_ar_deq_q_io_deq_bits_echo_real_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_r_ready = nodeIn_r_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign nodeOut_aw_deq_q_clock = clock;
  assign nodeOut_aw_deq_q_reset = reset;
  assign nodeOut_aw_deq_q_io_enq_valid = auto_in_aw_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_aw_deq_q_io_enq_bits_id = auto_in_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_aw_deq_q_io_enq_bits_addr = auto_in_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_aw_deq_q_io_enq_bits_echo_real_last = auto_in_aw_bits_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_aw_deq_q_io_deq_ready = auto_out_aw_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeOut_w_deq_q_clock = clock;
  assign nodeOut_w_deq_q_reset = reset;
  assign nodeOut_w_deq_q_io_enq_valid = auto_in_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_w_deq_q_io_enq_bits_data = auto_in_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_w_deq_q_io_enq_bits_strb = auto_in_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_w_deq_q_io_deq_ready = auto_out_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_deq_q_clock = clock;
  assign nodeIn_b_deq_q_reset = reset;
  assign nodeIn_b_deq_q_io_enq_valid = auto_out_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_deq_q_io_enq_bits_id = auto_out_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_deq_q_io_enq_bits_resp = auto_out_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_deq_q_io_enq_bits_echo_real_last = auto_out_b_bits_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_b_deq_q_io_deq_ready = auto_in_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_ar_deq_q_clock = clock;
  assign nodeOut_ar_deq_q_reset = reset;
  assign nodeOut_ar_deq_q_io_enq_valid = auto_in_ar_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_ar_deq_q_io_enq_bits_id = auto_in_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_ar_deq_q_io_enq_bits_addr = auto_in_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_ar_deq_q_io_enq_bits_echo_real_last = auto_in_ar_bits_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign nodeOut_ar_deq_q_io_deq_ready = auto_out_ar_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_clock = clock;
  assign nodeIn_r_deq_q_reset = reset;
  assign nodeIn_r_deq_q_io_enq_valid = auto_out_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_io_enq_bits_id = auto_out_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_io_enq_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_io_enq_bits_resp = auto_out_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_io_enq_bits_echo_real_last = auto_out_r_bits_echo_real_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign nodeIn_r_deq_q_io_deq_ready = auto_in_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
endmodule
module Queue_52(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_burst, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_burst // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_addr [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_len [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_burst [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_23 = io_deq_ready ? 1'h0 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 324:26 286:27 324:35]
  wire  do_enq = empty ? _GEN_23 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 286:27]
  wire  line_1299_clock;
  wire  line_1299_reset;
  wire  line_1299_valid;
  reg  line_1299_valid_reg;
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 323:14 287:27]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1300_clock;
  wire  line_1300_reset;
  wire  line_1300_valid;
  reg  line_1300_valid_reg;
  wire  line_1301_clock;
  wire  line_1301_reset;
  wire  line_1301_valid;
  reg  line_1301_valid_reg;
  wire  line_1302_clock;
  wire  line_1302_reset;
  wire  line_1302_valid;
  reg  line_1302_valid_reg;
  wire  line_1303_clock;
  wire  line_1303_reset;
  wire  line_1303_valid;
  reg  line_1303_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1299)) line_1299 (
    .clock(line_1299_clock),
    .reset(line_1299_reset),
    .valid(line_1299_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1300)) line_1300 (
    .clock(line_1300_clock),
    .reset(line_1300_reset),
    .valid(line_1300_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1301)) line_1301 (
    .clock(line_1301_clock),
    .reset(line_1301_reset),
    .valid(line_1301_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1302)) line_1302 (
    .clock(line_1302_clock),
    .reset(line_1302_reset),
    .valid(line_1302_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1303)) line_1303 (
    .clock(line_1303_clock),
    .reset(line_1303_reset),
    .valid(line_1303_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign line_1299_clock = clock;
  assign line_1299_reset = reset;
  assign line_1299_valid = do_enq ^ line_1299_valid_reg;
  assign line_1300_clock = clock;
  assign line_1300_reset = reset;
  assign line_1300_valid = _T ^ line_1300_valid_reg;
  assign line_1301_clock = clock;
  assign line_1301_reset = reset;
  assign line_1301_valid = io_enq_valid ^ line_1301_valid_reg;
  assign line_1302_clock = clock;
  assign line_1302_reset = reset;
  assign line_1302_valid = empty ^ line_1302_valid_reg;
  assign line_1303_clock = clock;
  assign line_1303_reset = reset;
  assign line_1303_valid = io_deq_ready ^ line_1303_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:16 320:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
        if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
          maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
        end else begin
          maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end
    if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
      if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
        line_1299_valid_reg <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
      end else begin
        line_1299_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end else begin
      line_1299_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
    end
    line_1300_valid_reg <= _T;
    line_1301_valid_reg <= io_enq_valid;
    line_1302_valid_reg <= empty;
    line_1303_valid_reg <= io_deq_ready;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1299_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1300_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1301_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1302_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1303_valid_reg = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_53(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [3:0]  io_enq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [31:0] io_enq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [2:0]  io_enq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [1:0]  io_enq_bits_burst, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [3:0]  io_deq_bits_id, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [31:0] io_deq_bits_addr, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_len, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [2:0]  io_deq_bits_size, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [1:0]  io_deq_bits_burst // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] ram_id [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [3:0] ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_id_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [31:0] ram_addr [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [31:0] ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_addr_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_len [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_len_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [2:0] ram_size [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [2:0] ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_size_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [1:0] ram_burst [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [1:0] ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_burst_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_23 = io_deq_ready ? 1'h0 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 324:26 286:27 324:35]
  wire  do_enq = empty ? _GEN_23 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 286:27]
  wire  line_1304_clock;
  wire  line_1304_reset;
  wire  line_1304_valid;
  reg  line_1304_valid_reg;
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 323:14 287:27]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1305_clock;
  wire  line_1305_reset;
  wire  line_1305_valid;
  reg  line_1305_valid_reg;
  wire  line_1306_clock;
  wire  line_1306_reset;
  wire  line_1306_valid;
  reg  line_1306_valid_reg;
  wire  line_1307_clock;
  wire  line_1307_reset;
  wire  line_1307_valid;
  reg  line_1307_valid_reg;
  wire  line_1308_clock;
  wire  line_1308_reset;
  wire  line_1308_valid;
  reg  line_1308_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1304)) line_1304 (
    .clock(line_1304_clock),
    .reset(line_1304_reset),
    .valid(line_1304_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1305)) line_1305 (
    .clock(line_1305_clock),
    .reset(line_1305_reset),
    .valid(line_1305_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1306)) line_1306 (
    .clock(line_1306_clock),
    .reset(line_1306_reset),
    .valid(line_1306_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1307)) line_1307 (
    .clock(line_1307_clock),
    .reset(line_1307_reset),
    .valid(line_1307_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1308)) line_1308 (
    .clock(line_1308_clock),
    .reset(line_1308_reset),
    .valid(line_1308_valid)
  );
  assign ram_id_io_deq_bits_MPORT_en = 1'h1;
  assign ram_id_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = 1'h0;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_size_io_deq_bits_MPORT_en = 1'h1;
  assign ram_size_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = 1'h0;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign ram_burst_io_deq_bits_MPORT_en = 1'h1;
  assign ram_burst_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_burst_io_deq_bits_MPORT_data = ram_burst[ram_burst_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_burst_MPORT_data = io_enq_bits_burst;
  assign ram_burst_MPORT_addr = 1'h0;
  assign ram_burst_MPORT_mask = 1'h1;
  assign ram_burst_MPORT_en = empty ? _GEN_23 : _do_enq_T;
  assign line_1304_clock = clock;
  assign line_1304_reset = reset;
  assign line_1304_valid = do_enq ^ line_1304_valid_reg;
  assign line_1305_clock = clock;
  assign line_1305_reset = reset;
  assign line_1305_valid = _T ^ line_1305_valid_reg;
  assign line_1306_clock = clock;
  assign line_1306_reset = reset;
  assign line_1306_valid = io_enq_valid ^ line_1306_valid_reg;
  assign line_1307_clock = clock;
  assign line_1307_reset = reset;
  assign line_1307_valid = empty ^ line_1307_valid_reg;
  assign line_1308_clock = clock;
  assign line_1308_reset = reset;
  assign line_1308_valid = io_deq_ready ^ line_1308_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:16 320:{24,39}]
  assign io_deq_bits_id = empty ? io_enq_bits_id : ram_id_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_addr = empty ? io_enq_bits_addr : ram_addr_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_len = empty ? io_enq_bits_len : ram_len_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_size = empty ? io_enq_bits_size : ram_size_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_burst = empty ? io_enq_bits_burst : ram_burst_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  always @(posedge clock) begin
    if (ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_burst_MPORT_en & ram_burst_MPORT_mask) begin
      ram_burst[ram_burst_MPORT_addr] <= ram_burst_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
        if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
          maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
        end else begin
          maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end
    if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
      if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
        line_1304_valid_reg <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
      end else begin
        line_1304_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end else begin
      line_1304_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
    end
    line_1305_valid_reg <= _T;
    line_1306_valid_reg <= io_enq_valid;
    line_1307_valid_reg <= empty;
    line_1308_valid_reg <= io_deq_ready;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1304_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1305_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1306_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_1307_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1308_valid_reg = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_54(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [63:0] io_enq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input  [7:0]  io_enq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_enq_bits_last, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  input         io_deq_ready, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_valid, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [63:0] io_deq_bits_data, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output [7:0]  io_deq_bits_strb, // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
  output        io_deq_bits_last // @[src/main/scala/chisel3/util/Decoupled.scala 278:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_data [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [63:0] ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_data_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg [7:0] ram_strb [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire [7:0] ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_strb_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  ram_last [0:0]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_mask; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  wire  ram_last_MPORT_en; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  reg  maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
  wire  empty = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 284:28]
  wire  _do_enq_T = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _do_deq_T = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_17 = io_deq_ready ? 1'h0 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 324:26 286:27 324:35]
  wire  do_enq = empty ? _GEN_17 : _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 286:27]
  wire  line_1309_clock;
  wire  line_1309_reset;
  wire  line_1309_valid;
  reg  line_1309_valid_reg;
  wire  do_deq = empty ? 1'h0 : _do_deq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 321:17 323:14 287:27]
  wire  _T = do_enq != do_deq; // @[src/main/scala/chisel3/util/Decoupled.scala 299:15]
  wire  line_1310_clock;
  wire  line_1310_reset;
  wire  line_1310_valid;
  reg  line_1310_valid_reg;
  wire  line_1311_clock;
  wire  line_1311_reset;
  wire  line_1311_valid;
  reg  line_1311_valid_reg;
  wire  line_1312_clock;
  wire  line_1312_reset;
  wire  line_1312_valid;
  reg  line_1312_valid_reg;
  wire  line_1313_clock;
  wire  line_1313_reset;
  wire  line_1313_valid;
  reg  line_1313_valid_reg;
  GEN_w1_line #(.COVER_INDEX(1309)) line_1309 (
    .clock(line_1309_clock),
    .reset(line_1309_reset),
    .valid(line_1309_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1310)) line_1310 (
    .clock(line_1310_clock),
    .reset(line_1310_reset),
    .valid(line_1310_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1311)) line_1311 (
    .clock(line_1311_clock),
    .reset(line_1311_reset),
    .valid(line_1311_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1312)) line_1312 (
    .clock(line_1312_clock),
    .reset(line_1312_reset),
    .valid(line_1312_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1313)) line_1313 (
    .clock(line_1313_clock),
    .reset(line_1313_reset),
    .valid(line_1313_valid)
  );
  assign ram_data_io_deq_bits_MPORT_en = 1'h1;
  assign ram_data_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = 1'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_strb_io_deq_bits_MPORT_en = 1'h1;
  assign ram_strb_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_strb_io_deq_bits_MPORT_data = ram_strb[ram_strb_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_strb_MPORT_data = io_enq_bits_strb;
  assign ram_strb_MPORT_addr = 1'h0;
  assign ram_strb_MPORT_mask = 1'h1;
  assign ram_strb_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign ram_last_io_deq_bits_MPORT_en = 1'h1;
  assign ram_last_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = 1'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = empty ? _GEN_17 : _do_enq_T;
  assign line_1309_clock = clock;
  assign line_1309_reset = reset;
  assign line_1309_valid = do_enq ^ line_1309_valid_reg;
  assign line_1310_clock = clock;
  assign line_1310_reset = reset;
  assign line_1310_valid = _T ^ line_1310_valid_reg;
  assign line_1311_clock = clock;
  assign line_1311_reset = reset;
  assign line_1311_valid = io_enq_valid ^ line_1311_valid_reg;
  assign line_1312_clock = clock;
  assign line_1312_reset = reset;
  assign line_1312_valid = empty ^ line_1312_valid_reg;
  assign line_1313_clock = clock;
  assign line_1313_reset = reset;
  assign line_1313_valid = io_deq_ready ^ line_1313_valid_reg;
  assign io_enq_ready = ~maybe_full; // @[src/main/scala/chisel3/util/Decoupled.scala 309:19]
  assign io_deq_valid = io_enq_valid | ~empty; // @[src/main/scala/chisel3/util/Decoupled.scala 308:16 320:{24,39}]
  assign io_deq_bits_data = empty ? io_enq_bits_data : ram_data_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_strb = empty ? io_enq_bits_strb : ram_strb_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  assign io_deq_bits_last = empty ? io_enq_bits_last : ram_last_io_deq_bits_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 316:17 321:17 322:19]
  always @(posedge clock) begin
    if (ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_strb_MPORT_en & ram_strb_MPORT_mask) begin
      ram_strb[ram_strb_MPORT_addr] <= ram_strb_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[src/main/scala/chisel3/util/Decoupled.scala 279:95]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
      maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 282:27]
    end else if (do_enq != do_deq) begin // @[src/main/scala/chisel3/util/Decoupled.scala 299:27]
      if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
        if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
          maybe_full <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
        end else begin
          maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
        end
      end else begin
        maybe_full <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end
    if (empty) begin // @[src/main/scala/chisel3/util/Decoupled.scala 321:17]
      if (io_deq_ready) begin // @[src/main/scala/chisel3/util/Decoupled.scala 324:26]
        line_1309_valid_reg <= 1'h0; // @[src/main/scala/chisel3/util/Decoupled.scala 324:35]
      end else begin
        line_1309_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
      end
    end else begin
      line_1309_valid_reg <= _do_enq_T; // @[src/main/scala/chisel3/util/Decoupled.scala 286:27]
    end
    line_1310_valid_reg <= _T;
    line_1311_valid_reg <= io_enq_valid;
    line_1312_valid_reg <= empty;
    line_1313_valid_reg <= io_deq_ready;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1309_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1310_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  line_1311_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  line_1312_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_1313_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  output        auto_in_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_aw_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_aw_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_aw_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_in_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_w_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_in_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [31:0] auto_in_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [7:0]  auto_in_ar_bits_len, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [2:0]  auto_in_ar_bits_size, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_in_ar_bits_burst, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_in_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_in_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_in_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [1:0]  auto_in_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_in_r_bits_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_aw_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_aw_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_aw_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_aw_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_w_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_w_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [63:0] auto_out_w_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [7:0]  auto_out_w_bits_strb, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_b_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_b_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_b_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_b_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_ar_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [3:0]  auto_out_ar_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output [31:0] auto_out_ar_bits_addr, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_ar_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  output        auto_out_r_ready, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_valid, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [3:0]  auto_out_r_bits_id, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [63:0] auto_out_r_bits_data, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input  [1:0]  auto_out_r_bits_resp, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_echo_real_last, // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
  input         auto_out_r_bits_last // @[src/main/scala/diplomacy/LazyModule.scala 366:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire  deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] deq_q_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] deq_q_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] deq_q_io_enq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] deq_q_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] deq_q_io_enq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] deq_q_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] deq_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] deq_q_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] deq_q_1_io_enq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] deq_q_1_io_enq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] deq_q_1_io_enq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] deq_q_1_io_enq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] deq_q_1_io_enq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  deq_q_1_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [3:0] deq_q_1_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [31:0] deq_q_1_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] deq_q_1_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [2:0] deq_q_1_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [1:0] deq_q_1_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_clock; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_reset; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_enq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] in_w_deq_q_io_enq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] in_w_deq_q_io_enq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_enq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_deq_ready; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [63:0] in_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire [7:0] in_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  wire  in_w_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
  reg  busy; // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
  reg [31:0] r_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 65:25]
  reg [7:0] r_len; // @[src/main/scala/amba/axi4/Fragmenter.scala 66:25]
  wire [7:0] irr_bits_len = deq_q_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [7:0] len = busy ? r_len : irr_bits_len; // @[src/main/scala/amba/axi4/Fragmenter.scala 68:23]
  wire [31:0] irr_bits_addr = deq_q_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [31:0] addr = busy ? r_addr : irr_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 69:23]
  wire [1:0] irr_bits_burst = deq_q_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire  fixed = irr_bits_burst == 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 96:34]
  wire [2:0] irr_bits_size = deq_q_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [15:0] _inc_addr_T = 16'h1 << irr_bits_size; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:38]
  wire [31:0] _GEN_92 = {{16'd0}, _inc_addr_T}; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:29]
  wire [31:0] inc_addr = addr + _GEN_92; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:29]
  wire [15:0] _wrapMask_T = {irr_bits_len,8'hff}; // @[src/main/scala/amba/axi4/Bundles.scala 33:9]
  wire [22:0] _GEN_45 = {{7'd0}, _wrapMask_T}; // @[src/main/scala/amba/axi4/Bundles.scala 33:21]
  wire [22:0] _wrapMask_T_1 = _GEN_45 << irr_bits_size; // @[src/main/scala/amba/axi4/Bundles.scala 33:21]
  wire [14:0] wrapMask = _wrapMask_T_1[22:8]; // @[src/main/scala/amba/axi4/Bundles.scala 33:30]
  wire  _T = irr_bits_burst == 2'h2; // @[src/main/scala/amba/axi4/Fragmenter.scala 107:28]
  wire  line_1314_clock;
  wire  line_1314_reset;
  wire  line_1314_valid;
  reg  line_1314_valid_reg;
  wire [31:0] _GEN_93 = {{17'd0}, wrapMask}; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:33]
  wire [31:0] _mux_addr_T = inc_addr & _GEN_93; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:33]
  wire [31:0] _mux_addr_T_1 = ~irr_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:49]
  wire [31:0] _mux_addr_T_2 = _mux_addr_T_1 | _GEN_93; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:62]
  wire [31:0] _mux_addr_T_3 = ~_mux_addr_T_2; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:47]
  wire [31:0] _mux_addr_T_4 = _mux_addr_T | _mux_addr_T_3; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:45]
  wire  line_1315_clock;
  wire  line_1315_reset;
  wire  line_1315_valid;
  reg  line_1315_valid_reg;
  wire  ar_last = 8'h0 == len; // @[src/main/scala/amba/axi4/Fragmenter.scala 114:27]
  wire [31:0] _out_bits_addr_T = ~addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:28]
  wire [9:0] _out_bits_addr_T_2 = 10'h7 << irr_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [2:0] _out_bits_addr_T_4 = ~_out_bits_addr_T_2[2:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [31:0] _GEN_95 = {{29'd0}, _out_bits_addr_T_4}; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:34]
  wire [31:0] _out_bits_addr_T_5 = _out_bits_addr_T | _GEN_95; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:34]
  wire  irr_valid = deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  wire  _T_2 = auto_out_ar_ready & irr_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1316_clock;
  wire  line_1316_reset;
  wire  line_1316_valid;
  reg  line_1316_valid_reg;
  wire [8:0] _GEN_96 = {{1'd0}, len}; // @[src/main/scala/amba/axi4/Fragmenter.scala 131:25]
  wire [8:0] _r_len_T_1 = _GEN_96 - 9'h1; // @[src/main/scala/amba/axi4/Fragmenter.scala 131:25]
  wire [8:0] _GEN_48 = _T_2 ? _r_len_T_1 : {{1'd0}, r_len}; // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25 131:18 66:25]
  reg  busy_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
  reg [31:0] r_addr_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 65:25]
  reg [7:0] r_len_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 66:25]
  wire [7:0] irr_1_bits_len = deq_q_1_io_deq_bits_len; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [7:0] len_1 = busy_1 ? r_len_1 : irr_1_bits_len; // @[src/main/scala/amba/axi4/Fragmenter.scala 68:23]
  wire [31:0] irr_1_bits_addr = deq_q_1_io_deq_bits_addr; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [31:0] addr_1 = busy_1 ? r_addr_1 : irr_1_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 69:23]
  wire [1:0] irr_1_bits_burst = deq_q_1_io_deq_bits_burst; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire  fixed_1 = irr_1_bits_burst == 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 96:34]
  wire [2:0] irr_1_bits_size = deq_q_1_io_deq_bits_size; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire [15:0] _inc_addr_T_2 = 16'h1 << irr_1_bits_size; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:38]
  wire [31:0] _GEN_101 = {{16'd0}, _inc_addr_T_2}; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:29]
  wire [31:0] inc_addr_1 = addr_1 + _GEN_101; // @[src/main/scala/amba/axi4/Fragmenter.scala 104:29]
  wire [15:0] _wrapMask_T_2 = {irr_1_bits_len,8'hff}; // @[src/main/scala/amba/axi4/Bundles.scala 33:9]
  wire [22:0] _GEN_47 = {{7'd0}, _wrapMask_T_2}; // @[src/main/scala/amba/axi4/Bundles.scala 33:21]
  wire [22:0] _wrapMask_T_3 = _GEN_47 << irr_1_bits_size; // @[src/main/scala/amba/axi4/Bundles.scala 33:21]
  wire [14:0] wrapMask_1 = _wrapMask_T_3[22:8]; // @[src/main/scala/amba/axi4/Bundles.scala 33:30]
  wire  _T_3 = irr_1_bits_burst == 2'h2; // @[src/main/scala/amba/axi4/Fragmenter.scala 107:28]
  wire  line_1317_clock;
  wire  line_1317_reset;
  wire  line_1317_valid;
  reg  line_1317_valid_reg;
  wire [31:0] _GEN_102 = {{17'd0}, wrapMask_1}; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:33]
  wire [31:0] _mux_addr_T_5 = inc_addr_1 & _GEN_102; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:33]
  wire [31:0] _mux_addr_T_6 = ~irr_1_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:49]
  wire [31:0] _mux_addr_T_7 = _mux_addr_T_6 | _GEN_102; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:62]
  wire [31:0] _mux_addr_T_8 = ~_mux_addr_T_7; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:47]
  wire [31:0] _mux_addr_T_9 = _mux_addr_T_5 | _mux_addr_T_8; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:45]
  wire  line_1318_clock;
  wire  line_1318_reset;
  wire  line_1318_valid;
  reg  line_1318_valid_reg;
  wire  aw_last = 8'h0 == len_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 114:27]
  reg [8:0] w_counter; // @[src/main/scala/amba/axi4/Fragmenter.scala 172:30]
  wire  w_idle = w_counter == 9'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 173:30]
  reg  wbeats_latched; // @[src/main/scala/amba/axi4/Fragmenter.scala 156:35]
  wire  _in_aw_ready_T = w_idle | wbeats_latched; // @[src/main/scala/amba/axi4/Fragmenter.scala 164:52]
  wire  in_aw_ready = auto_out_aw_ready & (w_idle | wbeats_latched); // @[src/main/scala/amba/axi4/Fragmenter.scala 164:35]
  wire [31:0] _out_bits_addr_T_7 = ~addr_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:28]
  wire [9:0] _out_bits_addr_T_9 = 10'h7 << irr_1_bits_size; // @[src/main/scala/util/package.scala 235:71]
  wire [2:0] _out_bits_addr_T_11 = ~_out_bits_addr_T_9[2:0]; // @[src/main/scala/util/package.scala 235:46]
  wire [31:0] _GEN_104 = {{29'd0}, _out_bits_addr_T_11}; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:34]
  wire [31:0] _out_bits_addr_T_12 = _out_bits_addr_T_7 | _GEN_104; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:34]
  wire  irr_1_valid = deq_q_1_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  wire  _T_5 = in_aw_ready & irr_1_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1319_clock;
  wire  line_1319_reset;
  wire  line_1319_valid;
  reg  line_1319_valid_reg;
  wire [8:0] _GEN_105 = {{1'd0}, len_1}; // @[src/main/scala/amba/axi4/Fragmenter.scala 131:25]
  wire [8:0] _r_len_T_3 = _GEN_105 - 9'h1; // @[src/main/scala/amba/axi4/Fragmenter.scala 131:25]
  wire [8:0] _GEN_53 = _T_5 ? _r_len_T_3 : {{1'd0}, r_len_1}; // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25 131:18 66:25]
  wire  wbeats_valid = irr_1_valid & ~wbeats_latched; // @[src/main/scala/amba/axi4/Fragmenter.scala 165:35]
  wire  _T_6 = wbeats_valid & w_idle; // @[src/main/scala/amba/axi4/Fragmenter.scala 159:26]
  wire  line_1320_clock;
  wire  line_1320_reset;
  wire  line_1320_valid;
  reg  line_1320_valid_reg;
  wire  _GEN_54 = wbeats_valid & w_idle | wbeats_latched; // @[src/main/scala/amba/axi4/Fragmenter.scala 156:35 159:{43,60}]
  wire  nodeOut_aw_valid = irr_1_valid & _in_aw_ready_T; // @[src/main/scala/amba/axi4/Fragmenter.scala 163:35]
  wire  _T_7 = auto_out_aw_ready & nodeOut_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  line_1321_clock;
  wire  line_1321_reset;
  wire  line_1321_valid;
  reg  line_1321_valid_reg;
  wire [8:0] _w_todo_T = wbeats_valid ? 9'h1 : 9'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 174:35]
  wire [8:0] w_todo = w_idle ? _w_todo_T : w_counter; // @[src/main/scala/amba/axi4/Fragmenter.scala 174:23]
  wire  w_last = w_todo == 9'h1; // @[src/main/scala/amba/axi4/Fragmenter.scala 175:27]
  wire  in_w_valid = in_w_deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  wire  _nodeOut_w_valid_T_1 = ~w_idle | wbeats_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 181:51]
  wire  nodeOut_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[src/main/scala/amba/axi4/Fragmenter.scala 181:33]
  wire  _w_counter_T = auto_out_w_ready & nodeOut_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [8:0] _GEN_106 = {{8'd0}, _w_counter_T}; // @[src/main/scala/amba/axi4/Fragmenter.scala 176:27]
  wire [8:0] _w_counter_T_2 = w_todo - _GEN_106; // @[src/main/scala/amba/axi4/Fragmenter.scala 176:27]
  wire  _T_13 = ~reset; // @[src/main/scala/amba/axi4/Fragmenter.scala 177:14]
  wire  line_1322_clock;
  wire  line_1322_reset;
  wire  line_1322_valid;
  reg  line_1322_valid_reg;
  wire  _T_14 = ~(~_w_counter_T | w_todo != 9'h0); // @[src/main/scala/amba/axi4/Fragmenter.scala 177:14]
  wire  line_1323_clock;
  wire  line_1323_reset;
  wire  line_1323_valid;
  reg  line_1323_valid_reg;
  wire  in_w_bits_last = in_w_deq_q_io_deq_bits_last; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  wire  line_1324_clock;
  wire  line_1324_reset;
  wire  line_1324_valid;
  reg  line_1324_valid_reg;
  wire  _T_21 = ~(~nodeOut_w_valid | ~in_w_bits_last | w_last); // @[src/main/scala/amba/axi4/Fragmenter.scala 186:14]
  wire  line_1325_clock;
  wire  line_1325_reset;
  wire  line_1325_valid;
  reg  line_1325_valid_reg;
  wire  nodeOut_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 204:33]
  reg [1:0] error_0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_2; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_3; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_4; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_5; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_6; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_7; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_8; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_9; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_10; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_11; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_12; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_13; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_14; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  reg [1:0] error_15; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
  wire  line_1326_clock;
  wire  line_1326_reset;
  wire  line_1326_valid;
  reg  line_1326_valid_reg;
  wire  line_1327_clock;
  wire  line_1327_reset;
  wire  line_1327_valid;
  reg  line_1327_valid_reg;
  wire [1:0] _GEN_57 = 4'h1 == auto_out_b_bits_id ? error_1 : error_0; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1328_clock;
  wire  line_1328_reset;
  wire  line_1328_valid;
  reg  line_1328_valid_reg;
  wire [1:0] _GEN_58 = 4'h2 == auto_out_b_bits_id ? error_2 : _GEN_57; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1329_clock;
  wire  line_1329_reset;
  wire  line_1329_valid;
  reg  line_1329_valid_reg;
  wire [1:0] _GEN_59 = 4'h3 == auto_out_b_bits_id ? error_3 : _GEN_58; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1330_clock;
  wire  line_1330_reset;
  wire  line_1330_valid;
  reg  line_1330_valid_reg;
  wire [1:0] _GEN_60 = 4'h4 == auto_out_b_bits_id ? error_4 : _GEN_59; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1331_clock;
  wire  line_1331_reset;
  wire  line_1331_valid;
  reg  line_1331_valid_reg;
  wire [1:0] _GEN_61 = 4'h5 == auto_out_b_bits_id ? error_5 : _GEN_60; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1332_clock;
  wire  line_1332_reset;
  wire  line_1332_valid;
  reg  line_1332_valid_reg;
  wire [1:0] _GEN_62 = 4'h6 == auto_out_b_bits_id ? error_6 : _GEN_61; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1333_clock;
  wire  line_1333_reset;
  wire  line_1333_valid;
  reg  line_1333_valid_reg;
  wire [1:0] _GEN_63 = 4'h7 == auto_out_b_bits_id ? error_7 : _GEN_62; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1334_clock;
  wire  line_1334_reset;
  wire  line_1334_valid;
  reg  line_1334_valid_reg;
  wire [1:0] _GEN_64 = 4'h8 == auto_out_b_bits_id ? error_8 : _GEN_63; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1335_clock;
  wire  line_1335_reset;
  wire  line_1335_valid;
  reg  line_1335_valid_reg;
  wire [1:0] _GEN_65 = 4'h9 == auto_out_b_bits_id ? error_9 : _GEN_64; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1336_clock;
  wire  line_1336_reset;
  wire  line_1336_valid;
  reg  line_1336_valid_reg;
  wire [1:0] _GEN_66 = 4'ha == auto_out_b_bits_id ? error_10 : _GEN_65; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1337_clock;
  wire  line_1337_reset;
  wire  line_1337_valid;
  reg  line_1337_valid_reg;
  wire [1:0] _GEN_67 = 4'hb == auto_out_b_bits_id ? error_11 : _GEN_66; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1338_clock;
  wire  line_1338_reset;
  wire  line_1338_valid;
  reg  line_1338_valid_reg;
  wire [1:0] _GEN_68 = 4'hc == auto_out_b_bits_id ? error_12 : _GEN_67; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1339_clock;
  wire  line_1339_reset;
  wire  line_1339_valid;
  reg  line_1339_valid_reg;
  wire [1:0] _GEN_69 = 4'hd == auto_out_b_bits_id ? error_13 : _GEN_68; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1340_clock;
  wire  line_1340_reset;
  wire  line_1340_valid;
  reg  line_1340_valid_reg;
  wire [1:0] _GEN_70 = 4'he == auto_out_b_bits_id ? error_14 : _GEN_69; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire  line_1341_clock;
  wire  line_1341_reset;
  wire  line_1341_valid;
  reg  line_1341_valid_reg;
  wire [1:0] _GEN_71 = 4'hf == auto_out_b_bits_id ? error_15 : _GEN_70; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:{41,41}]
  wire [15:0] _T_22 = 16'h1 << auto_out_b_bits_id; // @[src/main/scala/chisel3/util/OneHot.scala 65:12]
  wire  _T_40 = nodeOut_b_ready & auto_out_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_41 = _T_22[0] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1342_clock;
  wire  line_1342_reset;
  wire  line_1342_valid;
  reg  line_1342_valid_reg;
  wire [1:0] _error_0_T = error_0 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_43 = _T_22[1] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1343_clock;
  wire  line_1343_reset;
  wire  line_1343_valid;
  reg  line_1343_valid_reg;
  wire [1:0] _error_1_T = error_1 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_45 = _T_22[2] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1344_clock;
  wire  line_1344_reset;
  wire  line_1344_valid;
  reg  line_1344_valid_reg;
  wire [1:0] _error_2_T = error_2 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_47 = _T_22[3] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1345_clock;
  wire  line_1345_reset;
  wire  line_1345_valid;
  reg  line_1345_valid_reg;
  wire [1:0] _error_3_T = error_3 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_49 = _T_22[4] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1346_clock;
  wire  line_1346_reset;
  wire  line_1346_valid;
  reg  line_1346_valid_reg;
  wire [1:0] _error_4_T = error_4 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_51 = _T_22[5] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1347_clock;
  wire  line_1347_reset;
  wire  line_1347_valid;
  reg  line_1347_valid_reg;
  wire [1:0] _error_5_T = error_5 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_53 = _T_22[6] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1348_clock;
  wire  line_1348_reset;
  wire  line_1348_valid;
  reg  line_1348_valid_reg;
  wire [1:0] _error_6_T = error_6 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_55 = _T_22[7] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1349_clock;
  wire  line_1349_reset;
  wire  line_1349_valid;
  reg  line_1349_valid_reg;
  wire [1:0] _error_7_T = error_7 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_57 = _T_22[8] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1350_clock;
  wire  line_1350_reset;
  wire  line_1350_valid;
  reg  line_1350_valid_reg;
  wire [1:0] _error_8_T = error_8 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_59 = _T_22[9] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1351_clock;
  wire  line_1351_reset;
  wire  line_1351_valid;
  reg  line_1351_valid_reg;
  wire [1:0] _error_9_T = error_9 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_61 = _T_22[10] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1352_clock;
  wire  line_1352_reset;
  wire  line_1352_valid;
  reg  line_1352_valid_reg;
  wire [1:0] _error_10_T = error_10 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_63 = _T_22[11] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1353_clock;
  wire  line_1353_reset;
  wire  line_1353_valid;
  reg  line_1353_valid_reg;
  wire [1:0] _error_11_T = error_11 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_65 = _T_22[12] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1354_clock;
  wire  line_1354_reset;
  wire  line_1354_valid;
  reg  line_1354_valid_reg;
  wire [1:0] _error_12_T = error_12 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_67 = _T_22[13] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1355_clock;
  wire  line_1355_reset;
  wire  line_1355_valid;
  reg  line_1355_valid_reg;
  wire [1:0] _error_13_T = error_13 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_69 = _T_22[14] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1356_clock;
  wire  line_1356_reset;
  wire  line_1356_valid;
  reg  line_1356_valid_reg;
  wire [1:0] _error_14_T = error_14 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  wire  _T_71 = _T_22[15] & _T_40; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:19]
  wire  line_1357_clock;
  wire  line_1357_reset;
  wire  line_1357_valid;
  reg  line_1357_valid_reg;
  wire [1:0] _error_15_T = error_15 | auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 210:64]
  Queue_52 deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(deq_q_clock),
    .reset(deq_q_reset),
    .io_enq_ready(deq_q_io_enq_ready),
    .io_enq_valid(deq_q_io_enq_valid),
    .io_enq_bits_id(deq_q_io_enq_bits_id),
    .io_enq_bits_addr(deq_q_io_enq_bits_addr),
    .io_enq_bits_len(deq_q_io_enq_bits_len),
    .io_enq_bits_size(deq_q_io_enq_bits_size),
    .io_enq_bits_burst(deq_q_io_enq_bits_burst),
    .io_deq_ready(deq_q_io_deq_ready),
    .io_deq_valid(deq_q_io_deq_valid),
    .io_deq_bits_id(deq_q_io_deq_bits_id),
    .io_deq_bits_addr(deq_q_io_deq_bits_addr),
    .io_deq_bits_len(deq_q_io_deq_bits_len),
    .io_deq_bits_size(deq_q_io_deq_bits_size),
    .io_deq_bits_burst(deq_q_io_deq_bits_burst)
  );
  Queue_53 deq_q_1 ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(deq_q_1_clock),
    .reset(deq_q_1_reset),
    .io_enq_ready(deq_q_1_io_enq_ready),
    .io_enq_valid(deq_q_1_io_enq_valid),
    .io_enq_bits_id(deq_q_1_io_enq_bits_id),
    .io_enq_bits_addr(deq_q_1_io_enq_bits_addr),
    .io_enq_bits_len(deq_q_1_io_enq_bits_len),
    .io_enq_bits_size(deq_q_1_io_enq_bits_size),
    .io_enq_bits_burst(deq_q_1_io_enq_bits_burst),
    .io_deq_ready(deq_q_1_io_deq_ready),
    .io_deq_valid(deq_q_1_io_deq_valid),
    .io_deq_bits_id(deq_q_1_io_deq_bits_id),
    .io_deq_bits_addr(deq_q_1_io_deq_bits_addr),
    .io_deq_bits_len(deq_q_1_io_deq_bits_len),
    .io_deq_bits_size(deq_q_1_io_deq_bits_size),
    .io_deq_bits_burst(deq_q_1_io_deq_bits_burst)
  );
  Queue_54 in_w_deq_q ( // @[src/main/scala/chisel3/util/Decoupled.scala 381:21]
    .clock(in_w_deq_q_clock),
    .reset(in_w_deq_q_reset),
    .io_enq_ready(in_w_deq_q_io_enq_ready),
    .io_enq_valid(in_w_deq_q_io_enq_valid),
    .io_enq_bits_data(in_w_deq_q_io_enq_bits_data),
    .io_enq_bits_strb(in_w_deq_q_io_enq_bits_strb),
    .io_enq_bits_last(in_w_deq_q_io_enq_bits_last),
    .io_deq_ready(in_w_deq_q_io_deq_ready),
    .io_deq_valid(in_w_deq_q_io_deq_valid),
    .io_deq_bits_data(in_w_deq_q_io_deq_bits_data),
    .io_deq_bits_strb(in_w_deq_q_io_deq_bits_strb),
    .io_deq_bits_last(in_w_deq_q_io_deq_bits_last)
  );
  GEN_w1_line #(.COVER_INDEX(1314)) line_1314 (
    .clock(line_1314_clock),
    .reset(line_1314_reset),
    .valid(line_1314_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1315)) line_1315 (
    .clock(line_1315_clock),
    .reset(line_1315_reset),
    .valid(line_1315_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1316)) line_1316 (
    .clock(line_1316_clock),
    .reset(line_1316_reset),
    .valid(line_1316_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1317)) line_1317 (
    .clock(line_1317_clock),
    .reset(line_1317_reset),
    .valid(line_1317_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1318)) line_1318 (
    .clock(line_1318_clock),
    .reset(line_1318_reset),
    .valid(line_1318_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1319)) line_1319 (
    .clock(line_1319_clock),
    .reset(line_1319_reset),
    .valid(line_1319_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1320)) line_1320 (
    .clock(line_1320_clock),
    .reset(line_1320_reset),
    .valid(line_1320_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1321)) line_1321 (
    .clock(line_1321_clock),
    .reset(line_1321_reset),
    .valid(line_1321_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1322)) line_1322 (
    .clock(line_1322_clock),
    .reset(line_1322_reset),
    .valid(line_1322_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1323)) line_1323 (
    .clock(line_1323_clock),
    .reset(line_1323_reset),
    .valid(line_1323_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1324)) line_1324 (
    .clock(line_1324_clock),
    .reset(line_1324_reset),
    .valid(line_1324_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1325)) line_1325 (
    .clock(line_1325_clock),
    .reset(line_1325_reset),
    .valid(line_1325_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1326)) line_1326 (
    .clock(line_1326_clock),
    .reset(line_1326_reset),
    .valid(line_1326_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1327)) line_1327 (
    .clock(line_1327_clock),
    .reset(line_1327_reset),
    .valid(line_1327_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1328)) line_1328 (
    .clock(line_1328_clock),
    .reset(line_1328_reset),
    .valid(line_1328_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1329)) line_1329 (
    .clock(line_1329_clock),
    .reset(line_1329_reset),
    .valid(line_1329_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1330)) line_1330 (
    .clock(line_1330_clock),
    .reset(line_1330_reset),
    .valid(line_1330_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1331)) line_1331 (
    .clock(line_1331_clock),
    .reset(line_1331_reset),
    .valid(line_1331_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1332)) line_1332 (
    .clock(line_1332_clock),
    .reset(line_1332_reset),
    .valid(line_1332_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1333)) line_1333 (
    .clock(line_1333_clock),
    .reset(line_1333_reset),
    .valid(line_1333_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1334)) line_1334 (
    .clock(line_1334_clock),
    .reset(line_1334_reset),
    .valid(line_1334_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1335)) line_1335 (
    .clock(line_1335_clock),
    .reset(line_1335_reset),
    .valid(line_1335_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1336)) line_1336 (
    .clock(line_1336_clock),
    .reset(line_1336_reset),
    .valid(line_1336_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1337)) line_1337 (
    .clock(line_1337_clock),
    .reset(line_1337_reset),
    .valid(line_1337_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1338)) line_1338 (
    .clock(line_1338_clock),
    .reset(line_1338_reset),
    .valid(line_1338_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1339)) line_1339 (
    .clock(line_1339_clock),
    .reset(line_1339_reset),
    .valid(line_1339_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1340)) line_1340 (
    .clock(line_1340_clock),
    .reset(line_1340_reset),
    .valid(line_1340_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1341)) line_1341 (
    .clock(line_1341_clock),
    .reset(line_1341_reset),
    .valid(line_1341_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1342)) line_1342 (
    .clock(line_1342_clock),
    .reset(line_1342_reset),
    .valid(line_1342_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1343)) line_1343 (
    .clock(line_1343_clock),
    .reset(line_1343_reset),
    .valid(line_1343_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1344)) line_1344 (
    .clock(line_1344_clock),
    .reset(line_1344_reset),
    .valid(line_1344_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1345)) line_1345 (
    .clock(line_1345_clock),
    .reset(line_1345_reset),
    .valid(line_1345_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1346)) line_1346 (
    .clock(line_1346_clock),
    .reset(line_1346_reset),
    .valid(line_1346_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1347)) line_1347 (
    .clock(line_1347_clock),
    .reset(line_1347_reset),
    .valid(line_1347_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1348)) line_1348 (
    .clock(line_1348_clock),
    .reset(line_1348_reset),
    .valid(line_1348_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1349)) line_1349 (
    .clock(line_1349_clock),
    .reset(line_1349_reset),
    .valid(line_1349_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1350)) line_1350 (
    .clock(line_1350_clock),
    .reset(line_1350_reset),
    .valid(line_1350_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1351)) line_1351 (
    .clock(line_1351_clock),
    .reset(line_1351_reset),
    .valid(line_1351_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1352)) line_1352 (
    .clock(line_1352_clock),
    .reset(line_1352_reset),
    .valid(line_1352_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1353)) line_1353 (
    .clock(line_1353_clock),
    .reset(line_1353_reset),
    .valid(line_1353_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1354)) line_1354 (
    .clock(line_1354_clock),
    .reset(line_1354_reset),
    .valid(line_1354_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1355)) line_1355 (
    .clock(line_1355_clock),
    .reset(line_1355_reset),
    .valid(line_1355_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1356)) line_1356 (
    .clock(line_1356_clock),
    .reset(line_1356_reset),
    .valid(line_1356_valid)
  );
  GEN_w1_line #(.COVER_INDEX(1357)) line_1357 (
    .clock(line_1357_clock),
    .reset(line_1357_reset),
    .valid(line_1357_valid)
  );
  assign line_1314_clock = clock;
  assign line_1314_reset = reset;
  assign line_1314_valid = _T ^ line_1314_valid_reg;
  assign line_1315_clock = clock;
  assign line_1315_reset = reset;
  assign line_1315_valid = fixed ^ line_1315_valid_reg;
  assign line_1316_clock = clock;
  assign line_1316_reset = reset;
  assign line_1316_valid = _T_2 ^ line_1316_valid_reg;
  assign line_1317_clock = clock;
  assign line_1317_reset = reset;
  assign line_1317_valid = _T_3 ^ line_1317_valid_reg;
  assign line_1318_clock = clock;
  assign line_1318_reset = reset;
  assign line_1318_valid = fixed_1 ^ line_1318_valid_reg;
  assign line_1319_clock = clock;
  assign line_1319_reset = reset;
  assign line_1319_valid = _T_5 ^ line_1319_valid_reg;
  assign line_1320_clock = clock;
  assign line_1320_reset = reset;
  assign line_1320_valid = _T_6 ^ line_1320_valid_reg;
  assign line_1321_clock = clock;
  assign line_1321_reset = reset;
  assign line_1321_valid = _T_7 ^ line_1321_valid_reg;
  assign line_1322_clock = clock;
  assign line_1322_reset = reset;
  assign line_1322_valid = _T_13 ^ line_1322_valid_reg;
  assign line_1323_clock = clock;
  assign line_1323_reset = reset;
  assign line_1323_valid = _T_14 ^ line_1323_valid_reg;
  assign line_1324_clock = clock;
  assign line_1324_reset = reset;
  assign line_1324_valid = _T_13 ^ line_1324_valid_reg;
  assign line_1325_clock = clock;
  assign line_1325_reset = reset;
  assign line_1325_valid = _T_21 ^ line_1325_valid_reg;
  assign line_1326_clock = clock;
  assign line_1326_reset = reset;
  assign line_1326_valid = 4'h0 == auto_out_b_bits_id ^ line_1326_valid_reg;
  assign line_1327_clock = clock;
  assign line_1327_reset = reset;
  assign line_1327_valid = 4'h1 == auto_out_b_bits_id ^ line_1327_valid_reg;
  assign line_1328_clock = clock;
  assign line_1328_reset = reset;
  assign line_1328_valid = 4'h2 == auto_out_b_bits_id ^ line_1328_valid_reg;
  assign line_1329_clock = clock;
  assign line_1329_reset = reset;
  assign line_1329_valid = 4'h3 == auto_out_b_bits_id ^ line_1329_valid_reg;
  assign line_1330_clock = clock;
  assign line_1330_reset = reset;
  assign line_1330_valid = 4'h4 == auto_out_b_bits_id ^ line_1330_valid_reg;
  assign line_1331_clock = clock;
  assign line_1331_reset = reset;
  assign line_1331_valid = 4'h5 == auto_out_b_bits_id ^ line_1331_valid_reg;
  assign line_1332_clock = clock;
  assign line_1332_reset = reset;
  assign line_1332_valid = 4'h6 == auto_out_b_bits_id ^ line_1332_valid_reg;
  assign line_1333_clock = clock;
  assign line_1333_reset = reset;
  assign line_1333_valid = 4'h7 == auto_out_b_bits_id ^ line_1333_valid_reg;
  assign line_1334_clock = clock;
  assign line_1334_reset = reset;
  assign line_1334_valid = 4'h8 == auto_out_b_bits_id ^ line_1334_valid_reg;
  assign line_1335_clock = clock;
  assign line_1335_reset = reset;
  assign line_1335_valid = 4'h9 == auto_out_b_bits_id ^ line_1335_valid_reg;
  assign line_1336_clock = clock;
  assign line_1336_reset = reset;
  assign line_1336_valid = 4'ha == auto_out_b_bits_id ^ line_1336_valid_reg;
  assign line_1337_clock = clock;
  assign line_1337_reset = reset;
  assign line_1337_valid = 4'hb == auto_out_b_bits_id ^ line_1337_valid_reg;
  assign line_1338_clock = clock;
  assign line_1338_reset = reset;
  assign line_1338_valid = 4'hc == auto_out_b_bits_id ^ line_1338_valid_reg;
  assign line_1339_clock = clock;
  assign line_1339_reset = reset;
  assign line_1339_valid = 4'hd == auto_out_b_bits_id ^ line_1339_valid_reg;
  assign line_1340_clock = clock;
  assign line_1340_reset = reset;
  assign line_1340_valid = 4'he == auto_out_b_bits_id ^ line_1340_valid_reg;
  assign line_1341_clock = clock;
  assign line_1341_reset = reset;
  assign line_1341_valid = 4'hf == auto_out_b_bits_id ^ line_1341_valid_reg;
  assign line_1342_clock = clock;
  assign line_1342_reset = reset;
  assign line_1342_valid = _T_41 ^ line_1342_valid_reg;
  assign line_1343_clock = clock;
  assign line_1343_reset = reset;
  assign line_1343_valid = _T_43 ^ line_1343_valid_reg;
  assign line_1344_clock = clock;
  assign line_1344_reset = reset;
  assign line_1344_valid = _T_45 ^ line_1344_valid_reg;
  assign line_1345_clock = clock;
  assign line_1345_reset = reset;
  assign line_1345_valid = _T_47 ^ line_1345_valid_reg;
  assign line_1346_clock = clock;
  assign line_1346_reset = reset;
  assign line_1346_valid = _T_49 ^ line_1346_valid_reg;
  assign line_1347_clock = clock;
  assign line_1347_reset = reset;
  assign line_1347_valid = _T_51 ^ line_1347_valid_reg;
  assign line_1348_clock = clock;
  assign line_1348_reset = reset;
  assign line_1348_valid = _T_53 ^ line_1348_valid_reg;
  assign line_1349_clock = clock;
  assign line_1349_reset = reset;
  assign line_1349_valid = _T_55 ^ line_1349_valid_reg;
  assign line_1350_clock = clock;
  assign line_1350_reset = reset;
  assign line_1350_valid = _T_57 ^ line_1350_valid_reg;
  assign line_1351_clock = clock;
  assign line_1351_reset = reset;
  assign line_1351_valid = _T_59 ^ line_1351_valid_reg;
  assign line_1352_clock = clock;
  assign line_1352_reset = reset;
  assign line_1352_valid = _T_61 ^ line_1352_valid_reg;
  assign line_1353_clock = clock;
  assign line_1353_reset = reset;
  assign line_1353_valid = _T_63 ^ line_1353_valid_reg;
  assign line_1354_clock = clock;
  assign line_1354_reset = reset;
  assign line_1354_valid = _T_65 ^ line_1354_valid_reg;
  assign line_1355_clock = clock;
  assign line_1355_reset = reset;
  assign line_1355_valid = _T_67 ^ line_1355_valid_reg;
  assign line_1356_clock = clock;
  assign line_1356_reset = reset;
  assign line_1356_valid = _T_69 ^ line_1356_valid_reg;
  assign line_1357_clock = clock;
  assign line_1357_reset = reset;
  assign line_1357_valid = _T_71 ^ line_1357_valid_reg;
  assign auto_in_aw_ready = deq_q_1_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_w_ready = in_w_deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_b_valid = auto_out_b_valid & auto_out_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 203:33]
  assign auto_in_b_bits_id = auto_out_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp | _GEN_71; // @[src/main/scala/amba/axi4/Fragmenter.scala 208:41]
  assign auto_in_ar_ready = deq_q_io_enq_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/chisel3/util/Decoupled.scala 385:17]
  assign auto_in_r_valid = auto_out_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_id = auto_out_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 372:12]
  assign auto_in_r_bits_last = auto_out_r_bits_last & auto_out_r_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 194:41]
  assign auto_out_aw_valid = irr_1_valid & _in_aw_ready_T; // @[src/main/scala/amba/axi4/Fragmenter.scala 163:35]
  assign auto_out_aw_bits_id = deq_q_1_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_aw_bits_addr = ~_out_bits_addr_T_12; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:26]
  assign auto_out_aw_bits_echo_real_last = 8'h0 == len_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 114:27]
  assign auto_out_w_valid = in_w_valid & (~w_idle | wbeats_valid); // @[src/main/scala/amba/axi4/Fragmenter.scala 181:33]
  assign auto_out_w_bits_data = in_w_deq_q_io_deq_bits_data; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_w_bits_strb = in_w_deq_q_io_deq_bits_strb; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 204:33]
  assign auto_out_ar_valid = deq_q_io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 422:15]
  assign auto_out_ar_bits_id = deq_q_io_deq_bits_id; // @[src/main/scala/chisel3/util/Decoupled.scala 420:19 421:14]
  assign auto_out_ar_bits_addr = ~_out_bits_addr_T_5; // @[src/main/scala/amba/axi4/Fragmenter.scala 126:26]
  assign auto_out_ar_bits_echo_real_last = 8'h0 == len; // @[src/main/scala/amba/axi4/Fragmenter.scala 114:27]
  assign auto_out_r_ready = auto_in_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_clock = clock;
  assign deq_q_reset = reset;
  assign deq_q_io_enq_valid = auto_in_ar_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_enq_bits_id = auto_in_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_enq_bits_addr = auto_in_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_enq_bits_len = auto_in_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_enq_bits_size = auto_in_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_enq_bits_burst = auto_in_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_io_deq_ready = auto_out_ar_ready & ar_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 115:30]
  assign deq_q_1_clock = clock;
  assign deq_q_1_reset = reset;
  assign deq_q_1_io_enq_valid = auto_in_aw_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_enq_bits_id = auto_in_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_enq_bits_addr = auto_in_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_enq_bits_len = auto_in_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_enq_bits_size = auto_in_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_enq_bits_burst = auto_in_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign deq_q_1_io_deq_ready = in_aw_ready & aw_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 115:30]
  assign in_w_deq_q_clock = clock;
  assign in_w_deq_q_reset = reset;
  assign in_w_deq_q_io_enq_valid = auto_in_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign in_w_deq_q_io_enq_bits_data = auto_in_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign in_w_deq_q_io_enq_bits_strb = auto_in_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign in_w_deq_q_io_enq_bits_last = auto_in_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1214:17 src/main/scala/diplomacy/LazyModule.scala 370:16]
  assign in_w_deq_q_io_deq_ready = auto_out_w_ready & _nodeOut_w_valid_T_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 182:33]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
      busy <= 1'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
    end else if (_T_2) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25]
      busy <= ~ar_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 129:16]
    end
    if (_T_2) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25]
      if (fixed) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 110:60]
        r_addr <= irr_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 111:20]
      end else if (irr_bits_burst == 2'h2) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 107:59]
        r_addr <= _mux_addr_T_4; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:20]
      end else begin
        r_addr <= inc_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 106:35]
      end
    end
    r_len <= _GEN_48[7:0];
    line_1314_valid_reg <= _T;
    line_1315_valid_reg <= fixed;
    line_1316_valid_reg <= _T_2;
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
      busy_1 <= 1'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 64:29]
    end else if (_T_5) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25]
      busy_1 <= ~aw_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 129:16]
    end
    if (_T_5) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 128:25]
      if (fixed_1) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 110:60]
        r_addr_1 <= irr_1_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 111:20]
      end else if (irr_1_bits_burst == 2'h2) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 107:59]
        r_addr_1 <= _mux_addr_T_9; // @[src/main/scala/amba/axi4/Fragmenter.scala 108:20]
      end else begin
        r_addr_1 <= inc_addr_1; // @[src/main/scala/amba/axi4/Fragmenter.scala 106:35]
      end
    end
    r_len_1 <= _GEN_53[7:0];
    line_1317_valid_reg <= _T_3;
    line_1318_valid_reg <= fixed_1;
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 172:30]
      w_counter <= 9'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 172:30]
    end else begin
      w_counter <= _w_counter_T_2; // @[src/main/scala/amba/axi4/Fragmenter.scala 176:17]
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 156:35]
      wbeats_latched <= 1'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 156:35]
    end else if (_T_7) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 160:26]
      wbeats_latched <= 1'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 160:43]
    end else begin
      wbeats_latched <= _GEN_54;
    end
    line_1319_valid_reg <= _T_5;
    line_1320_valid_reg <= _T_6;
    line_1321_valid_reg <= _T_7;
    line_1322_valid_reg <= _T_13;
    line_1323_valid_reg <= _T_14;
    line_1324_valid_reg <= _T_13;
    line_1325_valid_reg <= _T_21;
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_0 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[0] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_0 <= 2'h0;
      end else begin
        error_0 <= _error_0_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_1 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[1] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_1 <= 2'h0;
      end else begin
        error_1 <= _error_1_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_2 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[2] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_2 <= 2'h0;
      end else begin
        error_2 <= _error_2_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_3 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[3] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_3 <= 2'h0;
      end else begin
        error_3 <= _error_3_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_4 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[4] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_4 <= 2'h0;
      end else begin
        error_4 <= _error_4_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_5 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[5] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_5 <= 2'h0;
      end else begin
        error_5 <= _error_5_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_6 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[6] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_6 <= 2'h0;
      end else begin
        error_6 <= _error_6_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_7 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[7] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_7 <= 2'h0;
      end else begin
        error_7 <= _error_7_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_8 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[8] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_8 <= 2'h0;
      end else begin
        error_8 <= _error_8_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_9 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[9] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_9 <= 2'h0;
      end else begin
        error_9 <= _error_9_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_10 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[10] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_10 <= 2'h0;
      end else begin
        error_10 <= _error_10_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_11 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[11] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_11 <= 2'h0;
      end else begin
        error_11 <= _error_11_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_12 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[12] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_12 <= 2'h0;
      end else begin
        error_12 <= _error_12_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_13 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[13] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_13 <= 2'h0;
      end else begin
        error_13 <= _error_13_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_14 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[14] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_14 <= 2'h0;
      end else begin
        error_14 <= _error_14_T;
      end
    end
    if (reset) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
      error_15 <= 2'h0; // @[src/main/scala/amba/axi4/Fragmenter.scala 207:26]
    end else if (_T_22[15] & _T_40) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:34]
      if (auto_out_b_bits_echo_real_last) begin // @[src/main/scala/amba/axi4/Fragmenter.scala 210:46]
        error_15 <= 2'h0;
      end else begin
        error_15 <= _error_15_T;
      end
    end
    line_1326_valid_reg <= 4'h0 == auto_out_b_bits_id;
    line_1327_valid_reg <= 4'h1 == auto_out_b_bits_id;
    line_1328_valid_reg <= 4'h2 == auto_out_b_bits_id;
    line_1329_valid_reg <= 4'h3 == auto_out_b_bits_id;
    line_1330_valid_reg <= 4'h4 == auto_out_b_bits_id;
    line_1331_valid_reg <= 4'h5 == auto_out_b_bits_id;
    line_1332_valid_reg <= 4'h6 == auto_out_b_bits_id;
    line_1333_valid_reg <= 4'h7 == auto_out_b_bits_id;
    line_1334_valid_reg <= 4'h8 == auto_out_b_bits_id;
    line_1335_valid_reg <= 4'h9 == auto_out_b_bits_id;
    line_1336_valid_reg <= 4'ha == auto_out_b_bits_id;
    line_1337_valid_reg <= 4'hb == auto_out_b_bits_id;
    line_1338_valid_reg <= 4'hc == auto_out_b_bits_id;
    line_1339_valid_reg <= 4'hd == auto_out_b_bits_id;
    line_1340_valid_reg <= 4'he == auto_out_b_bits_id;
    line_1341_valid_reg <= 4'hf == auto_out_b_bits_id;
    line_1342_valid_reg <= _T_41;
    line_1343_valid_reg <= _T_43;
    line_1344_valid_reg <= _T_45;
    line_1345_valid_reg <= _T_47;
    line_1346_valid_reg <= _T_49;
    line_1347_valid_reg <= _T_51;
    line_1348_valid_reg <= _T_53;
    line_1349_valid_reg <= _T_55;
    line_1350_valid_reg <= _T_57;
    line_1351_valid_reg <= _T_59;
    line_1352_valid_reg <= _T_61;
    line_1353_valid_reg <= _T_63;
    line_1354_valid_reg <= _T_65;
    line_1355_valid_reg <= _T_67;
    line_1356_valid_reg <= _T_69;
    line_1357_valid_reg <= _T_71;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~_w_counter_T | w_todo != 9'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:177 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n"
            ); // @[src/main/scala/amba/axi4/Fragmenter.scala 177:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~nodeOut_w_valid | ~in_w_bits_last | w_last)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:186 assert (!out.w.valid || !in_w.bits.last || w_last)\n"); // @[src/main/scala/amba/axi4/Fragmenter.scala 186:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  r_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  line_1314_valid_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  line_1315_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  line_1316_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  busy_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_addr_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_len_1 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  line_1317_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_1318_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  w_counter = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  wbeats_latched = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  line_1319_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  line_1320_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  line_1321_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  line_1322_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  line_1323_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  line_1324_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  line_1325_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  error_0 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  error_1 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  error_2 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  error_3 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  error_4 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  error_5 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  error_6 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  error_7 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  error_8 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  error_9 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  error_10 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  error_11 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  error_12 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  error_13 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  error_14 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  error_15 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  line_1326_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  line_1327_valid_reg = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  line_1328_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  line_1329_valid_reg = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  line_1330_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  line_1331_valid_reg = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  line_1332_valid_reg = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  line_1333_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  line_1334_valid_reg = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  line_1335_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  line_1336_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  line_1337_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  line_1338_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  line_1339_valid_reg = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  line_1340_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  line_1341_valid_reg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  line_1342_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  line_1343_valid_reg = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  line_1344_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  line_1345_valid_reg = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  line_1346_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  line_1347_valid_reg = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  line_1348_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  line_1349_valid_reg = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  line_1350_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  line_1351_valid_reg = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  line_1352_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  line_1353_valid_reg = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  line_1354_valid_reg = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  line_1355_valid_reg = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  line_1356_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  line_1357_valid_reg = _RAND_67[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~_w_counter_T | w_todo != 9'h0); // @[src/main/scala/amba/axi4/Fragmenter.scala 177:14]
    end
    //
    if (_T_13) begin
      assert(~nodeOut_w_valid | ~in_w_bits_last | w_last); // @[src/main/scala/amba/axi4/Fragmenter.scala 186:14]
    end
  end
endmodule
module SimAXIMem(
  input         clock,
  input         reset,
  output        io_axi4_0_aw_ready, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_aw_valid, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [3:0]  io_axi4_0_aw_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [31:0] io_axi4_0_aw_bits_addr, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [7:0]  io_axi4_0_aw_bits_len, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [2:0]  io_axi4_0_aw_bits_size, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [1:0]  io_axi4_0_aw_bits_burst, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output        io_axi4_0_w_ready, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_w_valid, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [63:0] io_axi4_0_w_bits_data, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [7:0]  io_axi4_0_w_bits_strb, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_w_bits_last, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_b_ready, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output        io_axi4_0_b_valid, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output [3:0]  io_axi4_0_b_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output [1:0]  io_axi4_0_b_bits_resp, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output        io_axi4_0_ar_ready, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_ar_valid, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [3:0]  io_axi4_0_ar_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [31:0] io_axi4_0_ar_bits_addr, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [7:0]  io_axi4_0_ar_bits_len, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [2:0]  io_axi4_0_ar_bits_size, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input  [1:0]  io_axi4_0_ar_bits_burst, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  input         io_axi4_0_r_ready, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output        io_axi4_0_r_valid, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output [3:0]  io_axi4_0_r_bits_id, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output [63:0] io_axi4_0_r_bits_data, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output [1:0]  io_axi4_0_r_bits_resp, // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
  output        io_axi4_0_r_bits_last // @[src/main/scala/diplomacy/Nodes.scala 1649:17]
);
  wire  srams_clock; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_reset; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_aw_ready; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_aw_valid; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [3:0] srams_auto_in_aw_bits_id; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [31:0] srams_auto_in_aw_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_aw_bits_echo_real_last; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_w_ready; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_w_valid; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [63:0] srams_auto_in_w_bits_data; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [7:0] srams_auto_in_w_bits_strb; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_b_ready; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_b_valid; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [3:0] srams_auto_in_b_bits_id; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [1:0] srams_auto_in_b_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_b_bits_echo_real_last; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_ar_ready; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_ar_valid; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [3:0] srams_auto_in_ar_bits_id; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [31:0] srams_auto_in_ar_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_ar_bits_echo_real_last; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_r_ready; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_r_valid; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [3:0] srams_auto_in_r_bits_id; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [63:0] srams_auto_in_r_bits_data; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire [1:0] srams_auto_in_r_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  srams_auto_in_r_bits_echo_real_last; // @[src/main/scala/system/SimAXIMem.scala 19:15]
  wire  axi4xbar_clock; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_reset; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_aw_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_aw_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [31:0] axi4xbar_auto_in_aw_bits_addr; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_in_aw_bits_len; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [2:0] axi4xbar_auto_in_aw_bits_size; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_in_aw_bits_burst; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_w_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_w_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [63:0] axi4xbar_auto_in_w_bits_data; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_in_w_bits_strb; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_w_bits_last; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_b_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_b_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_in_b_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_in_b_bits_resp; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_ar_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_ar_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [31:0] axi4xbar_auto_in_ar_bits_addr; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_in_ar_bits_len; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [2:0] axi4xbar_auto_in_ar_bits_size; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_in_ar_bits_burst; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_r_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_r_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_in_r_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [63:0] axi4xbar_auto_in_r_bits_data; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_in_r_bits_resp; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_in_r_bits_last; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_aw_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_aw_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_out_aw_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [31:0] axi4xbar_auto_out_aw_bits_addr; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_out_aw_bits_len; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [2:0] axi4xbar_auto_out_aw_bits_size; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_out_aw_bits_burst; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_w_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_w_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [63:0] axi4xbar_auto_out_w_bits_data; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_out_w_bits_strb; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_w_bits_last; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_b_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_b_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_out_b_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_ar_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_ar_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_out_ar_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [31:0] axi4xbar_auto_out_ar_bits_addr; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [7:0] axi4xbar_auto_out_ar_bits_len; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [2:0] axi4xbar_auto_out_ar_bits_size; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_out_ar_bits_burst; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_r_ready; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_r_valid; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [3:0] axi4xbar_auto_out_r_bits_id; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [63:0] axi4xbar_auto_out_r_bits_data; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire [1:0] axi4xbar_auto_out_r_bits_resp; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4xbar_auto_out_r_bits_last; // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
  wire  axi4buf_clock; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_reset; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [31:0] axi4buf_auto_in_aw_bits_addr; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_aw_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_w_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_w_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_in_w_bits_data; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_in_w_bits_strb; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_b_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_b_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_b_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [31:0] axi4buf_auto_in_ar_bits_addr; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_ar_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_in_r_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_in_r_bits_data; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_in_r_bits_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_aw_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [31:0] axi4buf_auto_out_aw_bits_addr; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_aw_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_w_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_w_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_out_w_bits_data; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [7:0] axi4buf_auto_out_w_bits_strb; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_b_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_b_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_b_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_ar_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [31:0] axi4buf_auto_out_ar_bits_addr; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_ar_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_ready; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_valid; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [3:0] axi4buf_auto_out_r_bits_id; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [63:0] axi4buf_auto_out_r_bits_data; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire [1:0] axi4buf_auto_out_r_bits_resp; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4buf_auto_out_r_bits_echo_real_last; // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
  wire  axi4frag_clock; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_reset; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_aw_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_aw_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_in_aw_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [31:0] axi4frag_auto_in_aw_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [7:0] axi4frag_auto_in_aw_bits_len; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [2:0] axi4frag_auto_in_aw_bits_size; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_in_aw_bits_burst; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_w_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_w_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [63:0] axi4frag_auto_in_w_bits_data; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [7:0] axi4frag_auto_in_w_bits_strb; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_w_bits_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_b_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_b_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_in_b_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_in_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_ar_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_ar_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_in_ar_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [31:0] axi4frag_auto_in_ar_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [7:0] axi4frag_auto_in_ar_bits_len; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [2:0] axi4frag_auto_in_ar_bits_size; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_in_ar_bits_burst; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_r_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_r_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_in_r_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [63:0] axi4frag_auto_in_r_bits_data; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_in_r_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_in_r_bits_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_aw_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_aw_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_out_aw_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [31:0] axi4frag_auto_out_aw_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_aw_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_w_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_w_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [63:0] axi4frag_auto_out_w_bits_data; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [7:0] axi4frag_auto_out_w_bits_strb; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_b_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_b_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_out_b_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_out_b_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_b_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_ar_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_ar_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_out_ar_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [31:0] axi4frag_auto_out_ar_bits_addr; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_ar_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_r_ready; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_r_valid; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [3:0] axi4frag_auto_out_r_bits_id; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [63:0] axi4frag_auto_out_r_bits_data; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire [1:0] axi4frag_auto_out_r_bits_resp; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_r_bits_echo_real_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  wire  axi4frag_auto_out_r_bits_last; // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
  AXI4RAM srams ( // @[src/main/scala/system/SimAXIMem.scala 19:15]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_aw_ready(srams_auto_in_aw_ready),
    .auto_in_aw_valid(srams_auto_in_aw_valid),
    .auto_in_aw_bits_id(srams_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(srams_auto_in_aw_bits_addr),
    .auto_in_aw_bits_echo_real_last(srams_auto_in_aw_bits_echo_real_last),
    .auto_in_w_ready(srams_auto_in_w_ready),
    .auto_in_w_valid(srams_auto_in_w_valid),
    .auto_in_w_bits_data(srams_auto_in_w_bits_data),
    .auto_in_w_bits_strb(srams_auto_in_w_bits_strb),
    .auto_in_b_ready(srams_auto_in_b_ready),
    .auto_in_b_valid(srams_auto_in_b_valid),
    .auto_in_b_bits_id(srams_auto_in_b_bits_id),
    .auto_in_b_bits_resp(srams_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_real_last(srams_auto_in_b_bits_echo_real_last),
    .auto_in_ar_ready(srams_auto_in_ar_ready),
    .auto_in_ar_valid(srams_auto_in_ar_valid),
    .auto_in_ar_bits_id(srams_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(srams_auto_in_ar_bits_addr),
    .auto_in_ar_bits_echo_real_last(srams_auto_in_ar_bits_echo_real_last),
    .auto_in_r_ready(srams_auto_in_r_ready),
    .auto_in_r_valid(srams_auto_in_r_valid),
    .auto_in_r_bits_id(srams_auto_in_r_bits_id),
    .auto_in_r_bits_data(srams_auto_in_r_bits_data),
    .auto_in_r_bits_resp(srams_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_real_last(srams_auto_in_r_bits_echo_real_last)
  );
  AXI4Xbar axi4xbar ( // @[src/main/scala/amba/axi4/Xbar.scala 230:30]
    .clock(axi4xbar_clock),
    .reset(axi4xbar_reset),
    .auto_in_aw_ready(axi4xbar_auto_in_aw_ready),
    .auto_in_aw_valid(axi4xbar_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4xbar_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4xbar_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4xbar_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4xbar_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4xbar_auto_in_aw_bits_burst),
    .auto_in_w_ready(axi4xbar_auto_in_w_ready),
    .auto_in_w_valid(axi4xbar_auto_in_w_valid),
    .auto_in_w_bits_data(axi4xbar_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4xbar_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4xbar_auto_in_w_bits_last),
    .auto_in_b_ready(axi4xbar_auto_in_b_ready),
    .auto_in_b_valid(axi4xbar_auto_in_b_valid),
    .auto_in_b_bits_id(axi4xbar_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4xbar_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4xbar_auto_in_ar_ready),
    .auto_in_ar_valid(axi4xbar_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4xbar_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4xbar_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4xbar_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4xbar_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4xbar_auto_in_ar_bits_burst),
    .auto_in_r_ready(axi4xbar_auto_in_r_ready),
    .auto_in_r_valid(axi4xbar_auto_in_r_valid),
    .auto_in_r_bits_id(axi4xbar_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4xbar_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4xbar_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4xbar_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4xbar_auto_out_aw_ready),
    .auto_out_aw_valid(axi4xbar_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4xbar_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4xbar_auto_out_aw_bits_addr),
    .auto_out_aw_bits_len(axi4xbar_auto_out_aw_bits_len),
    .auto_out_aw_bits_size(axi4xbar_auto_out_aw_bits_size),
    .auto_out_aw_bits_burst(axi4xbar_auto_out_aw_bits_burst),
    .auto_out_w_ready(axi4xbar_auto_out_w_ready),
    .auto_out_w_valid(axi4xbar_auto_out_w_valid),
    .auto_out_w_bits_data(axi4xbar_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4xbar_auto_out_w_bits_strb),
    .auto_out_w_bits_last(axi4xbar_auto_out_w_bits_last),
    .auto_out_b_ready(axi4xbar_auto_out_b_ready),
    .auto_out_b_valid(axi4xbar_auto_out_b_valid),
    .auto_out_b_bits_id(axi4xbar_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4xbar_auto_out_b_bits_resp),
    .auto_out_ar_ready(axi4xbar_auto_out_ar_ready),
    .auto_out_ar_valid(axi4xbar_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4xbar_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4xbar_auto_out_ar_bits_addr),
    .auto_out_ar_bits_len(axi4xbar_auto_out_ar_bits_len),
    .auto_out_ar_bits_size(axi4xbar_auto_out_ar_bits_size),
    .auto_out_ar_bits_burst(axi4xbar_auto_out_ar_bits_burst),
    .auto_out_r_ready(axi4xbar_auto_out_r_ready),
    .auto_out_r_valid(axi4xbar_auto_out_r_valid),
    .auto_out_r_bits_id(axi4xbar_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4xbar_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4xbar_auto_out_r_bits_resp),
    .auto_out_r_bits_last(axi4xbar_auto_out_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[src/main/scala/amba/axi4/Buffer.scala 63:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_echo_real_last(axi4buf_auto_in_aw_bits_echo_real_last),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_b_bits_echo_real_last(axi4buf_auto_in_b_bits_echo_real_last),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_echo_real_last(axi4buf_auto_in_ar_bits_echo_real_last),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_echo_real_last(axi4buf_auto_in_r_bits_echo_real_last),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_aw_bits_echo_real_last(axi4buf_auto_out_aw_bits_echo_real_last),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4buf_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_real_last(axi4buf_auto_out_b_bits_echo_real_last),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_echo_real_last(axi4buf_auto_out_ar_bits_echo_real_last),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4buf_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_real_last(axi4buf_auto_out_r_bits_echo_real_last)
  );
  AXI4Fragmenter axi4frag ( // @[src/main/scala/amba/axi4/Fragmenter.scala 220:30]
    .clock(axi4frag_clock),
    .reset(axi4frag_reset),
    .auto_in_aw_ready(axi4frag_auto_in_aw_ready),
    .auto_in_aw_valid(axi4frag_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4frag_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4frag_auto_in_aw_bits_addr),
    .auto_in_aw_bits_len(axi4frag_auto_in_aw_bits_len),
    .auto_in_aw_bits_size(axi4frag_auto_in_aw_bits_size),
    .auto_in_aw_bits_burst(axi4frag_auto_in_aw_bits_burst),
    .auto_in_w_ready(axi4frag_auto_in_w_ready),
    .auto_in_w_valid(axi4frag_auto_in_w_valid),
    .auto_in_w_bits_data(axi4frag_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4frag_auto_in_w_bits_strb),
    .auto_in_w_bits_last(axi4frag_auto_in_w_bits_last),
    .auto_in_b_ready(axi4frag_auto_in_b_ready),
    .auto_in_b_valid(axi4frag_auto_in_b_valid),
    .auto_in_b_bits_id(axi4frag_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4frag_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4frag_auto_in_ar_ready),
    .auto_in_ar_valid(axi4frag_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4frag_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4frag_auto_in_ar_bits_addr),
    .auto_in_ar_bits_len(axi4frag_auto_in_ar_bits_len),
    .auto_in_ar_bits_size(axi4frag_auto_in_ar_bits_size),
    .auto_in_ar_bits_burst(axi4frag_auto_in_ar_bits_burst),
    .auto_in_r_ready(axi4frag_auto_in_r_ready),
    .auto_in_r_valid(axi4frag_auto_in_r_valid),
    .auto_in_r_bits_id(axi4frag_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4frag_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4frag_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4frag_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4frag_auto_out_aw_ready),
    .auto_out_aw_valid(axi4frag_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4frag_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4frag_auto_out_aw_bits_addr),
    .auto_out_aw_bits_echo_real_last(axi4frag_auto_out_aw_bits_echo_real_last),
    .auto_out_w_ready(axi4frag_auto_out_w_ready),
    .auto_out_w_valid(axi4frag_auto_out_w_valid),
    .auto_out_w_bits_data(axi4frag_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4frag_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4frag_auto_out_b_ready),
    .auto_out_b_valid(axi4frag_auto_out_b_valid),
    .auto_out_b_bits_id(axi4frag_auto_out_b_bits_id),
    .auto_out_b_bits_resp(axi4frag_auto_out_b_bits_resp),
    .auto_out_b_bits_echo_real_last(axi4frag_auto_out_b_bits_echo_real_last),
    .auto_out_ar_ready(axi4frag_auto_out_ar_ready),
    .auto_out_ar_valid(axi4frag_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4frag_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4frag_auto_out_ar_bits_addr),
    .auto_out_ar_bits_echo_real_last(axi4frag_auto_out_ar_bits_echo_real_last),
    .auto_out_r_ready(axi4frag_auto_out_r_ready),
    .auto_out_r_valid(axi4frag_auto_out_r_valid),
    .auto_out_r_bits_id(axi4frag_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4frag_auto_out_r_bits_data),
    .auto_out_r_bits_resp(axi4frag_auto_out_r_bits_resp),
    .auto_out_r_bits_echo_real_last(axi4frag_auto_out_r_bits_echo_real_last),
    .auto_out_r_bits_last(axi4frag_auto_out_r_bits_last)
  );
  assign io_axi4_0_aw_ready = axi4xbar_auto_in_aw_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_w_ready = axi4xbar_auto_in_w_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_b_valid = axi4xbar_auto_in_b_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_b_bits_id = axi4xbar_auto_in_b_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_b_bits_resp = axi4xbar_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_ar_ready = axi4xbar_auto_in_ar_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_r_valid = axi4xbar_auto_in_r_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_r_bits_id = axi4xbar_auto_in_r_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_r_bits_data = axi4xbar_auto_in_r_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_r_bits_resp = axi4xbar_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign io_axi4_0_r_bits_last = axi4xbar_auto_in_r_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign srams_clock = clock;
  assign srams_reset = reset;
  assign srams_auto_in_aw_valid = axi4buf_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_aw_bits_echo_real_last = axi4buf_auto_out_aw_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_w_valid = axi4buf_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_b_ready = axi4buf_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_ar_valid = axi4buf_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_ar_bits_echo_real_last = axi4buf_auto_out_ar_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign srams_auto_in_r_ready = axi4buf_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4xbar_clock = clock;
  assign axi4xbar_reset = reset;
  assign axi4xbar_auto_in_aw_valid = io_axi4_0_aw_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_aw_bits_id = io_axi4_0_aw_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_aw_bits_addr = io_axi4_0_aw_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_aw_bits_len = io_axi4_0_aw_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_aw_bits_size = io_axi4_0_aw_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_aw_bits_burst = io_axi4_0_aw_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_w_valid = io_axi4_0_w_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_w_bits_data = io_axi4_0_w_bits_data; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_w_bits_strb = io_axi4_0_w_bits_strb; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_w_bits_last = io_axi4_0_w_bits_last; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_b_ready = io_axi4_0_b_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_valid = io_axi4_0_ar_valid; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_bits_id = io_axi4_0_ar_bits_id; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_bits_addr = io_axi4_0_ar_bits_addr; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_bits_len = io_axi4_0_ar_bits_len; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_bits_size = io_axi4_0_ar_bits_size; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_ar_bits_burst = io_axi4_0_ar_bits_burst; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_in_r_ready = io_axi4_0_r_ready; // @[src/main/scala/diplomacy/Nodes.scala 1205:17 1651:60]
  assign axi4xbar_auto_out_aw_ready = axi4frag_auto_in_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_w_ready = axi4frag_auto_in_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_b_valid = axi4frag_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_b_bits_id = axi4frag_auto_in_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_b_bits_resp = axi4frag_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_ar_ready = axi4frag_auto_in_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_r_valid = axi4frag_auto_in_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_r_bits_id = axi4frag_auto_in_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_r_bits_data = axi4frag_auto_in_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_r_bits_resp = axi4frag_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4xbar_auto_out_r_bits_last = axi4frag_auto_in_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = axi4frag_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_aw_bits_id = axi4frag_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_aw_bits_addr = axi4frag_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_aw_bits_echo_real_last = axi4frag_auto_out_aw_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_w_valid = axi4frag_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_w_bits_data = axi4frag_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_w_bits_strb = axi4frag_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_b_ready = axi4frag_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_ar_valid = axi4frag_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_ar_bits_id = axi4frag_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_ar_bits_addr = axi4frag_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_ar_bits_echo_real_last = axi4frag_auto_out_ar_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_in_r_ready = axi4frag_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_aw_ready = srams_auto_in_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_w_ready = srams_auto_in_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_b_valid = srams_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_b_bits_id = srams_auto_in_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_b_bits_resp = srams_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_b_bits_echo_real_last = srams_auto_in_b_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_ar_ready = srams_auto_in_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_r_valid = srams_auto_in_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_r_bits_id = srams_auto_in_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_r_bits_data = srams_auto_in_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_r_bits_resp = srams_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4buf_auto_out_r_bits_echo_real_last = srams_auto_in_r_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_clock = clock;
  assign axi4frag_reset = reset;
  assign axi4frag_auto_in_aw_valid = axi4xbar_auto_out_aw_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_aw_bits_id = axi4xbar_auto_out_aw_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_aw_bits_addr = axi4xbar_auto_out_aw_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_aw_bits_len = axi4xbar_auto_out_aw_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_aw_bits_size = axi4xbar_auto_out_aw_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_aw_bits_burst = axi4xbar_auto_out_aw_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_w_valid = axi4xbar_auto_out_w_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_w_bits_data = axi4xbar_auto_out_w_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_w_bits_strb = axi4xbar_auto_out_w_bits_strb; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_w_bits_last = axi4xbar_auto_out_w_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_b_ready = axi4xbar_auto_out_b_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_valid = axi4xbar_auto_out_ar_valid; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_bits_id = axi4xbar_auto_out_ar_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_bits_addr = axi4xbar_auto_out_ar_bits_addr; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_bits_len = axi4xbar_auto_out_ar_bits_len; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_bits_size = axi4xbar_auto_out_ar_bits_size; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_ar_bits_burst = axi4xbar_auto_out_ar_bits_burst; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_in_r_ready = axi4xbar_auto_out_r_ready; // @[src/main/scala/diplomacy/LazyModule.scala 357:18]
  assign axi4frag_auto_out_aw_ready = axi4buf_auto_in_aw_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_w_ready = axi4buf_auto_in_w_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_b_valid = axi4buf_auto_in_b_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_b_bits_id = axi4buf_auto_in_b_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_b_bits_echo_real_last = axi4buf_auto_in_b_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_ar_ready = axi4buf_auto_in_ar_ready; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_valid = axi4buf_auto_in_r_valid; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_bits_id = axi4buf_auto_in_r_bits_id; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_bits_data = axi4buf_auto_in_r_bits_data; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_bits_echo_real_last = axi4buf_auto_in_r_bits_echo_real_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
  assign axi4frag_auto_out_r_bits_last = axi4buf_auto_in_r_bits_last; // @[src/main/scala/diplomacy/LazyModule.scala 355:18]
endmodule
module SimTop(
  input         clock,
  input         reset,
  output [63:0] difftest_exit, // @[difftest/src/main/scala/Difftest.scala 502:22]
  output [63:0] difftest_step, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input         difftest_perfCtrl_clean, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input         difftest_perfCtrl_dump, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input  [63:0] difftest_logCtrl_begin, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input  [63:0] difftest_logCtrl_end, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input  [63:0] difftest_logCtrl_level, // @[difftest/src/main/scala/Difftest.scala 502:22]
  output        difftest_uart_out_valid, // @[difftest/src/main/scala/Difftest.scala 502:22]
  output [7:0]  difftest_uart_out_ch, // @[difftest/src/main/scala/Difftest.scala 502:22]
  output        difftest_uart_in_valid, // @[difftest/src/main/scala/Difftest.scala 502:22]
  input  [7:0]  difftest_uart_in_ch // @[difftest/src/main/scala/Difftest.scala 502:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  ldut_clock; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_reset; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_aw_ready; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_aw_valid; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [3:0] ldut_mem_axi4_0_aw_bits_id; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [31:0] ldut_mem_axi4_0_aw_bits_addr; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [7:0] ldut_mem_axi4_0_aw_bits_len; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [2:0] ldut_mem_axi4_0_aw_bits_size; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [1:0] ldut_mem_axi4_0_aw_bits_burst; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_w_ready; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_w_valid; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [63:0] ldut_mem_axi4_0_w_bits_data; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [7:0] ldut_mem_axi4_0_w_bits_strb; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_w_bits_last; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_b_ready; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_b_valid; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [3:0] ldut_mem_axi4_0_b_bits_id; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [1:0] ldut_mem_axi4_0_b_bits_resp; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_ar_ready; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_ar_valid; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [3:0] ldut_mem_axi4_0_ar_bits_id; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [31:0] ldut_mem_axi4_0_ar_bits_addr; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [7:0] ldut_mem_axi4_0_ar_bits_len; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [2:0] ldut_mem_axi4_0_ar_bits_size; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [1:0] ldut_mem_axi4_0_ar_bits_burst; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_r_ready; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_r_valid; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [3:0] ldut_mem_axi4_0_r_bits_id; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [63:0] ldut_mem_axi4_0_r_bits_data; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire [1:0] ldut_mem_axi4_0_r_bits_resp; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  ldut_mem_axi4_0_r_bits_last; // @[src/main/scala/system/FuzzHarness.scala 28:19]
  wire  mem_clock; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_reset; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_aw_ready; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_aw_valid; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [3:0] mem_io_axi4_0_aw_bits_id; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [31:0] mem_io_axi4_0_aw_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [7:0] mem_io_axi4_0_aw_bits_len; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [2:0] mem_io_axi4_0_aw_bits_size; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [1:0] mem_io_axi4_0_aw_bits_burst; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_w_ready; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_w_valid; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [63:0] mem_io_axi4_0_w_bits_data; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [7:0] mem_io_axi4_0_w_bits_strb; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_w_bits_last; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_b_ready; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_b_valid; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [3:0] mem_io_axi4_0_b_bits_id; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [1:0] mem_io_axi4_0_b_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_ar_ready; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_ar_valid; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [3:0] mem_io_axi4_0_ar_bits_id; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [31:0] mem_io_axi4_0_ar_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [7:0] mem_io_axi4_0_ar_bits_len; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [2:0] mem_io_axi4_0_ar_bits_size; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [1:0] mem_io_axi4_0_ar_bits_burst; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_r_ready; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_r_valid; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [3:0] mem_io_axi4_0_r_bits_id; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [63:0] mem_io_axi4_0_r_bits_data; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire [1:0] mem_io_axi4_0_r_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  wire  mem_io_axi4_0_r_bits_last; // @[src/main/scala/system/SimAXIMem.scala 47:13]
  reg [63:0] difftest_timer; // @[difftest/src/main/scala/Difftest.scala 507:24]
  wire [63:0] _difftest_timer_T_1 = difftest_timer + 64'h1; // @[difftest/src/main/scala/Difftest.scala 508:20]
  wire  difftest_log_enable = difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end; // @[difftest/src/main/scala/Difftest.scala 656:26]
  ExampleFuzzSystem ldut ( // @[src/main/scala/system/FuzzHarness.scala 28:19]
    .clock(ldut_clock),
    .reset(ldut_reset),
    .mem_axi4_0_aw_ready(ldut_mem_axi4_0_aw_ready),
    .mem_axi4_0_aw_valid(ldut_mem_axi4_0_aw_valid),
    .mem_axi4_0_aw_bits_id(ldut_mem_axi4_0_aw_bits_id),
    .mem_axi4_0_aw_bits_addr(ldut_mem_axi4_0_aw_bits_addr),
    .mem_axi4_0_aw_bits_len(ldut_mem_axi4_0_aw_bits_len),
    .mem_axi4_0_aw_bits_size(ldut_mem_axi4_0_aw_bits_size),
    .mem_axi4_0_aw_bits_burst(ldut_mem_axi4_0_aw_bits_burst),
    .mem_axi4_0_w_ready(ldut_mem_axi4_0_w_ready),
    .mem_axi4_0_w_valid(ldut_mem_axi4_0_w_valid),
    .mem_axi4_0_w_bits_data(ldut_mem_axi4_0_w_bits_data),
    .mem_axi4_0_w_bits_strb(ldut_mem_axi4_0_w_bits_strb),
    .mem_axi4_0_w_bits_last(ldut_mem_axi4_0_w_bits_last),
    .mem_axi4_0_b_ready(ldut_mem_axi4_0_b_ready),
    .mem_axi4_0_b_valid(ldut_mem_axi4_0_b_valid),
    .mem_axi4_0_b_bits_id(ldut_mem_axi4_0_b_bits_id),
    .mem_axi4_0_b_bits_resp(ldut_mem_axi4_0_b_bits_resp),
    .mem_axi4_0_ar_ready(ldut_mem_axi4_0_ar_ready),
    .mem_axi4_0_ar_valid(ldut_mem_axi4_0_ar_valid),
    .mem_axi4_0_ar_bits_id(ldut_mem_axi4_0_ar_bits_id),
    .mem_axi4_0_ar_bits_addr(ldut_mem_axi4_0_ar_bits_addr),
    .mem_axi4_0_ar_bits_len(ldut_mem_axi4_0_ar_bits_len),
    .mem_axi4_0_ar_bits_size(ldut_mem_axi4_0_ar_bits_size),
    .mem_axi4_0_ar_bits_burst(ldut_mem_axi4_0_ar_bits_burst),
    .mem_axi4_0_r_ready(ldut_mem_axi4_0_r_ready),
    .mem_axi4_0_r_valid(ldut_mem_axi4_0_r_valid),
    .mem_axi4_0_r_bits_id(ldut_mem_axi4_0_r_bits_id),
    .mem_axi4_0_r_bits_data(ldut_mem_axi4_0_r_bits_data),
    .mem_axi4_0_r_bits_resp(ldut_mem_axi4_0_r_bits_resp),
    .mem_axi4_0_r_bits_last(ldut_mem_axi4_0_r_bits_last)
  );
  SimAXIMem mem ( // @[src/main/scala/system/SimAXIMem.scala 47:13]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_axi4_0_aw_ready(mem_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(mem_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(mem_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(mem_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(mem_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(mem_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(mem_io_axi4_0_aw_bits_burst),
    .io_axi4_0_w_ready(mem_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(mem_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(mem_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(mem_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(mem_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(mem_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(mem_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(mem_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(mem_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(mem_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(mem_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(mem_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(mem_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(mem_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(mem_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(mem_io_axi4_0_ar_bits_burst),
    .io_axi4_0_r_ready(mem_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(mem_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(mem_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(mem_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(mem_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(mem_io_axi4_0_r_bits_last)
  );
  assign difftest_exit = 64'h0; // @[difftest/src/main/scala/Difftest.scala 504:19]
  assign difftest_step = 64'h1; // @[difftest/src/main/scala/Difftest.scala 505:19]
  assign difftest_uart_out_valid = 1'h0;
  assign difftest_uart_out_ch = 8'h0;
  assign difftest_uart_in_valid = 1'h0;
  assign ldut_clock = clock;
  assign ldut_reset = reset; // @[src/main/scala/system/FuzzHarness.scala 31:109]
  assign ldut_mem_axi4_0_aw_ready = mem_io_axi4_0_aw_ready; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_w_ready = mem_io_axi4_0_w_ready; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_b_valid = mem_io_axi4_0_b_valid; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_b_bits_id = mem_io_axi4_0_b_bits_id; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_b_bits_resp = mem_io_axi4_0_b_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_ar_ready = mem_io_axi4_0_ar_ready; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_r_valid = mem_io_axi4_0_r_valid; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_r_bits_id = mem_io_axi4_0_r_bits_id; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_r_bits_data = mem_io_axi4_0_r_bits_data; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_r_bits_resp = mem_io_axi4_0_r_bits_resp; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign ldut_mem_axi4_0_r_bits_last = mem_io_axi4_0_r_bits_last; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_axi4_0_aw_valid = ldut_mem_axi4_0_aw_valid; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_aw_bits_id = ldut_mem_axi4_0_aw_bits_id; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_aw_bits_addr = ldut_mem_axi4_0_aw_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_aw_bits_len = ldut_mem_axi4_0_aw_bits_len; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_aw_bits_size = ldut_mem_axi4_0_aw_bits_size; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_aw_bits_burst = ldut_mem_axi4_0_aw_bits_burst; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_w_valid = ldut_mem_axi4_0_w_valid; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_w_bits_data = ldut_mem_axi4_0_w_bits_data; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_w_bits_strb = ldut_mem_axi4_0_w_bits_strb; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_w_bits_last = ldut_mem_axi4_0_w_bits_last; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_b_ready = ldut_mem_axi4_0_b_ready; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_valid = ldut_mem_axi4_0_ar_valid; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_bits_id = ldut_mem_axi4_0_ar_bits_id; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_bits_addr = ldut_mem_axi4_0_ar_bits_addr; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_bits_len = ldut_mem_axi4_0_ar_bits_len; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_bits_size = ldut_mem_axi4_0_ar_bits_size; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_ar_bits_burst = ldut_mem_axi4_0_ar_bits_burst; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  assign mem_io_axi4_0_r_ready = ldut_mem_axi4_0_r_ready; // @[src/main/scala/system/SimAXIMem.scala 48:24]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/Difftest.scala 507:24]
      difftest_timer <= 64'h0; // @[difftest/src/main/scala/Difftest.scala 507:24]
    end else begin
      difftest_timer <= _difftest_timer_T_1; // @[difftest/src/main/scala/Difftest.scala 508:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_timer = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
