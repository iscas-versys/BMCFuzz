module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [28:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [1:0]  io_r_resp_data_0__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [38:0] io_r_resp_data_0_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [2:0]  io_r_resp_data_0_brIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [28:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [1:0]  io_w_req_bits_data__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [38:0] io_w_req_bits_data_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [2:0]  io_w_req_bits_data_brIdx // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_0_R0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_R0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_W0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_W0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire [73:0] _wdataword_T = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,
    io_w_req_bits_data_brIdx,1'h1}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  reg  rdata_REG; // @[src/main/scala/utils/Hold.scala 28:106]
  reg [73:0] rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [73:0] _GEN_14 = rdata_REG ? array_0_R0_data : rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  array_0 array_0 ( // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    .R0_addr(array_0_R0_addr),
    .R0_en(array_0_R0_en),
    .R0_clk(array_0_R0_clk),
    .R0_data(array_0_R0_data),
    .W0_addr(array_0_W0_addr),
    .W0_en(array_0_W0_en),
    .W0_clk(array_0_W0_clk),
    .W0_data(array_0_W0_data)
  );
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _GEN_14[73:45]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0__type = _GEN_14[44:43]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_target = _GEN_14[42:4]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_brIdx = _GEN_14[3:1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _GEN_14[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign array_0_R0_addr = io_r_req_bits_setIdx; // @[src/main/scala/utils/Hold.scala 28:87]
  assign array_0_R0_en = io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
  assign array_0_R0_clk = clock; // @[src/main/scala/utils/Hold.scala 28:{87,87}]
  assign array_0_W0_addr = resetState ? resetSet : io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 91:19]
  assign array_0_W0_en = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  assign array_0_W0_clk = clock; // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
  assign array_0_W0_data = resetState ? 74'h0 : _wdataword_T; // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
  always @(posedge clock) begin
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    rdata_REG <= io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= 74'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (rdata_REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= array_0_R0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  rdata_REG = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  rdata_r_0 = _RAND_3[73:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input  [38:0] io_in_pc_bits, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [38:0] io_out_target, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [2:0]  io_brIdx, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_crosslineJump, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushICache,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_reset; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  reg [38:0] ras [0:15]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_rasTarget_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_rasTarget_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_MPORT_1_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  reg  flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire [28:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  _btbHit_T_7 = btb_io_r_req_ready & btb_io_r_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:10] & ~flush & btbHit_REG & ~(pcLatch[1] & btbRead_brIdx[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  reg [3:0] sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [38:0] rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire  _btbWrite_brIdx_T_3 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/BPU.scala 367:46]
  wire  _btbWrite_brIdx_T_6 = ~bpuUpdateReq_pc[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 367:72]
  wire [1:0] btbWrite_brIdx_hi = {_btbWrite_brIdx_T_3,bpuUpdateReq_pc[1]}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  wire  _T_27 = bpuUpdateReq_fuOpType == 7'h5c; // @[src/main/scala/nutcore/frontend/BPU.scala 403:24]
  wire [3:0] _T_29 = sp_value + 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 404:26]
  wire [38:0] _T_31 = bpuUpdateReq_pc + 39'h2; // @[src/main/scala/nutcore/frontend/BPU.scala 404:55]
  wire [38:0] _T_33 = bpuUpdateReq_pc + 39'h4; // @[src/main/scala/nutcore/frontend/BPU.scala 404:69]
  wire [3:0] _value_T_4 = sp_value - 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 412:53]
  wire [3:0] _value_T_5 = sp_value == 4'h0 ? 4'h0 : _value_T_4; // @[src/main/scala/nutcore/frontend/BPU.scala 412:22]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [1:0] _io_brIdx_T = io_out_valid ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 419:63]
  wire [3:0] _io_brIdx_T_1 = {1'h1,crosslineJump,_io_brIdx_T}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:35]
  wire [3:0] _GEN_3 = {{1'd0}, btbRead_brIdx}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  wire [3:0] _io_brIdx_T_2 = _GEN_3 & _io_brIdx_T_1; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  SRAMTemplate btb ( // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  assign ras_rasTarget_MPORT_en = 1'h1;
  assign ras_rasTarget_MPORT_addr = sp_value;
  assign ras_rasTarget_MPORT_data = ras[ras_rasTarget_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  assign ras_MPORT_1_data = bpuUpdateReq_isRVC ? _T_31 : _T_33;
  assign ras_MPORT_1_addr = sp_value + 4'h1;
  assign ras_MPORT_1_mask = 1'h1;
  assign ras_MPORT_1_en = bpuUpdateReq_valid & _T_27;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[src/main/scala/nutcore/frontend/BPU.scala 416:23]
  assign io_out_valid = 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 420:16]
  assign io_brIdx = _io_brIdx_T_2[2:0]; // @[src/main/scala/nutcore/frontend/BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 375:43]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:10]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_brIdx = {btbWrite_brIdx_hi,_btbWrite_brIdx_T_6}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  always @(posedge clock) begin
    if (ras_MPORT_1_en & ras_MPORT_1_mask) begin
      ras[ras_MPORT_1_addr] <= ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      flush <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
      pcLatch <= io_in_pc_bits; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
      btbHit_REG <= 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end else begin
      btbHit_REG <= _btbHit_T_7; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      sp_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        sp_value <= _T_29; // @[src/main/scala/nutcore/frontend/BPU.scala 406:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[src/main/scala/nutcore/frontend/BPU.scala 408:48]
        sp_value <= _value_T_5; // @[src/main/scala/nutcore/frontend/BPU.scala 412:16]
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      rasTarget <= ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_0[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flush = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  pcLatch = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  btbHit_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sp_value = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  rasTarget = _RAND_5[38:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [81:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [81:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input         flushICache,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_reset; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_in_pc_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_in_pc_bits; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_out_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [2:0] bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_crosslineJump; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushICache; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushTLB; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  reg [38:0] pc; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
  wire  _pcUpdate_T = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  pcUpdate = io_redirect_valid | _pcUpdate_T; // @[src/main/scala/nutcore/frontend/IFU.scala 324:36]
  wire [38:0] _snpc_T_2 = pc + 39'h2; // @[src/main/scala/nutcore/frontend/IFU.scala 325:28]
  wire [38:0] _snpc_T_4 = pc + 39'h4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:38]
  wire [38:0] snpc = pc[1] ? _snpc_T_2 : _snpc_T_4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:17]
  reg  crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
  reg [38:0] crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
  wire [38:0] _npc_T_1 = crosslineJumpLatch ? crosslineJumpTarget : snpc; // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  wire  _npcIsSeq_T_2 = crosslineJumpLatch ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/frontend/IFU.scala 342:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _npcIsSeq_T_2; // @[src/main/scala/nutcore/frontend/IFU.scala 342:21]
  wire [2:0] _brIdx_T = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 350:29]
  wire [42:0] x8_hi = {npcIsSeq,_brIdx_T,npc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  wire  _T_3 = io_imem_resp_ready & io_imem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_4 = |io_flushVec; // @[src/main/scala/nutcore/frontend/IFU.scala 396:37]
  BPU_inorder bp1 ( // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushICache(bp1_MOUFlushICache),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[src/main/scala/nutcore/frontend/IFU.scala 373:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[src/main/scala/nutcore/frontend/IFU.scala 371:36]
  assign io_imem_req_bits_user = {x8_hi,pc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 375:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 393:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/IFU.scala 385:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[src/main/scala/nutcore/frontend/IFU.scala 387:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[src/main/scala/nutcore/frontend/IFU.scala 388:26]
  assign io_out_bits_exceptionVec_1 = io_iaf; // @[src/main/scala/nutcore/frontend/IFU.scala 392:46]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[src/main/scala/nutcore/frontend/IFU.scala 389:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 368:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  assign bp1_io_flush = io_redirect_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
  assign bp1_bpuUpdateReq_valid = REG_valid;
  assign bp1_bpuUpdateReq_pc = REG_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_actualTarget;
  assign bp1_bpuUpdateReq_fuOpType = REG_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_isRVC;
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
      pc <= 39'h80000000; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end else if (pcUpdate) begin // @[src/main/scala/nutcore/frontend/IFU.scala 361:19]
      if (io_redirect_valid) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= snpc;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
      crosslineJumpLatch <= 1'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 331:34]
      if (bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 332:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
      crosslineJumpTarget <= bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_3) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  r = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_0, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_2, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_3, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_4, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_5, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_6, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_7, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_8, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_9, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_10, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_11, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_13, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_14, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_15, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_flush // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
  wire  _instr_T = state == 2'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:23]
  wire  _instr_T_1 = state == 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 44:19]
  reg [15:0] specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
  wire [31:0] _instr_T_4 = {instIn[15:0],specialInstR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:73]
  wire  _pcOffset_T = state == 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:28]
  reg [2:0] pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:21]
  wire  _instr_T_9 = 3'h0 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_13 = _instr_T_9 ? instIn[31:0] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_10 = 3'h2 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_14 = _instr_T_10 ? instIn[47:16] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_17 = _instr_T_13 | _instr_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_11 = 3'h4 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_15 = _instr_T_11 ? instIn[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_18 = _instr_T_17 | _instr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_12 = 3'h6 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_16 = _instr_T_12 ? instIn[79:48] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_19 = _instr_T_18 | _instr_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _instr_T_4 : _instr_T_19; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 34:27]
  wire [7:0] hasException_lo = {io_in_bits_exceptionVec_7,io_in_bits_exceptionVec_6,io_in_bits_exceptionVec_5,
    io_in_bits_exceptionVec_4,io_in_bits_exceptionVec_3,io_in_bits_exceptionVec_2,io_in_bits_exceptionVec_1,
    io_in_bits_exceptionVec_0}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire [15:0] _hasException_T = {io_in_bits_exceptionVec_15,io_in_bits_exceptionVec_14,io_in_bits_exceptionVec_13,
    io_in_bits_exceptionVec_12,io_in_bits_exceptionVec_11,io_in_bits_exceptionVec_10,io_in_bits_exceptionVec_9,
    io_in_bits_exceptionVec_8,hasException_lo}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire  hasException = io_in_valid & |_hasException_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:34]
  wire  _rvcFinish_T = pcOffset == 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:28]
  wire  _rvcFinish_T_1 = ~isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:40]
  wire  _rvcFinish_T_5 = pcOffset == 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:72]
  wire  _rvcFinish_T_11 = pcOffset == 3'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:116]
  wire  _rvcFinish_T_16 = pcOffset == 3'h6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:147]
  wire  _rvcNext_T_13 = _rvcFinish_T_11 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:122]
  wire  _rvcNext_T_15 = ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:135]
  wire  rvcNext = _rvcFinish_T & (isRVC & ~io_in_bits_brIdx[0]) | _rvcFinish_T_5 & (isRVC & ~io_in_bits_brIdx[0]) |
    _rvcFinish_T_11 & _rvcFinish_T_1 & ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:102]
  wire  _rvcSpecial_T_2 = _rvcFinish_T_16 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:37]
  wire  rvcSpecial = _rvcFinish_T_16 & _rvcFinish_T_1 & ~io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:47]
  wire  rvcSpecialJump = _rvcSpecial_T_2 & io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 55:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 56:24]
  wire  _flushIFU_T_2 = _pcOffset_T | state == 2'h1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:36]
  wire  flushIFU = (_pcOffset_T | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:87]
  wire  loadNextInstline = _flushIFU_T_2 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 62:115]
  reg [38:0] specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
  reg [38:0] specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
  reg  specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
  wire  hasCrossBoundaryFault = io_in_bits_exceptionVec_1 | io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 70:73]
  wire  rvcForceLoadNext = _rvcNext_T_13 & io_in_bits_pnpc[2:0] == 3'h4 & _rvcNext_T_15; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 72:86]
  wire  _canGo_T = rvcFinish | rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:28]
  wire  _canIn_T = rvcFinish | rvcForceLoadNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 104:28]
  wire [38:0] _pnpcOut_T_1 = io_in_bits_pc + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:76]
  wire [38:0] _pnpcOut_T_3 = io_in_bits_pc + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:95]
  wire [38:0] _pnpcOut_T_4 = isRVC ? _pnpcOut_T_1 : _pnpcOut_T_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:55]
  wire [38:0] _pnpcOut_T_5 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:23]
  wire  _T_6 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_0 = _T_6 & rvcFinish ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:{39,46} 41:22]
  wire [2:0] _pcOffsetR_T = isRVC ? 3'h2 : 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:38]
  wire [2:0] _pcOffsetR_T_2 = pcOffset + _pcOffsetR_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:33]
  wire [1:0] _GEN_1 = _T_6 & rvcNext ? 2'h1 : _GEN_0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 109:17]
  wire [2:0] _GEN_2 = _T_6 & rvcNext ? _pcOffsetR_T_2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 110:21 42:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 113:17]
  wire [38:0] _pcOut_T_2 = {io_in_bits_pc[38:3],pcOffsetR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 129:21]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 164:15 64:23]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 152:15]
  wire [38:0] _GEN_40 = 2'h1 == state ? _pcOut_T_2 : _GEN_32; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 129:15]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 114:22 66:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 115:24 68:25]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? hasCrossBoundaryFault : specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 116:23 69:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 119:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 120:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 121:23 67:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 122:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? hasCrossBoundaryFault : _GEN_6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 123:23]
  wire [38:0] _pnpcOut_T_7 = pcOut + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:68]
  wire [38:0] _pnpcOut_T_9 = pcOut + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:79]
  wire [38:0] _pnpcOut_T_10 = isRVC ? _pnpcOut_T_7 : _pnpcOut_T_9; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:55]
  wire [38:0] _pnpcOut_T_11 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_10; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:23]
  wire [38:0] _pnpcOut_T_13 = specialPCR + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 153:31]
  wire [1:0] _GEN_24 = _T_6 ? 2'h1 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 158:17 41:22]
  wire [2:0] _GEN_25 = _T_6 ? 3'h2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 159:21 42:26]
  wire [1:0] _GEN_26 = _T_6 ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 169:26 170:17 41:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 165:17 65:25]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 167:15 46:23]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 41:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _pnpcOut_T_13 : _GEN_28; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 153:17]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 155:15]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 156:15]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 42:26]
  wire  _GEN_38 = 2'h1 == state ? _canGo_T : _GEN_34; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 127:15]
  wire  _GEN_39 = 2'h1 == state ? _canIn_T : _GEN_35; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 128:15]
  wire [38:0] _GEN_41 = 2'h1 == state ? _pnpcOut_T_11 : _GEN_33; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 130:17]
  wire [1:0] _GEN_42 = 2'h1 == state ? _GEN_7 : _GEN_36; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire  _GEN_48 = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 103:15]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 104:15]
  wire [38:0] pnpcOut = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  wire  canGo = hasException | _GEN_48; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23 184:11]
  wire  _io_out_bits_brIdx_T_10 = pnpcOut == _pnpcOut_T_9 & _rvcFinish_T_1 | pnpcOut == _pnpcOut_T_7 & isRVC ? 1'h0 : 1'h1
    ; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:27]
  wire  _io_out_bits_exceptionVec_12_T_2 = _instr_T_1 | _instr_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:133]
  assign io_in_ready = ~io_in_valid | _T_6 & canIn | loadNextInstline; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 196:58]
  assign io_out_valid = io_in_valid & canGo; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 195:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 192:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  assign io_out_bits_pnpc = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  assign io_out_bits_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 198:28]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_instr_T_1 | _instr_T); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:87]
  assign io_out_bits_brIdx = {{3'd0}, _io_out_bits_brIdx_T_10}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:21]
  assign io_out_bits_crossBoundaryFault = hasCrossBoundaryFault & _io_out_bits_exceptionVec_12_T_2 & ~specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 200:115]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 183:11]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_42;
      end
    end else begin
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 175:11]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
      pcOffsetR <= 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
      specialIPFR <= 1'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_11;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~flushIFU)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:61 assert(!flushIFU)\n"); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~flushIFU); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
    end
  end
endmodule
module RVCExpander(
  input  [31:0] io_in, // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
  output [31:0] io_out_bits // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
);
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 50:20]
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 51:15]
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 33:18]
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 55:23]
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 32:18]
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 54:22]
  wire [27:0] _io_out_s_T_51 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 53:22]
  wire [26:0] _io_out_s_T_73 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f}; // @[src/main/scala/nutcore/frontend/RVC.scala 60:25]
  wire [27:0] _io_out_s_T_93 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 63:23]
  wire [26:0] _io_out_s_T_115 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 62:22]
  wire [27:0] _io_out_s_T_135 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 61:22]
  wire [6:0] _io_out_s_T_144 = io_in[12] ? 7'h7f : 7'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 40:25]
  wire [11:0] _io_out_s_T_146 = {_io_out_s_T_144,io_in[6:2]}; // @[src/main/scala/nutcore/frontend/RVC.scala 40:20]
  wire [31:0] io_out_s_res_8_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 72:24]
  wire  _io_out_s_opc_T_3 = |io_in[11:7]; // @[src/main/scala/nutcore/frontend/RVC.scala 74:24]
  wire [6:0] io_out_s_opc_1 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 74:20]
  wire [31:0] io_out_s_res_9_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],io_out_s_opc_1}; // @[src/main/scala/nutcore/frontend/RVC.scala 75:15]
  wire [31:0] io_out_s_res_10_bits = {_io_out_s_T_144,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 81:22]
  wire  _io_out_s_opc_T_8 = |_io_out_s_T_146; // @[src/main/scala/nutcore/frontend/RVC.scala 87:29]
  wire [6:0] io_out_s_opc_2 = |_io_out_s_T_146 ? 7'h37 : 7'h3f; // @[src/main/scala/nutcore/frontend/RVC.scala 87:20]
  wire [14:0] _io_out_s_me_T_1 = io_in[12] ? 15'h7fff : 15'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 38:24]
  wire [31:0] _io_out_s_me_T_3 = {_io_out_s_me_T_1,io_in[6:2],12'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 38:19]
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_3[31:12],io_in[11:7],io_out_s_opc_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 88:24]
  wire [6:0] io_out_s_opc_3 = _io_out_s_opc_T_8 ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 83:20]
  wire [2:0] _io_out_s_T_183 = io_in[12] ? 3'h7 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 39:29]
  wire [31:0] io_out_s_res_11_bits = {_io_out_s_T_183,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[
    11:7],io_out_s_opc_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 84:15]
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_11_bits : io_out_s_me_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 89:10]
  wire [25:0] _io_out_s_T_205 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 95:21]
  wire [30:0] _GEN_44 = {{5'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [30:0] _io_out_s_T_214 = _GEN_44 | 31'h40000000; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [31:0] _io_out_s_T_223 = {_io_out_s_T_144,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 97:21]
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]}; // @[src/main/scala/nutcore/frontend/RVC.scala 99:77]
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 100:22]
  wire [6:0] io_out_s_opc_4 = io_in[12] ? 7'h3b : 7'h33; // @[src/main/scala/nutcore/frontend/RVC.scala 101:22]
  wire [2:0] _GEN_1 = 3'h1 == _io_out_s_funct_T_2 ? 3'h4 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_2 = 3'h2 == _io_out_s_funct_T_2 ? 3'h6 : _GEN_1; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_3 = 3'h3 == _io_out_s_funct_T_2 ? 3'h7 : _GEN_2; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_4 = 3'h4 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_3; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_5 = 3'h5 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_4; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_6 = 3'h6 == _io_out_s_funct_T_2 ? 3'h2 : _GEN_5; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_7 = 3'h7 == _io_out_s_funct_T_2 ? 3'h3 : _GEN_6; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [24:0] _io_out_s_T_230 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_GEN_7,2'h1,io_in[9:7],io_out_s_opc_4}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:12]
  wire [30:0] _GEN_45 = {{6'd0}, _io_out_s_T_230}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire [30:0] _io_out_s_T_231 = _GEN_45 | io_out_s_sub; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire [31:0] _io_out_s_WIRE_0 = {{6'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] _io_out_s_WIRE_1 = {{1'd0}, _io_out_s_T_214}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] _GEN_9 = 2'h1 == io_in[11:10] ? _io_out_s_WIRE_1 : _io_out_s_WIRE_0; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [31:0] _GEN_10 = 2'h2 == io_in[11:10] ? _io_out_s_T_223 : _GEN_9; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [31:0] _io_out_s_WIRE_3 = {{1'd0}, _io_out_s_T_231}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] io_out_s_res_12_bits = 2'h3 == io_in[11:10] ? _io_out_s_WIRE_3 : _GEN_10; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [9:0] _io_out_s_T_241 = io_in[12] ? 10'h3ff : 10'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 41:22]
  wire [20:0] _io_out_s_T_249 = {_io_out_s_T_241,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    }; // @[src/main/scala/nutcore/frontend/RVC.scala 41:17]
  wire [31:0] io_out_s_res_13_bits = {_io_out_s_T_249[20],_io_out_s_T_249[10:1],_io_out_s_T_249[11],_io_out_s_T_249[19:
    12],5'h0,7'h6f}; // @[src/main/scala/nutcore/frontend/RVC.scala 91:21]
  wire [4:0] _io_out_s_T_291 = io_in[12] ? 5'h1f : 5'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 42:22]
  wire [12:0] _io_out_s_T_296 = {_io_out_s_T_291,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 42:17]
  wire [31:0] io_out_s_res_14_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h0,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 92:24]
  wire [31:0] io_out_s_res_15_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h1,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 93:24]
  wire [6:0] io_out_s_load_opc = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 110:23]
  wire [25:0] _io_out_s_T_373 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 111:24]
  wire [28:0] _io_out_s_T_383 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 114:25]
  wire [27:0] _io_out_s_T_392 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 113:24]
  wire [28:0] _io_out_s_T_401 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 112:24]
  wire [19:0] _io_out_s_mv_T_2 = {io_in[6:2],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 127:24]
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[src/main/scala/nutcore/frontend/RVC.scala 128:25]
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[src/main/scala/nutcore/frontend/RVC.scala 129:19]
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f}; // @[src/main/scala/nutcore/frontend/RVC.scala 130:25]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[src/main/scala/nutcore/frontend/RVC.scala 131:33]
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2]; // @[src/main/scala/nutcore/frontend/RVC.scala 132:27]
  wire [31:0] io_out_s_mv_bits = {{12'd0}, _io_out_s_mv_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 132:22]
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[src/main/scala/nutcore/frontend/RVC.scala 133:21]
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73}; // @[src/main/scala/nutcore/frontend/RVC.scala 134:23]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000; // @[src/main/scala/nutcore/frontend/RVC.scala 134:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[src/main/scala/nutcore/frontend/RVC.scala 135:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 136:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 137:10]
  wire [8:0] _io_out_s_T_409 = {io_in[9:7],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 37:20]
  wire [28:0] _io_out_s_T_416 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 121:25]
  wire [7:0] _io_out_s_T_422 = {io_in[8:7],io_in[12:9],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 36:20]
  wire [27:0] _io_out_s_T_429 = {_io_out_s_T_422[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_422[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 120:24]
  wire [28:0] _io_out_s_T_442 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 119:24]
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]}; // @[src/main/scala/nutcore/frontend/RVC.scala 148:10]
  wire [31:0] io_out_s_res_bits = {{2'd0}, _io_out_s_T_7}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_res_1_bits = {{4'd0}, _io_out_s_T_20}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_13 = 5'h1 == _io_out_T_2 ? io_out_s_res_1_bits : io_out_s_res_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_2_bits = {{5'd0}, _io_out_s_T_36}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_14 = 5'h2 == _io_out_T_2 ? io_out_s_res_2_bits : _GEN_13; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_3_bits = {{4'd0}, _io_out_s_T_51}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_15 = 5'h3 == _io_out_T_2 ? io_out_s_res_3_bits : _GEN_14; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_4_bits = {{5'd0}, _io_out_s_T_73}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_16 = 5'h4 == _io_out_T_2 ? io_out_s_res_4_bits : _GEN_15; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_5_bits = {{4'd0}, _io_out_s_T_93}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_17 = 5'h5 == _io_out_T_2 ? io_out_s_res_5_bits : _GEN_16; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_6_bits = {{5'd0}, _io_out_s_T_115}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_18 = 5'h6 == _io_out_T_2 ? io_out_s_res_6_bits : _GEN_17; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_7_bits = {{4'd0}, _io_out_s_T_135}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_19 = 5'h7 == _io_out_T_2 ? io_out_s_res_7_bits : _GEN_18; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_20 = 5'h8 == _io_out_T_2 ? io_out_s_res_8_bits : _GEN_19; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_21 = 5'h9 == _io_out_T_2 ? io_out_s_res_9_bits : _GEN_20; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_22 = 5'ha == _io_out_T_2 ? io_out_s_res_10_bits : _GEN_21; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_23 = 5'hb == _io_out_T_2 ? io_out_s_11_bits : _GEN_22; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_24 = 5'hc == _io_out_T_2 ? io_out_s_res_12_bits : _GEN_23; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_25 = 5'hd == _io_out_T_2 ? io_out_s_res_13_bits : _GEN_24; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_26 = 5'he == _io_out_T_2 ? io_out_s_res_14_bits : _GEN_25; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_27 = 5'hf == _io_out_T_2 ? io_out_s_res_15_bits : _GEN_26; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_16_bits = {{6'd0}, _io_out_s_T_373}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_28 = 5'h10 == _io_out_T_2 ? io_out_s_res_16_bits : _GEN_27; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_17_bits = {{3'd0}, _io_out_s_T_383}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_29 = 5'h11 == _io_out_T_2 ? io_out_s_res_17_bits : _GEN_28; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_18_bits = {{4'd0}, _io_out_s_T_392}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_30 = 5'h12 == _io_out_T_2 ? io_out_s_res_18_bits : _GEN_29; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_19_bits = {{3'd0}, _io_out_s_T_401}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_31 = 5'h13 == _io_out_T_2 ? io_out_s_res_19_bits : _GEN_30; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_32 = 5'h14 == _io_out_T_2 ? io_out_s_20_bits : _GEN_31; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_20_bits = {{3'd0}, _io_out_s_T_416}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_33 = 5'h15 == _io_out_T_2 ? io_out_s_res_20_bits : _GEN_32; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_21_bits = {{4'd0}, _io_out_s_T_429}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_34 = 5'h16 == _io_out_T_2 ? io_out_s_res_21_bits : _GEN_33; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_22_bits = {{3'd0}, _io_out_s_T_442}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_35 = 5'h17 == _io_out_T_2 ? io_out_s_res_22_bits : _GEN_34; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_36 = 5'h18 == _io_out_T_2 ? io_in : _GEN_35; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_37 = 5'h19 == _io_out_T_2 ? io_in : _GEN_36; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_38 = 5'h1a == _io_out_T_2 ? io_in : _GEN_37; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_39 = 5'h1b == _io_out_T_2 ? io_in : _GEN_38; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_40 = 5'h1c == _io_out_T_2 ? io_in : _GEN_39; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_41 = 5'h1d == _io_out_T_2 ? io_in : _GEN_40; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_42 = 5'h1e == _io_out_T_2 ? io_in : _GEN_41; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  assign io_out_bits = 5'h1f == _io_out_T_2 ? io_in : _GEN_42; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
endmodule
module Decoder(
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_isWFI, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [11:0] intrVecIDU
);
  wire [31:0] expander_io_in; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] expander_io_out_bits; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] _decodeList_T = expander_io_out_bits & 32'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_1 = 32'h13 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_2 = expander_io_out_bits & 32'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_3 = 32'h1013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_5 = 32'h2013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_7 = 32'h3013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_9 = 32'h4013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_11 = 32'h5013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_13 = 32'h6013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_15 = 32'h7013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_17 = 32'h40005013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_18 = expander_io_out_bits & 32'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_19 = 32'h33 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_21 = 32'h1033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_23 = 32'h2033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_25 = 32'h3033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_27 = 32'h4033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_29 = 32'h5033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_31 = 32'h6033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_33 = 32'h7033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_35 = 32'h40000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_37 = 32'h40005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_38 = expander_io_out_bits & 32'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_39 = 32'h17 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_41 = 32'h37 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_43 = 32'h6f == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_45 = 32'h67 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_47 = 32'h63 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_49 = 32'h1063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_51 = 32'h4063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_53 = 32'h5063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_55 = 32'h6063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_57 = 32'h7063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_59 = 32'h3 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_61 = 32'h1003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_63 = 32'h2003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_65 = 32'h4003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_67 = 32'h5003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_69 = 32'h23 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_71 = 32'h1023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_73 = 32'h2023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_75 = 32'h1b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_77 = 32'h101b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_79 = 32'h501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_81 = 32'h4000501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_83 = 32'h103b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_85 = 32'h503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_87 = 32'h4000503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_89 = 32'h3b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_91 = 32'h4000003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_93 = 32'h6003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_95 = 32'h3003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_97 = 32'h3023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_99 = 32'h6b == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_101 = 32'h2000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_103 = 32'h2001033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_105 = 32'h2002033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_107 = 32'h2003033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_109 = 32'h2004033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_111 = 32'h2005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_113 = 32'h2006033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_115 = 32'h2007033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_117 = 32'h200003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_119 = 32'h200403b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_121 = 32'h200503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_123 = 32'h200603b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_125 = 32'h200703b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_126 = expander_io_out_bits; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_127 = 32'h73 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_129 = 32'h100073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_131 = 32'h30200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_133 = 32'hf == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_135 = 32'h10500073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_137 = 32'h10200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_138 = expander_io_out_bits & 32'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_139 = 32'h12000073 == _decodeList_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_140 = expander_io_out_bits & 32'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_141 = 32'h1000302f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_143 = 32'h1000202f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_144 = expander_io_out_bits & 32'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_145 = 32'h1800302f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_147 = 32'h1800202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_148 = expander_io_out_bits & 32'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_149 = 32'h800202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_151 = 32'h202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_153 = 32'h2000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_155 = 32'h6000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_157 = 32'h4000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_159 = 32'h8000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_161 = 32'ha000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_163 = 32'hc000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_165 = 32'he000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_167 = 32'h1073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_169 = 32'h2073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_171 = 32'h3073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_173 = 32'h5073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_175 = 32'h6073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_177 = 32'h7073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_179 = 32'h100f == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _decodeList_T_181 = _decodeList_T_177 ? 3'h4 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_182 = _decodeList_T_175 ? 3'h4 : _decodeList_T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_183 = _decodeList_T_173 ? 3'h4 : _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_184 = _decodeList_T_171 ? 3'h4 : _decodeList_T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_185 = _decodeList_T_169 ? 3'h4 : _decodeList_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_186 = _decodeList_T_167 ? 3'h4 : _decodeList_T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_187 = _decodeList_T_165 ? 3'h5 : _decodeList_T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_188 = _decodeList_T_163 ? 3'h5 : _decodeList_T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_189 = _decodeList_T_161 ? 3'h5 : _decodeList_T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_190 = _decodeList_T_159 ? 3'h5 : _decodeList_T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_191 = _decodeList_T_157 ? 3'h5 : _decodeList_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_192 = _decodeList_T_155 ? 3'h5 : _decodeList_T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_193 = _decodeList_T_153 ? 3'h5 : _decodeList_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_194 = _decodeList_T_151 ? 3'h5 : _decodeList_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_195 = _decodeList_T_149 ? 3'h5 : _decodeList_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_196 = _decodeList_T_147 ? 4'hf : {{1'd0}, _decodeList_T_195}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_197 = _decodeList_T_145 ? 4'hf : _decodeList_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_198 = _decodeList_T_143 ? 4'h5 : _decodeList_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_199 = _decodeList_T_141 ? 4'h5 : _decodeList_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_200 = _decodeList_T_139 ? 4'h5 : _decodeList_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_201 = _decodeList_T_137 ? 4'h4 : _decodeList_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_202 = _decodeList_T_135 ? 4'h4 : _decodeList_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_203 = _decodeList_T_133 ? 4'h2 : _decodeList_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_204 = _decodeList_T_131 ? 4'h4 : _decodeList_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_205 = _decodeList_T_129 ? 4'h4 : _decodeList_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_206 = _decodeList_T_127 ? 4'h4 : _decodeList_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_207 = _decodeList_T_125 ? 4'h5 : _decodeList_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_208 = _decodeList_T_123 ? 4'h5 : _decodeList_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_209 = _decodeList_T_121 ? 4'h5 : _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_210 = _decodeList_T_119 ? 4'h5 : _decodeList_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_211 = _decodeList_T_117 ? 4'h5 : _decodeList_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_212 = _decodeList_T_115 ? 4'h5 : _decodeList_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_213 = _decodeList_T_113 ? 4'h5 : _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_214 = _decodeList_T_111 ? 4'h5 : _decodeList_T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_215 = _decodeList_T_109 ? 4'h5 : _decodeList_T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_216 = _decodeList_T_107 ? 4'h5 : _decodeList_T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_217 = _decodeList_T_105 ? 4'h5 : _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_218 = _decodeList_T_103 ? 4'h5 : _decodeList_T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_219 = _decodeList_T_101 ? 4'h5 : _decodeList_T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_220 = _decodeList_T_99 ? 4'h4 : _decodeList_T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_221 = _decodeList_T_97 ? 4'h2 : _decodeList_T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_222 = _decodeList_T_95 ? 4'h4 : _decodeList_T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_223 = _decodeList_T_93 ? 4'h4 : _decodeList_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_224 = _decodeList_T_91 ? 4'h5 : _decodeList_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_225 = _decodeList_T_89 ? 4'h5 : _decodeList_T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_226 = _decodeList_T_87 ? 4'h5 : _decodeList_T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_227 = _decodeList_T_85 ? 4'h5 : _decodeList_T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_228 = _decodeList_T_83 ? 4'h5 : _decodeList_T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_229 = _decodeList_T_81 ? 4'h4 : _decodeList_T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_230 = _decodeList_T_79 ? 4'h4 : _decodeList_T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_231 = _decodeList_T_77 ? 4'h4 : _decodeList_T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_232 = _decodeList_T_75 ? 4'h4 : _decodeList_T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_233 = _decodeList_T_73 ? 4'h2 : _decodeList_T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_234 = _decodeList_T_71 ? 4'h2 : _decodeList_T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_235 = _decodeList_T_69 ? 4'h2 : _decodeList_T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_236 = _decodeList_T_67 ? 4'h4 : _decodeList_T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_237 = _decodeList_T_65 ? 4'h4 : _decodeList_T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_238 = _decodeList_T_63 ? 4'h4 : _decodeList_T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_239 = _decodeList_T_61 ? 4'h4 : _decodeList_T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_240 = _decodeList_T_59 ? 4'h4 : _decodeList_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_241 = _decodeList_T_57 ? 4'h1 : _decodeList_T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_242 = _decodeList_T_55 ? 4'h1 : _decodeList_T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_243 = _decodeList_T_53 ? 4'h1 : _decodeList_T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_244 = _decodeList_T_51 ? 4'h1 : _decodeList_T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_245 = _decodeList_T_49 ? 4'h1 : _decodeList_T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_246 = _decodeList_T_47 ? 4'h1 : _decodeList_T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_247 = _decodeList_T_45 ? 4'h4 : _decodeList_T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_248 = _decodeList_T_43 ? 4'h7 : _decodeList_T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_249 = _decodeList_T_41 ? 4'h6 : _decodeList_T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_250 = _decodeList_T_39 ? 4'h6 : _decodeList_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_251 = _decodeList_T_37 ? 4'h5 : _decodeList_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_252 = _decodeList_T_35 ? 4'h5 : _decodeList_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_253 = _decodeList_T_33 ? 4'h5 : _decodeList_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_254 = _decodeList_T_31 ? 4'h5 : _decodeList_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_255 = _decodeList_T_29 ? 4'h5 : _decodeList_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_256 = _decodeList_T_27 ? 4'h5 : _decodeList_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_257 = _decodeList_T_25 ? 4'h5 : _decodeList_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_258 = _decodeList_T_23 ? 4'h5 : _decodeList_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_259 = _decodeList_T_21 ? 4'h5 : _decodeList_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_260 = _decodeList_T_19 ? 4'h5 : _decodeList_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_261 = _decodeList_T_17 ? 4'h4 : _decodeList_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_262 = _decodeList_T_15 ? 4'h4 : _decodeList_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_263 = _decodeList_T_13 ? 4'h4 : _decodeList_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_264 = _decodeList_T_11 ? 4'h4 : _decodeList_T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_265 = _decodeList_T_9 ? 4'h4 : _decodeList_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_266 = _decodeList_T_7 ? 4'h4 : _decodeList_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_267 = _decodeList_T_5 ? 4'h4 : _decodeList_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_268 = _decodeList_T_3 ? 4'h4 : _decodeList_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] decodeList_0 = _decodeList_T_1 ? 4'h4 : _decodeList_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_269 = _decodeList_T_179 ? 3'h4 : 3'h3; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_270 = _decodeList_T_177 ? 3'h3 : _decodeList_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_271 = _decodeList_T_175 ? 3'h3 : _decodeList_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_272 = _decodeList_T_173 ? 3'h3 : _decodeList_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_273 = _decodeList_T_171 ? 3'h3 : _decodeList_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_274 = _decodeList_T_169 ? 3'h3 : _decodeList_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_275 = _decodeList_T_167 ? 3'h3 : _decodeList_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_276 = _decodeList_T_165 ? 3'h1 : _decodeList_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_277 = _decodeList_T_163 ? 3'h1 : _decodeList_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_278 = _decodeList_T_161 ? 3'h1 : _decodeList_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_279 = _decodeList_T_159 ? 3'h1 : _decodeList_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_280 = _decodeList_T_157 ? 3'h1 : _decodeList_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_281 = _decodeList_T_155 ? 3'h1 : _decodeList_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_282 = _decodeList_T_153 ? 3'h1 : _decodeList_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_283 = _decodeList_T_151 ? 3'h1 : _decodeList_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_284 = _decodeList_T_149 ? 3'h1 : _decodeList_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_285 = _decodeList_T_147 ? 3'h1 : _decodeList_T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_286 = _decodeList_T_145 ? 3'h1 : _decodeList_T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_287 = _decodeList_T_143 ? 3'h1 : _decodeList_T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_288 = _decodeList_T_141 ? 3'h1 : _decodeList_T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_289 = _decodeList_T_139 ? 3'h4 : _decodeList_T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_290 = _decodeList_T_137 ? 3'h3 : _decodeList_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_291 = _decodeList_T_135 ? 3'h0 : _decodeList_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_292 = _decodeList_T_133 ? 3'h4 : _decodeList_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_293 = _decodeList_T_131 ? 3'h3 : _decodeList_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_294 = _decodeList_T_129 ? 3'h3 : _decodeList_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_295 = _decodeList_T_127 ? 3'h3 : _decodeList_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_296 = _decodeList_T_125 ? 3'h2 : _decodeList_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_297 = _decodeList_T_123 ? 3'h2 : _decodeList_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_298 = _decodeList_T_121 ? 3'h2 : _decodeList_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_299 = _decodeList_T_119 ? 3'h2 : _decodeList_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_300 = _decodeList_T_117 ? 3'h2 : _decodeList_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_301 = _decodeList_T_115 ? 3'h2 : _decodeList_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_302 = _decodeList_T_113 ? 3'h2 : _decodeList_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_303 = _decodeList_T_111 ? 3'h2 : _decodeList_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_304 = _decodeList_T_109 ? 3'h2 : _decodeList_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_305 = _decodeList_T_107 ? 3'h2 : _decodeList_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_306 = _decodeList_T_105 ? 3'h2 : _decodeList_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_307 = _decodeList_T_103 ? 3'h2 : _decodeList_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_308 = _decodeList_T_101 ? 3'h2 : _decodeList_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_309 = _decodeList_T_99 ? 3'h3 : _decodeList_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_310 = _decodeList_T_97 ? 3'h1 : _decodeList_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_311 = _decodeList_T_95 ? 3'h1 : _decodeList_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_312 = _decodeList_T_93 ? 3'h1 : _decodeList_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_313 = _decodeList_T_91 ? 3'h0 : _decodeList_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_314 = _decodeList_T_89 ? 3'h0 : _decodeList_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_315 = _decodeList_T_87 ? 3'h0 : _decodeList_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_316 = _decodeList_T_85 ? 3'h0 : _decodeList_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_317 = _decodeList_T_83 ? 3'h0 : _decodeList_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_318 = _decodeList_T_81 ? 3'h0 : _decodeList_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_319 = _decodeList_T_79 ? 3'h0 : _decodeList_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_320 = _decodeList_T_77 ? 3'h0 : _decodeList_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_321 = _decodeList_T_75 ? 3'h0 : _decodeList_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_322 = _decodeList_T_73 ? 3'h1 : _decodeList_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_323 = _decodeList_T_71 ? 3'h1 : _decodeList_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_324 = _decodeList_T_69 ? 3'h1 : _decodeList_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_325 = _decodeList_T_67 ? 3'h1 : _decodeList_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_326 = _decodeList_T_65 ? 3'h1 : _decodeList_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_327 = _decodeList_T_63 ? 3'h1 : _decodeList_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_328 = _decodeList_T_61 ? 3'h1 : _decodeList_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_329 = _decodeList_T_59 ? 3'h1 : _decodeList_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_330 = _decodeList_T_57 ? 3'h0 : _decodeList_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_331 = _decodeList_T_55 ? 3'h0 : _decodeList_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_332 = _decodeList_T_53 ? 3'h0 : _decodeList_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_333 = _decodeList_T_51 ? 3'h0 : _decodeList_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_334 = _decodeList_T_49 ? 3'h0 : _decodeList_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_335 = _decodeList_T_47 ? 3'h0 : _decodeList_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_336 = _decodeList_T_45 ? 3'h0 : _decodeList_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_337 = _decodeList_T_43 ? 3'h0 : _decodeList_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_338 = _decodeList_T_41 ? 3'h0 : _decodeList_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_339 = _decodeList_T_39 ? 3'h0 : _decodeList_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_340 = _decodeList_T_37 ? 3'h0 : _decodeList_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_341 = _decodeList_T_35 ? 3'h0 : _decodeList_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_342 = _decodeList_T_33 ? 3'h0 : _decodeList_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_343 = _decodeList_T_31 ? 3'h0 : _decodeList_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_344 = _decodeList_T_29 ? 3'h0 : _decodeList_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_345 = _decodeList_T_27 ? 3'h0 : _decodeList_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_346 = _decodeList_T_25 ? 3'h0 : _decodeList_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_347 = _decodeList_T_23 ? 3'h0 : _decodeList_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_348 = _decodeList_T_21 ? 3'h0 : _decodeList_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_349 = _decodeList_T_19 ? 3'h0 : _decodeList_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_350 = _decodeList_T_17 ? 3'h0 : _decodeList_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_351 = _decodeList_T_15 ? 3'h0 : _decodeList_T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_352 = _decodeList_T_13 ? 3'h0 : _decodeList_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_353 = _decodeList_T_11 ? 3'h0 : _decodeList_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_354 = _decodeList_T_9 ? 3'h0 : _decodeList_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_355 = _decodeList_T_7 ? 3'h0 : _decodeList_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_356 = _decodeList_T_5 ? 3'h0 : _decodeList_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_357 = _decodeList_T_3 ? 3'h0 : _decodeList_T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] decodeList_1 = _decodeList_T_1 ? 3'h0 : _decodeList_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_359 = _decodeList_T_177 ? 3'h7 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_360 = _decodeList_T_175 ? 3'h6 : _decodeList_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_361 = _decodeList_T_173 ? 3'h5 : _decodeList_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_362 = _decodeList_T_171 ? 3'h3 : _decodeList_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_363 = _decodeList_T_169 ? 3'h2 : _decodeList_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_364 = _decodeList_T_167 ? 3'h1 : _decodeList_T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_365 = _decodeList_T_165 ? 6'h32 : {{3'd0}, _decodeList_T_364}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_366 = _decodeList_T_163 ? 6'h31 : _decodeList_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_367 = _decodeList_T_161 ? 6'h30 : _decodeList_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_368 = _decodeList_T_159 ? 6'h37 : _decodeList_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_369 = _decodeList_T_157 ? 6'h26 : _decodeList_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_370 = _decodeList_T_155 ? 6'h25 : _decodeList_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_371 = _decodeList_T_153 ? 6'h24 : _decodeList_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_372 = _decodeList_T_151 ? 7'h63 : {{1'd0}, _decodeList_T_371}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_373 = _decodeList_T_149 ? 7'h22 : _decodeList_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_374 = _decodeList_T_147 ? 7'h21 : _decodeList_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_375 = _decodeList_T_145 ? 7'h21 : _decodeList_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_376 = _decodeList_T_143 ? 7'h20 : _decodeList_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_377 = _decodeList_T_141 ? 7'h20 : _decodeList_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_378 = _decodeList_T_139 ? 7'h2 : _decodeList_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_379 = _decodeList_T_137 ? 7'h0 : _decodeList_T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_380 = _decodeList_T_135 ? 7'h40 : _decodeList_T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_381 = _decodeList_T_133 ? 7'h0 : _decodeList_T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_382 = _decodeList_T_131 ? 7'h0 : _decodeList_T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_383 = _decodeList_T_129 ? 7'h0 : _decodeList_T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_384 = _decodeList_T_127 ? 7'h0 : _decodeList_T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_385 = _decodeList_T_125 ? 7'hf : _decodeList_T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_386 = _decodeList_T_123 ? 7'he : _decodeList_T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_387 = _decodeList_T_121 ? 7'hd : _decodeList_T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_388 = _decodeList_T_119 ? 7'hc : _decodeList_T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_389 = _decodeList_T_117 ? 7'h8 : _decodeList_T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_390 = _decodeList_T_115 ? 7'h7 : _decodeList_T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_391 = _decodeList_T_113 ? 7'h6 : _decodeList_T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_392 = _decodeList_T_111 ? 7'h5 : _decodeList_T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_393 = _decodeList_T_109 ? 7'h4 : _decodeList_T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_394 = _decodeList_T_107 ? 7'h3 : _decodeList_T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_395 = _decodeList_T_105 ? 7'h2 : _decodeList_T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_396 = _decodeList_T_103 ? 7'h1 : _decodeList_T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_397 = _decodeList_T_101 ? 7'h0 : _decodeList_T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_398 = _decodeList_T_99 ? 7'h2 : _decodeList_T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_399 = _decodeList_T_97 ? 7'hb : _decodeList_T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_400 = _decodeList_T_95 ? 7'h3 : _decodeList_T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_401 = _decodeList_T_93 ? 7'h6 : _decodeList_T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_402 = _decodeList_T_91 ? 7'h28 : _decodeList_T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_403 = _decodeList_T_89 ? 7'h60 : _decodeList_T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_404 = _decodeList_T_87 ? 7'h2d : _decodeList_T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_405 = _decodeList_T_85 ? 7'h25 : _decodeList_T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_406 = _decodeList_T_83 ? 7'h21 : _decodeList_T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_407 = _decodeList_T_81 ? 7'h2d : _decodeList_T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_408 = _decodeList_T_79 ? 7'h25 : _decodeList_T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_409 = _decodeList_T_77 ? 7'h21 : _decodeList_T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_410 = _decodeList_T_75 ? 7'h60 : _decodeList_T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_411 = _decodeList_T_73 ? 7'ha : _decodeList_T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_412 = _decodeList_T_71 ? 7'h9 : _decodeList_T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_413 = _decodeList_T_69 ? 7'h8 : _decodeList_T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_414 = _decodeList_T_67 ? 7'h5 : _decodeList_T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_415 = _decodeList_T_65 ? 7'h4 : _decodeList_T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_416 = _decodeList_T_63 ? 7'h2 : _decodeList_T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_417 = _decodeList_T_61 ? 7'h1 : _decodeList_T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_418 = _decodeList_T_59 ? 7'h0 : _decodeList_T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_419 = _decodeList_T_57 ? 7'h17 : _decodeList_T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_420 = _decodeList_T_55 ? 7'h16 : _decodeList_T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_421 = _decodeList_T_53 ? 7'h15 : _decodeList_T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_422 = _decodeList_T_51 ? 7'h14 : _decodeList_T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_423 = _decodeList_T_49 ? 7'h11 : _decodeList_T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_424 = _decodeList_T_47 ? 7'h10 : _decodeList_T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_425 = _decodeList_T_45 ? 7'h5a : _decodeList_T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_426 = _decodeList_T_43 ? 7'h58 : _decodeList_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_427 = _decodeList_T_41 ? 7'h40 : _decodeList_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_428 = _decodeList_T_39 ? 7'h40 : _decodeList_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_429 = _decodeList_T_37 ? 7'hd : _decodeList_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_430 = _decodeList_T_35 ? 7'h8 : _decodeList_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_431 = _decodeList_T_33 ? 7'h7 : _decodeList_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_432 = _decodeList_T_31 ? 7'h6 : _decodeList_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_433 = _decodeList_T_29 ? 7'h5 : _decodeList_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_434 = _decodeList_T_27 ? 7'h4 : _decodeList_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_435 = _decodeList_T_25 ? 7'h3 : _decodeList_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_436 = _decodeList_T_23 ? 7'h2 : _decodeList_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_437 = _decodeList_T_21 ? 7'h1 : _decodeList_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_438 = _decodeList_T_19 ? 7'h40 : _decodeList_T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_439 = _decodeList_T_17 ? 7'hd : _decodeList_T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_440 = _decodeList_T_15 ? 7'h7 : _decodeList_T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_441 = _decodeList_T_13 ? 7'h6 : _decodeList_T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_442 = _decodeList_T_11 ? 7'h5 : _decodeList_T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_443 = _decodeList_T_9 ? 7'h4 : _decodeList_T_442; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_444 = _decodeList_T_7 ? 7'h3 : _decodeList_T_443; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_445 = _decodeList_T_5 ? 7'h2 : _decodeList_T_444; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_446 = _decodeList_T_3 ? 7'h1 : _decodeList_T_445; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] decodeList_2 = _decodeList_T_1 ? 7'h40 : _decodeList_T_446; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  hasIntr = |intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 130:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire  _src1Type_T = 4'h4 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = expander_io_out_bits[19:15]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:28]
  wire [4:0] rt = expander_io_out_bits[24:20]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:43]
  wire [4:0] rd = expander_io_out_bits[11:7]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:58]
  wire  imm_signBit = expander_io_out_bits[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_1 = imm_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_2 = {_imm_T_1,expander_io_out_bits[31:20]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [11:0] _imm_T_5 = {expander_io_out_bits[31:25],rd}; // @[src/main/scala/nutcore/frontend/IDU.scala 82:27]
  wire  imm_signBit_1 = _imm_T_5[11]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_6 = imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_7 = {_imm_T_6,expander_io_out_bits[31:25],rd}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [12:0] _imm_T_17 = {expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 84:27]
  wire  imm_signBit_3 = _imm_T_17[12]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [50:0] _imm_T_18 = imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_19 = {_imm_T_18,expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [31:0] _imm_T_21 = {expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 85:27]
  wire  imm_signBit_4 = _imm_T_21[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _imm_T_22 = imm_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_23 = {_imm_T_22,expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [20:0] _imm_T_28 = {expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 86:27]
  wire  imm_signBit_5 = _imm_T_28[20]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [42:0] _imm_T_29 = imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_30 = {_imm_T_29,expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imm_T_37 = _src1Type_T ? _imm_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_38 = _src1Type_T_2 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_39 = _src1Type_T_3 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_40 = _src1Type_T_4 ? _imm_T_19 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_41 = _src1Type_T_5 ? _imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_42 = _src1Type_T_6 ? _imm_T_30 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_43 = _imm_T_37 | _imm_T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_44 = _imm_T_43 | _imm_T_39; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_45 = _imm_T_44 | _imm_T_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_46 = _imm_T_45 | _imm_T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_9 = rd == 5'h1 | rd == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire [6:0] _GEN_0 = _T_9 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 92:{57,85}]
  wire  _T_15 = rs == 5'h1 | rs == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire [6:0] _GEN_1 = _T_15 ? 7'h5e : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 94:{29,57}]
  wire [6:0] _GEN_2 = _T_9 ? 7'h5c : _GEN_1; // @[src/main/scala/nutcore/frontend/IDU.scala 95:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 93:40]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  is_sfence_vma = fuType == 3'h4 & fuOpType == 7'h2; // @[src/main/scala/nutcore/frontend/IDU.scala 136:45]
  wire  sfence_vma_illegal = is_sfence_vma & io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 137:42]
  wire  wfi_illegal = io_isWFI & io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 138:30]
  wire  illegal_instr = instrType == 4'h0 | sfence_vma_illegal | wfi_illegal; // @[src/main/scala/nutcore/frontend/IDU.scala 139:82]
  RVCExpander expander ( // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
    .io_in(expander_io_in),
    .io_out_bits(expander_io_out_bits)
  );
  assign io_in_ready = ~io_in_valid | _io_in_ready_T_1; // @[src/main/scala/nutcore/frontend/IDU.scala 120:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 119:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 142:49]
  assign io_out_bits_cf_exceptionVec_2 = illegal_instr & ~hasIntr & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 140:74]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 141:47]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_ctrl_src1Type = expander_io_out_bits[6:0] == 7'h37 ? 1'h0 : src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 99:35]
  assign io_out_bits_ctrl_src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 90:32]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rs; // @[src/main/scala/nutcore/frontend/IDU.scala 74:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rt : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 75:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[src/main/scala/nutcore/Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rd : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 77:33]
  assign io_out_bits_ctrl_isNutCoreTrap = _decodeList_T_99 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 144:66]
  assign io_out_bits_data_imm = _imm_T_46 | _imm_T_42; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_isWFI = _decodeList_T_135 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 145:43]
  assign expander_io_in = io_in_bits_instr[31:0]; // @[src/main/scala/nutcore/frontend/IDU.scala 36:18]
endmodule
module IDU(
  output        io_in_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [63:0] io_in_0_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [3:0]  io_in_0_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        isWFI_0,
  input  [11:0] intrVecIDU
);
  wire  decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [2:0] decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [6:0] decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [11:0] decoder_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  isWFI = decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 175:{23,23}]
  Decoder decoder ( // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
    .io_in_ready(decoder_io_in_ready),
    .io_in_valid(decoder_io_in_valid),
    .io_in_bits_instr(decoder_io_in_bits_instr),
    .io_in_bits_pc(decoder_io_in_bits_pc),
    .io_in_bits_pnpc(decoder_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_1(decoder_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_12(decoder_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder_io_in_bits_brIdx),
    .io_in_bits_crossBoundaryFault(decoder_io_in_bits_crossBoundaryFault),
    .io_out_ready(decoder_io_out_ready),
    .io_out_valid(decoder_io_out_valid),
    .io_out_bits_cf_instr(decoder_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(decoder_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(decoder_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(decoder_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(decoder_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(decoder_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(decoder_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(decoder_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_src1Type(decoder_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(decoder_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_imm(decoder_io_out_bits_data_imm),
    .io_isWFI(decoder_io_isWFI),
    .io_sfence_vma_invalid(decoder_io_sfence_vma_invalid),
    .io_wfi_invalid(decoder_io_wfi_invalid),
    .intrVecIDU(decoder_intrVecIDU)
  );
  assign io_in_0_ready = decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign io_out_0_valid = decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_instr = decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pc = decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pnpc = decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_brIdx = decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_crossBoundaryFault = decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src1Type = decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src2Type = decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuType = decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfWen = decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfDest = decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_isNutCoreTrap = decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_data_imm = decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign isWFI_0 = isWFI;
  assign decoder_io_in_valid = io_in_0_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_instr = io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pc = io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_1 = io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_crossBoundaryFault = io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_out_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign decoder_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 171:33]
  assign decoder_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 172:26]
  assign decoder_intrVecIDU = intrVecIDU;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [63:0] io_enq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [3:0]  io_enq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_deq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [63:0] io_deq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_0, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_2, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_3, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_4, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_5, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_6, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_7, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_8, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_9, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_10, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_11, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_12, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_13, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_14, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_15, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [3:0]  io_deq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_flush // @[src/main/scala/utils/FlushableQueue.scala 21:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pnpc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_0 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_1 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_2 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_3 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_4 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_5 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_6 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_7 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_8 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_9 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_10 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_11 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_12 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_13 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_14 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_15 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [3:0] ram_brIdx [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/utils/FlushableQueue.scala 28:41]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 29:33]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 30:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pnpc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pnpc_io_deq_bits_MPORT_data = ram_pnpc[ram_pnpc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign ram_pnpc_MPORT_addr = enq_ptr_value;
  assign ram_pnpc_MPORT_mask = 1'h1;
  assign ram_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_data = ram_exceptionVec_0[ram_exceptionVec_0_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_0_MPORT_data = 1'h0;
  assign ram_exceptionVec_0_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_0_MPORT_mask = 1'h1;
  assign ram_exceptionVec_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_data = ram_exceptionVec_1[ram_exceptionVec_1_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_1_MPORT_data = io_enq_bits_exceptionVec_1;
  assign ram_exceptionVec_1_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_1_MPORT_mask = 1'h1;
  assign ram_exceptionVec_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_data = ram_exceptionVec_2[ram_exceptionVec_2_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_2_MPORT_data = 1'h0;
  assign ram_exceptionVec_2_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_2_MPORT_mask = 1'h1;
  assign ram_exceptionVec_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_data = ram_exceptionVec_3[ram_exceptionVec_3_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_3_MPORT_data = 1'h0;
  assign ram_exceptionVec_3_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_3_MPORT_mask = 1'h1;
  assign ram_exceptionVec_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_data = ram_exceptionVec_4[ram_exceptionVec_4_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_4_MPORT_data = 1'h0;
  assign ram_exceptionVec_4_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_4_MPORT_mask = 1'h1;
  assign ram_exceptionVec_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_data = ram_exceptionVec_5[ram_exceptionVec_5_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_5_MPORT_data = 1'h0;
  assign ram_exceptionVec_5_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_5_MPORT_mask = 1'h1;
  assign ram_exceptionVec_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_data = ram_exceptionVec_6[ram_exceptionVec_6_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_6_MPORT_data = 1'h0;
  assign ram_exceptionVec_6_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_6_MPORT_mask = 1'h1;
  assign ram_exceptionVec_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_data = ram_exceptionVec_7[ram_exceptionVec_7_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_7_MPORT_data = 1'h0;
  assign ram_exceptionVec_7_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_7_MPORT_mask = 1'h1;
  assign ram_exceptionVec_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_data = ram_exceptionVec_8[ram_exceptionVec_8_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_8_MPORT_data = 1'h0;
  assign ram_exceptionVec_8_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_8_MPORT_mask = 1'h1;
  assign ram_exceptionVec_8_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_data = ram_exceptionVec_9[ram_exceptionVec_9_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_9_MPORT_data = 1'h0;
  assign ram_exceptionVec_9_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_9_MPORT_mask = 1'h1;
  assign ram_exceptionVec_9_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_data = ram_exceptionVec_10[ram_exceptionVec_10_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_10_MPORT_data = 1'h0;
  assign ram_exceptionVec_10_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_10_MPORT_mask = 1'h1;
  assign ram_exceptionVec_10_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_data = ram_exceptionVec_11[ram_exceptionVec_11_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_11_MPORT_data = 1'h0;
  assign ram_exceptionVec_11_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_11_MPORT_mask = 1'h1;
  assign ram_exceptionVec_11_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_data = ram_exceptionVec_12[ram_exceptionVec_12_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_12_MPORT_data = 1'h0;
  assign ram_exceptionVec_12_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_12_MPORT_mask = 1'h1;
  assign ram_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_data = ram_exceptionVec_13[ram_exceptionVec_13_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_13_MPORT_data = 1'h0;
  assign ram_exceptionVec_13_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_13_MPORT_mask = 1'h1;
  assign ram_exceptionVec_13_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_data = ram_exceptionVec_14[ram_exceptionVec_14_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_14_MPORT_data = 1'h0;
  assign ram_exceptionVec_14_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_14_MPORT_mask = 1'h1;
  assign ram_exceptionVec_14_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_data = ram_exceptionVec_15[ram_exceptionVec_15_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_15_MPORT_data = 1'h0;
  assign ram_exceptionVec_15_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_15_MPORT_mask = 1'h1;
  assign ram_exceptionVec_15_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx_io_deq_bits_MPORT_en = 1'h1;
  assign ram_brIdx_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_brIdx_io_deq_bits_MPORT_data = ram_brIdx[ram_brIdx_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign ram_brIdx_MPORT_addr = enq_ptr_value;
  assign ram_brIdx_MPORT_mask = 1'h1;
  assign ram_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/utils/FlushableQueue.scala 46:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/utils/FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_0 = ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_1 = ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_2 = ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_3 = ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_4 = ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_5 = ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_6 = ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_7 = ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_8 = ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_9 = ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_10 = ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_11 = ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_13 = ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_14 = ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_15 = ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  always @(posedge clock) begin
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pnpc_MPORT_en & ram_pnpc_MPORT_mask) begin
      ram_pnpc[ram_pnpc_MPORT_addr] <= ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_0_MPORT_en & ram_exceptionVec_0_MPORT_mask) begin
      ram_exceptionVec_0[ram_exceptionVec_0_MPORT_addr] <= ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_1_MPORT_en & ram_exceptionVec_1_MPORT_mask) begin
      ram_exceptionVec_1[ram_exceptionVec_1_MPORT_addr] <= ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_2_MPORT_en & ram_exceptionVec_2_MPORT_mask) begin
      ram_exceptionVec_2[ram_exceptionVec_2_MPORT_addr] <= ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_3_MPORT_en & ram_exceptionVec_3_MPORT_mask) begin
      ram_exceptionVec_3[ram_exceptionVec_3_MPORT_addr] <= ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_4_MPORT_en & ram_exceptionVec_4_MPORT_mask) begin
      ram_exceptionVec_4[ram_exceptionVec_4_MPORT_addr] <= ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_5_MPORT_en & ram_exceptionVec_5_MPORT_mask) begin
      ram_exceptionVec_5[ram_exceptionVec_5_MPORT_addr] <= ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_6_MPORT_en & ram_exceptionVec_6_MPORT_mask) begin
      ram_exceptionVec_6[ram_exceptionVec_6_MPORT_addr] <= ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_7_MPORT_en & ram_exceptionVec_7_MPORT_mask) begin
      ram_exceptionVec_7[ram_exceptionVec_7_MPORT_addr] <= ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_8_MPORT_en & ram_exceptionVec_8_MPORT_mask) begin
      ram_exceptionVec_8[ram_exceptionVec_8_MPORT_addr] <= ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_9_MPORT_en & ram_exceptionVec_9_MPORT_mask) begin
      ram_exceptionVec_9[ram_exceptionVec_9_MPORT_addr] <= ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_10_MPORT_en & ram_exceptionVec_10_MPORT_mask) begin
      ram_exceptionVec_10[ram_exceptionVec_10_MPORT_addr] <= ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_11_MPORT_en & ram_exceptionVec_11_MPORT_mask) begin
      ram_exceptionVec_11[ram_exceptionVec_11_MPORT_addr] <= ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_12_MPORT_en & ram_exceptionVec_12_MPORT_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12_MPORT_addr] <= ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_13_MPORT_en & ram_exceptionVec_13_MPORT_mask) begin
      ram_exceptionVec_13[ram_exceptionVec_13_MPORT_addr] <= ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_14_MPORT_en & ram_exceptionVec_14_MPORT_mask) begin
      ram_exceptionVec_14[ram_exceptionVec_14_MPORT_addr] <= ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_15_MPORT_en & ram_exceptionVec_15_MPORT_mask) begin
      ram_exceptionVec_15[ram_exceptionVec_15_MPORT_addr] <= ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_brIdx_MPORT_en & ram_brIdx_MPORT_mask) begin
      ram_brIdx[ram_brIdx_MPORT_addr] <= ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      enq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 64:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      deq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 65:21]
    end else if (do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 38:17]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/FlushableQueue.scala 26:35]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 67:16]
    end else if (do_enq != do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 41:28]
      maybe_full <= do_enq; // @[src/main/scala/utils/FlushableQueue.scala 42:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_0[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_1[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_2[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_3[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_4[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_5[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_6[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_7[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_8[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_9[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_10[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_11[initvar] = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_13[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_14[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_15[initvar] = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_19[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  enq_ptr_value = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  deq_ptr_value = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  maybe_full = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [86:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [86:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  output        isWFI,
  input         flushICache,
  input         flushTLB,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isMissPredict; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_actualTarget; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [6:0] ifu_REG_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [1:0] ifu_REG_btbType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isRVC; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushICache; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushTLB; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ibf_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_flush; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  idu_io_in_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_isWFI_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [11:0] idu_intrVecIDU; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  ibf_io_in_q_clock; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_reset; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_flush; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  IFU_inorder ifu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ifu_io_out_bits_exceptionVec_1),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_iaf(ifu_io_iaf),
    .REG_valid(ifu_REG_valid),
    .REG_pc(ifu_REG_pc),
    .REG_isMissPredict(ifu_REG_isMissPredict),
    .REG_actualTarget(ifu_REG_actualTarget),
    .REG_fuOpType(ifu_REG_fuOpType),
    .REG_btbType(ifu_REG_btbType),
    .REG_isRVC(ifu_REG_isRVC),
    .flushICache(ifu_flushICache),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_0(ibf_io_in_bits_exceptionVec_0),
    .io_in_bits_exceptionVec_1(ibf_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_2(ibf_io_in_bits_exceptionVec_2),
    .io_in_bits_exceptionVec_3(ibf_io_in_bits_exceptionVec_3),
    .io_in_bits_exceptionVec_4(ibf_io_in_bits_exceptionVec_4),
    .io_in_bits_exceptionVec_5(ibf_io_in_bits_exceptionVec_5),
    .io_in_bits_exceptionVec_6(ibf_io_in_bits_exceptionVec_6),
    .io_in_bits_exceptionVec_7(ibf_io_in_bits_exceptionVec_7),
    .io_in_bits_exceptionVec_8(ibf_io_in_bits_exceptionVec_8),
    .io_in_bits_exceptionVec_9(ibf_io_in_bits_exceptionVec_9),
    .io_in_bits_exceptionVec_10(ibf_io_in_bits_exceptionVec_10),
    .io_in_bits_exceptionVec_11(ibf_io_in_bits_exceptionVec_11),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_exceptionVec_13(ibf_io_in_bits_exceptionVec_13),
    .io_in_bits_exceptionVec_14(ibf_io_in_bits_exceptionVec_14),
    .io_in_bits_exceptionVec_15(ibf_io_in_bits_exceptionVec_15),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ibf_io_out_bits_exceptionVec_1),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossBoundaryFault(ibf_io_out_bits_crossBoundaryFault),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_1(idu_io_in_0_bits_exceptionVec_1),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossBoundaryFault(idu_io_in_0_bits_crossBoundaryFault),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(idu_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(idu_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_sfence_vma_invalid(idu_io_sfence_vma_invalid),
    .io_wfi_invalid(idu_io_wfi_invalid),
    .isWFI_0(idu_isWFI_0),
    .intrVecIDU(idu_intrVecIDU)
  );
  FlushableQueue ibf_io_in_q ( // @[src/main/scala/utils/FlushableQueue.scala 94:21]
    .clock(ibf_io_in_q_clock),
    .reset(ibf_io_in_q_reset),
    .io_enq_ready(ibf_io_in_q_io_enq_ready),
    .io_enq_valid(ibf_io_in_q_io_enq_valid),
    .io_enq_bits_instr(ibf_io_in_q_io_enq_bits_instr),
    .io_enq_bits_pc(ibf_io_in_q_io_enq_bits_pc),
    .io_enq_bits_pnpc(ibf_io_in_q_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_1(ibf_io_in_q_io_enq_bits_exceptionVec_1),
    .io_enq_bits_brIdx(ibf_io_in_q_io_enq_bits_brIdx),
    .io_deq_ready(ibf_io_in_q_io_deq_ready),
    .io_deq_valid(ibf_io_in_q_io_deq_valid),
    .io_deq_bits_instr(ibf_io_in_q_io_deq_bits_instr),
    .io_deq_bits_pc(ibf_io_in_q_io_deq_bits_pc),
    .io_deq_bits_pnpc(ibf_io_in_q_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_0(ibf_io_in_q_io_deq_bits_exceptionVec_0),
    .io_deq_bits_exceptionVec_1(ibf_io_in_q_io_deq_bits_exceptionVec_1),
    .io_deq_bits_exceptionVec_2(ibf_io_in_q_io_deq_bits_exceptionVec_2),
    .io_deq_bits_exceptionVec_3(ibf_io_in_q_io_deq_bits_exceptionVec_3),
    .io_deq_bits_exceptionVec_4(ibf_io_in_q_io_deq_bits_exceptionVec_4),
    .io_deq_bits_exceptionVec_5(ibf_io_in_q_io_deq_bits_exceptionVec_5),
    .io_deq_bits_exceptionVec_6(ibf_io_in_q_io_deq_bits_exceptionVec_6),
    .io_deq_bits_exceptionVec_7(ibf_io_in_q_io_deq_bits_exceptionVec_7),
    .io_deq_bits_exceptionVec_8(ibf_io_in_q_io_deq_bits_exceptionVec_8),
    .io_deq_bits_exceptionVec_9(ibf_io_in_q_io_deq_bits_exceptionVec_9),
    .io_deq_bits_exceptionVec_10(ibf_io_in_q_io_deq_bits_exceptionVec_10),
    .io_deq_bits_exceptionVec_11(ibf_io_in_q_io_deq_bits_exceptionVec_11),
    .io_deq_bits_exceptionVec_12(ibf_io_in_q_io_deq_bits_exceptionVec_12),
    .io_deq_bits_exceptionVec_13(ibf_io_in_q_io_deq_bits_exceptionVec_13),
    .io_deq_bits_exceptionVec_14(ibf_io_in_q_io_deq_bits_exceptionVec_14),
    .io_deq_bits_exceptionVec_15(ibf_io_in_q_io_deq_bits_exceptionVec_15),
    .io_deq_bits_brIdx(ibf_io_in_q_io_deq_bits_brIdx),
    .io_flush(ibf_io_in_q_io_flush)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_crossBoundaryFault = idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_isNutCoreTrap = idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_flushVec = ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:15]
  assign isWFI = idu_isWFI_0;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_out_ready = ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_iaf = io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 122:10]
  assign ifu_REG_valid = REG_valid;
  assign ifu_REG_pc = REG_pc;
  assign ifu_REG_isMissPredict = REG_isMissPredict;
  assign ifu_REG_actualTarget = REG_actualTarget;
  assign ifu_REG_fuOpType = REG_fuOpType;
  assign ifu_REG_btbType = REG_btbType;
  assign ifu_REG_isRVC = REG_isRVC;
  assign ifu_flushICache = flushICache;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = ibf_io_in_q_io_deq_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_instr = ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pc = ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pnpc = ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_0 = ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_1 = ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_2 = ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_3 = ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_4 = ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_5 = ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_6 = ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_7 = ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_8 = ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_9 = ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_10 = ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_11 = ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_12 = ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_13 = ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_14 = ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_15 = ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_brIdx = ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[src/main/scala/nutcore/frontend/Frontend.scala 116:34]
  assign idu_io_in_0_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_1 = idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossBoundaryFault = idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign idu_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 113:29]
  assign idu_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:22]
  assign idu_intrVecIDU = intrVecIDU;
  assign ibf_io_in_q_clock = clock;
  assign ibf_io_in_q_reset = reset;
  assign ibf_io_in_q_io_enq_valid = ifu_io_out_valid; // @[src/main/scala/utils/FlushableQueue.scala 95:22]
  assign ibf_io_in_q_io_enq_bits_instr = ifu_io_out_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pc = ifu_io_out_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_exceptionVec_1 = ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_deq_ready = ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_q_io_flush = ifu_io_flushVec[0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:58]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_instr <= ibf_io_out_bits_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pc <= ibf_io_out_bits_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pnpc <= ibf_io_out_bits_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_1 <= ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_brIdx <= ibf_io_out_bits_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_crossBoundaryFault <= ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  idu_io_in_0_bits_r_crossBoundaryFault = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper(
  input         clock,
  input  [63:0] io_bits_value_1, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_2, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_3, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_4, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_5, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_6, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_7, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_8, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_9, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_10, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_11, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_12, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_13, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_14, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_15, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_16, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_17, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_18, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_19, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_20, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_21, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_22, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_23, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_24, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_25, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_26, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_27, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_28, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_29, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_30, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_31 // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_0; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_1; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_2; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_3; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_4; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_5; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_6; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_7; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_8; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_9; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_10; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_11; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_12; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_13; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_14; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_15; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_16; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_17; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_18; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_19; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_20; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_21; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_22; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_23; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_24; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_25; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_26; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_27; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_28; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_29; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_30; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_31; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchIntRegState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_value_0(dpic_io_value_0),
    .io_value_1(dpic_io_value_1),
    .io_value_2(dpic_io_value_2),
    .io_value_3(dpic_io_value_3),
    .io_value_4(dpic_io_value_4),
    .io_value_5(dpic_io_value_5),
    .io_value_6(dpic_io_value_6),
    .io_value_7(dpic_io_value_7),
    .io_value_8(dpic_io_value_8),
    .io_value_9(dpic_io_value_9),
    .io_value_10(dpic_io_value_10),
    .io_value_11(dpic_io_value_11),
    .io_value_12(dpic_io_value_12),
    .io_value_13(dpic_io_value_13),
    .io_value_14(dpic_io_value_14),
    .io_value_15(dpic_io_value_15),
    .io_value_16(dpic_io_value_16),
    .io_value_17(dpic_io_value_17),
    .io_value_18(dpic_io_value_18),
    .io_value_19(dpic_io_value_19),
    .io_value_20(dpic_io_value_20),
    .io_value_21(dpic_io_value_21),
    .io_value_22(dpic_io_value_22),
    .io_value_23(dpic_io_value_23),
    .io_value_24(dpic_io_value_24),
    .io_value_25(dpic_io_value_25),
    .io_value_26(dpic_io_value_26),
    .io_value_27(dpic_io_value_27),
    .io_value_28(dpic_io_value_28),
    .io_value_29(dpic_io_value_29),
    .io_value_30(dpic_io_value_30),
    .io_value_31(dpic_io_value_31),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_value_0 = 64'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_1 = io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_2 = io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_3 = io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_4 = io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_5 = io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_6 = io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_7 = io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_8 = io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_9 = io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_10 = io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_11 = io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_12 = io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_13 = io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_14 = io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_15 = io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_16 = io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_17 = io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_18 = io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_19 = io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_20 = io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_21 = io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_22 = io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_23 = io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_24 = io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_25 = io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_26 = io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_27 = io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_28 = io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_29 = io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_30 = io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_31 = io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_flush // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  _src1ForwardNextCycle_T = ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _src1ForwardNextCycle_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 51:43]
  wire  _src1Forward_T_1 = dontForward1 ? ~src1DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _src1Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:34]
  wire  _src2Forward_T_1 = dontForward1 ? ~src2DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _src2Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:34]
  reg [31:0] busy; // @[src/main/scala/nutcore/RF.scala 37:21]
  wire [31:0] _src1Ready_T = busy >> io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/RF.scala 38:37]
  wire  src1Ready = ~_src1Ready_T[0] | src1ForwardNextCycle | src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 56:62]
  wire [31:0] _src2Ready_T = busy >> io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/RF.scala 38:37]
  wire  src2Ready = ~_src2Ready_T[0] | src2ForwardNextCycle | src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 57:62]
  reg [63:0] rf_0; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_1; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_2; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_3; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_4; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_5; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_6; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_7; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_8; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_9; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_10; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_11; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_12; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_13; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_14; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_15; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_16; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_17; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_18; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_19; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_20; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_21; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_22; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_23; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_24; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_25; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_26; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_27; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_28; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_29; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_30; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_31; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  io_out_bits_data_src1_signBit = io_in_0_bits_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _io_out_bits_data_src1_T_1 = io_out_bits_data_src1_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_data_src1_T_2 = {_io_out_bits_data_src1_T_1,io_in_0_bits_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _io_out_bits_data_src1_T_3 = ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:21]
  wire  _io_out_bits_data_src1_T_4 = src1Forward & ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:18]
  wire  _io_out_bits_data_src1_T_9 = ~io_in_0_bits_ctrl_src1Type & _io_out_bits_data_src1_T_3 & ~src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 67:76]
  wire [63:0] _GEN_1 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_2 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? rf_2 : _GEN_1; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_3 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? rf_3 : _GEN_2; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_4 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? rf_4 : _GEN_3; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_5 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? rf_5 : _GEN_4; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_6 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? rf_6 : _GEN_5; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_7 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? rf_7 : _GEN_6; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_8 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? rf_8 : _GEN_7; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_9 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? rf_9 : _GEN_8; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_10 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? rf_10 : _GEN_9; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_11 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? rf_11 : _GEN_10; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_12 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? rf_12 : _GEN_11; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_13 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? rf_13 : _GEN_12; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_14 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? rf_14 : _GEN_13; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_15 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? rf_15 : _GEN_14; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_16 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? rf_16 : _GEN_15; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_17 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? rf_17 : _GEN_16; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_18 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? rf_18 : _GEN_17; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_19 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? rf_19 : _GEN_18; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_20 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? rf_20 : _GEN_19; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_21 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? rf_21 : _GEN_20; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_22 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? rf_22 : _GEN_21; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_23 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? rf_23 : _GEN_22; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_24 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? rf_24 : _GEN_23; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_25 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? rf_25 : _GEN_24; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_26 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? rf_26 : _GEN_25; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_27 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? rf_27 : _GEN_26; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_28 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? rf_28 : _GEN_27; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_29 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? rf_29 : _GEN_28; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_30 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? rf_30 : _GEN_29; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_31 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? rf_31 : _GEN_30; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _io_out_bits_data_src1_T_11 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : _GEN_31; // @[src/main/scala/nutcore/RF.scala 32:36]
  wire [63:0] _io_out_bits_data_src1_T_12 = io_in_0_bits_ctrl_src1Type ? _io_out_bits_data_src1_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_13 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_14 = _io_out_bits_data_src1_T_4 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_15 = _io_out_bits_data_src1_T_9 ? _io_out_bits_data_src1_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_16 = _io_out_bits_data_src1_T_12 | _io_out_bits_data_src1_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_17 = _io_out_bits_data_src1_T_16 | _io_out_bits_data_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_bits_data_src2_T_1 = ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:21]
  wire  _io_out_bits_data_src2_T_2 = src2Forward & ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:18]
  wire  _io_out_bits_data_src2_T_7 = ~io_in_0_bits_ctrl_src2Type & _io_out_bits_data_src2_T_1 & ~src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 73:77]
  wire [63:0] _GEN_33 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_34 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? rf_2 : _GEN_33; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_35 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? rf_3 : _GEN_34; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_36 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? rf_4 : _GEN_35; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_37 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? rf_5 : _GEN_36; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_38 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? rf_6 : _GEN_37; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_39 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? rf_7 : _GEN_38; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_40 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? rf_8 : _GEN_39; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_41 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? rf_9 : _GEN_40; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_42 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? rf_10 : _GEN_41; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_43 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? rf_11 : _GEN_42; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_44 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? rf_12 : _GEN_43; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_45 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? rf_13 : _GEN_44; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_46 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? rf_14 : _GEN_45; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_47 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? rf_15 : _GEN_46; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_48 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? rf_16 : _GEN_47; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_49 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? rf_17 : _GEN_48; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_50 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? rf_18 : _GEN_49; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_51 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? rf_19 : _GEN_50; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_52 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? rf_20 : _GEN_51; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_53 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? rf_21 : _GEN_52; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_54 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? rf_22 : _GEN_53; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_55 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? rf_23 : _GEN_54; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_56 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? rf_24 : _GEN_55; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_57 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? rf_25 : _GEN_56; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_58 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? rf_26 : _GEN_57; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_59 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? rf_27 : _GEN_58; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_60 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? rf_28 : _GEN_59; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_61 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? rf_29 : _GEN_60; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_62 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? rf_30 : _GEN_61; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_63 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? rf_31 : _GEN_62; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _io_out_bits_data_src2_T_9 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : _GEN_63; // @[src/main/scala/nutcore/RF.scala 32:36]
  wire [63:0] _io_out_bits_data_src2_T_10 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_11 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_12 = _io_out_bits_data_src2_T_2 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_13 = _io_out_bits_data_src2_T_7 ? _io_out_bits_data_src2_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_14 = _io_out_bits_data_src2_T_10 | _io_out_bits_data_src2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_15 = _io_out_bits_data_src2_T_14 | _io_out_bits_data_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wbClearMask_T_3 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire [62:0] _wbClearMask_T_6 = 63'h1 << io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 39:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_wbClearMask_T_3 ? _wbClearMask_T_6[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 85:24]
  wire  _isuFireSetMask_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [62:0] _isuFireSetMask_T_1 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/RF.scala 39:39]
  wire [31:0] isuFireSetMask = _isuFireSetMask_T ? _isuFireSetMask_T_1[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 87:27]
  wire [31:0] _busy_T_5 = ~wbClearMask; // @[src/main/scala/nutcore/RF.scala 45:26]
  wire [31:0] _busy_T_6 = busy & _busy_T_5; // @[src/main/scala/nutcore/RF.scala 45:24]
  wire [31:0] _busy_T_7 = _busy_T_6 | isuFireSetMask; // @[src/main/scala/nutcore/RF.scala 45:38]
  wire [31:0] _busy_T_9 = {_busy_T_7[31:1],1'h0}; // @[src/main/scala/nutcore/RF.scala 45:16]
  wire  _T_3 = io_in_0_valid & ~io_out_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 97:40]
  wire  _T_6 = io_out_valid & ~_isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 98:38]
  wire  _T_7 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  DummyDPICWrapper difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .io_bits_value_1(difftest_module_io_bits_value_1),
    .io_bits_value_2(difftest_module_io_bits_value_2),
    .io_bits_value_3(difftest_module_io_bits_value_3),
    .io_bits_value_4(difftest_module_io_bits_value_4),
    .io_bits_value_5(difftest_module_io_bits_value_5),
    .io_bits_value_6(difftest_module_io_bits_value_6),
    .io_bits_value_7(difftest_module_io_bits_value_7),
    .io_bits_value_8(difftest_module_io_bits_value_8),
    .io_bits_value_9(difftest_module_io_bits_value_9),
    .io_bits_value_10(difftest_module_io_bits_value_10),
    .io_bits_value_11(difftest_module_io_bits_value_11),
    .io_bits_value_12(difftest_module_io_bits_value_12),
    .io_bits_value_13(difftest_module_io_bits_value_13),
    .io_bits_value_14(difftest_module_io_bits_value_14),
    .io_bits_value_15(difftest_module_io_bits_value_15),
    .io_bits_value_16(difftest_module_io_bits_value_16),
    .io_bits_value_17(difftest_module_io_bits_value_17),
    .io_bits_value_18(difftest_module_io_bits_value_18),
    .io_bits_value_19(difftest_module_io_bits_value_19),
    .io_bits_value_20(difftest_module_io_bits_value_20),
    .io_bits_value_21(difftest_module_io_bits_value_21),
    .io_bits_value_22(difftest_module_io_bits_value_22),
    .io_bits_value_23(difftest_module_io_bits_value_23),
    .io_bits_value_24(difftest_module_io_bits_value_24),
    .io_bits_value_25(difftest_module_io_bits_value_25),
    .io_bits_value_26(difftest_module_io_bits_value_26),
    .io_bits_value_27(difftest_module_io_bits_value_27),
    .io_bits_value_28(difftest_module_io_bits_value_28),
    .io_bits_value_29(difftest_module_io_bits_value_29),
    .io_bits_value_30(difftest_module_io_bits_value_30),
    .io_bits_value_31(difftest_module_io_bits_value_31)
  );
  assign io_in_0_ready = ~io_in_0_valid | _isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[src/main/scala/nutcore/backend/seq/ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_data_src1 = _io_out_bits_data_src1_T_17 | _io_out_bits_data_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_src2 = _io_out_bits_data_src2_T_15 | _io_out_bits_data_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/ISU.scala 75:25]
  assign difftest_module_clock = clock;
  assign difftest_module_io_bits_value_1 = rf_1; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_2 = rf_2; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_3 = rf_3; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_4 = rf_4; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_5 = rf_5; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_6 = rf_6; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_7 = rf_7; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_8 = rf_8; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_9 = rf_9; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_10 = rf_10; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_11 = rf_11; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_12 = rf_12; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_13 = rf_13; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_14 = rf_14; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_15 = rf_15; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_16 = rf_16; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_17 = rf_17; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_18 = rf_18; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_19 = rf_19; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_20 = rf_20; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_21 = rf_21; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_22 = rf_22; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_23 = rf_23; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_24 = rf_24; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_25 = rf_25; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_26 = rf_26; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_27 = rf_27; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_28 = rf_28; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_29 = rf_29; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_30 = rf_30; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_31 = rf_31; // @[src/main/scala/nutcore/RF.scala 32:36]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 37:21]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 37:21]
    end else if (io_flush) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 88:19]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 45:10]
    end else begin
      busy <= _busy_T_9; // @[src/main/scala/nutcore/RF.scala 45:10]
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h0 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_0 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_1 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_1 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_2 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h2 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_2 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_3 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h3 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_3 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_4 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h4 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_4 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_5 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h5 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_5 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_6 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h6 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_6 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_7 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h7 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_7 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_8 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h8 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_8 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_9 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h9 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_9 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_10 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'ha == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_10 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_11 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hb == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_11 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_12 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hc == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_12 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_13 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hd == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_13 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_14 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'he == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_14 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_15 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hf == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_15 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_16 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h10 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_16 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_17 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h11 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_17 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_18 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h12 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_18 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_19 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h13 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_19 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_20 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h14 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_20 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_21 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h15 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_21 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_22 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h16 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_22 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_23 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h17 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_23 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_24 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h18 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_24 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_25 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h19 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_25 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_26 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1a == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_26 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_27 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1b == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_27 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_28 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1c == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_28 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_29 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1d == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_29 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_30 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1e == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_30 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_31 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1f == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_31 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  rf_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  rf_31 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pnpc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [3:0]  io_cfIn_brIdx, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_offset, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_iVmEnable, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_jumpIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_jumpIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_jumpIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 89:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:39]
  wire [63:0] _adderRes_T_1 = io_in_bits_src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:33]
  wire [64:0] _adderRes_T_2 = io_in_bits_src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:24]
  wire [64:0] _GEN_3 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 91:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 92:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/ALU.scala 93:28]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  shsrc1_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _shsrc1_T_4 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _shsrc1_T_5 = {_shsrc1_T_4,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _shsrc1_T_7 = 7'h25 == io_in_bits_func ? _shsrc1_T_2 : io_in_bits_src1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:18]
  wire [126:0] _GEN_6 = {{63'd0}, shsrc1}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [126:0] _res_T_1 = _GEN_6 << shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 105:32]
  wire [63:0] _res_T_6 = io_in_bits_src1 | io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:30]
  wire [63:0] _res_T_7 = io_in_bits_src1 & io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 107:30]
  wire [63:0] _res_T_8 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:32]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:49]
  wire [64:0] _res_T_12 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_1[63:0]} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_3} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_4} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_5} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_7} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  aluRes_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _aluRes_T_2 = aluRes_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _aluRes_T_3 = {_aluRes_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _aluRes_T_3} : res; // @[src/main/scala/nutcore/backend/fu/ALU.scala 110:19]
  wire  _T_1 = ~(|xorRes); // @[src/main/scala/nutcore/backend/fu/ALU.scala 113:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _taken_T_1 = 2'h0 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_2 = 2'h2 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_3 = 2'h3 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_8 = _taken_T_1 & _T_1 | _taken_T_2 & slt | _taken_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  taken = _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
  wire  target_signBit = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _target_T = target_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _target_T_1 = {_target_T,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _target_T_3 = _target_T_1 + io_offset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:56]
  wire [63:0] _target_T_5 = {adderRes[63:1],1'h0}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:72]
  wire [63:0] target = isBranch ? _target_T_3 : _target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
  wire  _predictWrong_T_1 = ~taken & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
  wire [38:0] _io_redirect_target_T_3 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:71]
  wire [38:0] _io_redirect_target_T_5 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:89]
  wire [38:0] _io_redirect_target_T_6 = isRVC ? _io_redirect_target_T_3 : _io_redirect_target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:52]
  wire [63:0] _io_redirect_target_T_7 = _predictWrong_T_1 ? {{25'd0}, _io_redirect_target_T_6} : target; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:28]
  wire  _io_redirect_valid_T = io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:30]
  wire  _io_redirect_valid_T_1 = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  wire  _io_out_bits_T = ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:33]
  wire [63:0] _io_out_bits_T_4 = _target_T_1 + 64'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:71]
  wire [63:0] _io_out_bits_T_8 = _target_T_1 + 64'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:108]
  wire [63:0] _io_out_bits_T_9 = ~isRVC ? _io_out_bits_T_4 : _io_out_bits_T_8; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:32]
  wire [64:0] _io_out_bits_T_10 = isBru ? {{1'd0}, _io_out_bits_T_9} : aluRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:21]
  reg  hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
  wire  addrNotLegal_signBit = target[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,target[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  addrNotLegal = io_iVmEnable ? target != _addrNotLegal_T_2 : |target[63:39]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 139:25]
  wire  isIllegalJumpAddr = io_redirect_valid & ~isBranch & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/ALU.scala 140:58]
  wire  _T_15 = io_jumpIsIllegal_ready & io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_0 = _T_15 ? 1'h0 : hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:38 144:24 138:35]
  wire  _GEN_1 = isIllegalJumpAddr | _GEN_0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 141:28 142:24]
  reg [63:0] io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
  wire  _bpuUpdateReq_btbType_T_6 = 7'h5c == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _bpuUpdateReq_btbType_T_7 = 7'h5e == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _bpuUpdateReq_btbType_T_8 = 7'h58 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _bpuUpdateReq_btbType_T_9 = 7'h5a == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [1:0] _bpuUpdateReq_btbType_T_17 = _bpuUpdateReq_btbType_T_7 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _bpuUpdateReq_btbType_T_19 = _bpuUpdateReq_btbType_T_9 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_4 = {{1'd0}, _bpuUpdateReq_btbType_T_6}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _bpuUpdateReq_btbType_T_26 = _GEN_4 | _bpuUpdateReq_btbType_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_5 = {{1'd0}, _bpuUpdateReq_btbType_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _bpuUpdateReq_btbType_T_27 = _bpuUpdateReq_btbType_T_26 | _GEN_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [6:0] REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [1:0] REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  right = _io_redirect_valid_T & ~predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:32]
  wire  _T_55 = right & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:33]
  wire  _T_56 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 179:33]
  wire  _T_60 = _T_56 & io_cfIn_pc[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:45]
  wire  _T_61 = _T_56 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:73]
  wire  _T_67 = _T_60 & _io_out_bits_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 181:73]
  wire  _T_71 = _T_56 & io_cfIn_pc[2:0] == 3'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:45]
  wire  _T_72 = _T_56 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:73]
  wire  _T_78 = _T_71 & _io_out_bits_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 183:73]
  wire  _T_82 = _T_56 & io_cfIn_pc[2:0] == 3'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:45]
  wire  _T_83 = _T_56 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:73]
  wire  _T_89 = _T_82 & _io_out_bits_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 185:73]
  wire  _T_93 = _T_56 & io_cfIn_pc[2:0] == 3'h6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:45]
  wire  _T_94 = _T_56 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:73]
  wire  _T_100 = _T_93 & _io_out_bits_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 187:73]
  wire  _T_103 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[src/main/scala/nutcore/backend/fu/ALU.scala 188:60]
  wire  _T_104 = right & (io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c); // @[src/main/scala/nutcore/backend/fu/ALU.scala 188:33]
  wire  _T_108 = _io_redirect_valid_T_1 & _T_103; // @[src/main/scala/nutcore/backend/fu/ALU.scala 189:33]
  wire  _T_109 = io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 190:41]
  wire  _T_110 = right & io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 190:33]
  wire  _T_112 = _io_redirect_valid_T_1 & _T_109; // @[src/main/scala/nutcore/backend/fu/ALU.scala 191:33]
  wire  _T_113 = io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 192:41]
  wire  _T_114 = right & io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 192:33]
  wire  _T_116 = _io_redirect_valid_T_1 & _T_113; // @[src/main/scala/nutcore/backend/fu/ALU.scala 193:33]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 161:16]
  assign io_out_bits = _io_out_bits_T_10[63:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:15]
  assign io_redirect_target = _io_redirect_target_T_7[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:22]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  assign io_jumpIsIllegal_valid = hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 146:26]
  assign io_jumpIsIllegal_bits = io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:25]
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
      hasIllegalJumpAddr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
    end else begin
      hasIllegalJumpAddr <= _GEN_1;
    end
    if (isIllegalJumpAddr) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
      if (isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
        io_jumpIsIllegal_bits_r <= _target_T_3;
      end else begin
        io_jumpIsIllegal_bits_r <= _target_T_5;
      end
    end
    REG_valid <= io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 164:31]
    REG_pc <= io_cfIn_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 165:19]
    if (~taken & isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= target[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 167:29]
    REG_actualTaken <= _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
    REG_fuOpType <= io_in_bits_func; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 169:25]
    REG_btbType <= _bpuUpdateReq_btbType_T_27 | _bpuUpdateReq_btbType_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:124 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasIllegalJumpAddr = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  io_jumpIsIllegal_bits_r = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  REG_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  REG_pc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  REG_actualTarget = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  REG_actualTaken = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_fuOpType = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  REG_btbType = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  REG_isRVC = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
    end
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_resp_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         DTLBPF,
  input         scIsSuccess_0,
  input         vmEnable_0,
  input         ISAMO2,
  input         DTLBFINISH,
  input         DTLBAF
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  _io_vaddr_T = io__in_ready & io__in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 423:23]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 424:30]
  reg [1:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
  wire [5:0] vaddrPF_lo_lo = {io__vaddr[58] != io__vaddr[38],io__vaddr[59] != io__vaddr[38],io__vaddr[60] != io__vaddr[
    38],io__vaddr[61] != io__vaddr[38],io__vaddr[62] != io__vaddr[38],io__vaddr[63] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [11:0] vaddrPF_lo = {io__vaddr[52] != io__vaddr[38],io__vaddr[53] != io__vaddr[38],io__vaddr[54] != io__vaddr[38]
    ,io__vaddr[55] != io__vaddr[38],io__vaddr[56] != io__vaddr[38],io__vaddr[57] != io__vaddr[38],vaddrPF_lo_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [5:0] vaddrPF_hi_lo = {io__vaddr[46] != io__vaddr[38],io__vaddr[47] != io__vaddr[38],io__vaddr[48] != io__vaddr[
    38],io__vaddr[49] != io__vaddr[38],io__vaddr[50] != io__vaddr[38],io__vaddr[51] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [24:0] _vaddrPF_T_76 = {io__vaddr[39] != io__vaddr[38],io__vaddr[40] != io__vaddr[38],io__vaddr[41] != io__vaddr[
    38],io__vaddr[42] != io__vaddr[38],io__vaddr[43] != io__vaddr[38],io__vaddr[44] != io__vaddr[38],io__vaddr[45] !=
    io__vaddr[38],vaddrPF_hi_lo,vaddrPF_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire  vaddrPF = io__in_valid & vmEnable_0 & |_vaddrPF_T_76; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:37]
  wire  dtlbHasException = DTLBPF | DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 446:33]
  wire  _T_1 = io__dmem_req_ready & io__dmem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_4 = ~vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:32]
  wire [1:0] _GEN_3 = DTLBFINISH & (dtlbHasException | ~scIsSuccess_0) ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 454:{63,71}]
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _state_T = partialLoad ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 457:62]
  wire [1:0] _GEN_5 = _T_14 ? _state_T : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 457:{48,56}]
  wire [1:0] _GEN_6 = 2'h3 == state ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18 427:22 458:32]
  wire [1:0] size = io__in_bits_func[1:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 465:18]
  wire [63:0] _reqWdata_T_3 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]
    ,io__wdata[7:0],io__wdata[7:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 399:22]
  wire [63:0] _reqWdata_T_6 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 400:22]
  wire [63:0] _reqWdata_T_8 = {io__wdata[31:0],io__wdata[31:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 401:22]
  wire  _reqWdata_T_9 = 2'h0 == size; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_10 = 2'h1 == size; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_11 = 2'h2 == size; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_12 = 2'h3 == size; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _reqWdata_T_13 = _reqWdata_T_9 ? _reqWdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_14 = _reqWdata_T_10 ? _reqWdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_15 = _reqWdata_T_11 ? _reqWdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_16 = _reqWdata_T_12 ? io__wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_17 = _reqWdata_T_13 | _reqWdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_18 = _reqWdata_T_17 | _reqWdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_5 = _reqWdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_6 = _reqWdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_7 = _reqWdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_14 = {{1'd0}, _reqWdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_8 = _GEN_14 | _reqWmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_15 = {{2'd0}, _reqWmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_9 = _GEN_15 | _reqWmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_16 = {{4'd0}, _reqWmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_10 = _GEN_16 | _reqWmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_24 = {{7'd0}, _reqWmask_T_10}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire [14:0] reqWmask = _GEN_24 << io__in_bits_src1[2:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire  hasException = io__loadAccessFault | io__storeAccessFault | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 476:64]
  wire  _io_dmem_req_valid_T = state == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:37]
  wire  _io_out_valid_T_3 = state == 2'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 483:13]
  wire  _io_out_valid_T_6 = _T_14 & state == 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 484:22]
  wire  _io_out_valid_T_7 = partialLoad ? _io_out_valid_T_3 : _io_out_valid_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 482:8]
  reg [63:0] rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
  wire  _rdataSel64_T_9 = 3'h0 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_10 = 3'h1 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_11 = 3'h2 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_12 = 3'h3 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_13 = 3'h4 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_14 = 3'h5 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_15 = 3'h6 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_16 = 3'h7 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataSel64_T_17 = _rdataSel64_T_9 ? rdataLatch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdataSel64_T_18 = _rdataSel64_T_10 ? rdataLatch[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdataSel64_T_19 = _rdataSel64_T_11 ? rdataLatch[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdataSel64_T_20 = _rdataSel64_T_12 ? rdataLatch[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdataSel64_T_21 = _rdataSel64_T_13 ? rdataLatch[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdataSel64_T_22 = _rdataSel64_T_14 ? rdataLatch[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdataSel64_T_23 = _rdataSel64_T_15 ? rdataLatch[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdataSel64_T_24 = _rdataSel64_T_16 ? rdataLatch[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_17 = {{8'd0}, _rdataSel64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_25 = _rdataSel64_T_17 | _GEN_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_18 = {{16'd0}, _rdataSel64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_26 = _rdataSel64_T_25 | _GEN_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_19 = {{24'd0}, _rdataSel64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_27 = _rdataSel64_T_26 | _GEN_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_20 = {{32'd0}, _rdataSel64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_28 = _rdataSel64_T_27 | _GEN_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_21 = {{40'd0}, _rdataSel64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_29 = _rdataSel64_T_28 | _GEN_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_22 = {{48'd0}, _rdataSel64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_30 = _rdataSel64_T_29 | _GEN_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_23 = {{56'd0}, _rdataSel64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataSel64 = _rdataSel64_T_30 | _GEN_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdataPartialLoad_signBit = rdataSel64[7]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [55:0] _rdataPartialLoad_T_1 = rdataPartialLoad_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_2 = {_rdataPartialLoad_T_1,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_1 = rdataSel64[15]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [47:0] _rdataPartialLoad_T_4 = rdataPartialLoad_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_5 = {_rdataPartialLoad_T_4,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_2 = rdataSel64[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _rdataPartialLoad_T_7 = rdataPartialLoad_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_8 = {_rdataPartialLoad_T_7,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _rdataPartialLoad_T_10 = {56'h0,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_12 = {48'h0,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_14 = {32'h0,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdataPartialLoad_T_15 = 7'h0 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_16 = 7'h1 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_17 = 7'h2 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_18 = 7'h4 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_19 = 7'h5 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_20 = 7'h6 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataPartialLoad_T_21 = _rdataPartialLoad_T_15 ? _rdataPartialLoad_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_22 = _rdataPartialLoad_T_16 ? _rdataPartialLoad_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_23 = _rdataPartialLoad_T_17 ? _rdataPartialLoad_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_24 = _rdataPartialLoad_T_18 ? _rdataPartialLoad_T_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_25 = _rdataPartialLoad_T_19 ? _rdataPartialLoad_T_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_26 = _rdataPartialLoad_T_20 ? _rdataPartialLoad_T_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_27 = _rdataPartialLoad_T_21 | _rdataPartialLoad_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_28 = _rdataPartialLoad_T_27 | _rdataPartialLoad_T_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_29 = _rdataPartialLoad_T_28 | _rdataPartialLoad_T_24; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_30 = _rdataPartialLoad_T_29 | _rdataPartialLoad_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataPartialLoad = _rdataPartialLoad_T_30 | _rdataPartialLoad_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_loadAccessFault_T_1 = io__in_valid & _T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:32]
  wire  _io_loadAccessFault_T_7 = io__in_bits_src1 >= 64'h38000000 & io__in_bits_src1 < 64'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_10 = io__in_bits_src1 >= 64'h3c000000 & io__in_bits_src1 < 64'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_13 = io__in_bits_src1 >= 64'h40600000 & io__in_bits_src1 < 64'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_16 = io__in_bits_src1 >= 64'h50000000 & io__in_bits_src1 < 64'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_19 = io__in_bits_src1 >= 64'h40001000 & io__in_bits_src1 < 64'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_22 = io__in_bits_src1 >= 64'h40000000 & io__in_bits_src1 < 64'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_25 = io__in_bits_src1 >= 64'h40002000 & io__in_bits_src1 < 64'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_28 = io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _io_loadAccessFault_T_29 = {_io_loadAccessFault_T_28,_io_loadAccessFault_T_25,_io_loadAccessFault_T_22,
    _io_loadAccessFault_T_19,_io_loadAccessFault_T_16,_io_loadAccessFault_T_13,_io_loadAccessFault_T_10,
    _io_loadAccessFault_T_7}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _io_loadAccessFault_T_30 = |_io_loadAccessFault_T_29; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _io_loadAccessFault_T_31 = ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:71]
  wire  _io_storeAccessFault_T_33 = |(io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _T_30 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_31 = io__dmem_req_valid & _T_30; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  wire  _T_33 = _T_31 & _T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 534:39]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_10 = _T_31 | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_42 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  reg  r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_12 = _T_42 | r_1; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  assign io__in_ready = _io_dmem_req_valid_T | dtlbHasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 487:37]
  assign io__out_valid = dtlbHasException & state != 2'h0 | hasException | _io_out_valid_T_7; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 480:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 520:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:49]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 466:68]
  assign io__dmem_req_bits_size = {{1'd0}, size}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _reqWdata_T_18 | _reqWdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__dmem_resp_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 478:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 443:23]
  assign io__dtlbAF = DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 431:24]
  assign io__vaddr = _io_vaddr_T ? io__in_bits_src1 : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io__loadAccessFault = io__in_valid & _T_4 & ~(isStore | ISAMO2) & ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:68]
  assign io__storeAccessFault = _io_loadAccessFault_T_1 & (isStore & _io_loadAccessFault_T_31 | ISAMO2 & ~
    _io_storeAccessFault_T_33); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 532:45]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= io__in_bits_src1; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    addrLatch <= io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
      state <= 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    end else if (2'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (_T_1 & ~vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:45]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:53]
      end else if (_T_1 & vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:45]
        state <= 2'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:53]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (DTLBFINISH & ~dtlbHasException & scIsSuccess_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:61]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:69]
      end else begin
        state <= _GEN_3;
      end
    end else if (2'h2 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      state <= _GEN_5;
    end else begin
      state <= _GEN_6;
    end
    rdataLatch <= io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_10;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r_1 <= _GEN_12;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  addrLatch = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  rdataLatch = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AtomALU(
  input  [63:0] io_src1, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [63:0] io_src2, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [6:0]  io_func, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input         io_isWordOp, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  output [63:0] io_result // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
);
  wire  src1_signBit = io_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src1_T_1 = src1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src1_T_2 = {_src1_T_1,io_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src1 = io_isWordOp ? _src1_T_2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 183:17]
  wire  src2_signBit = io_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src2_T_1 = src2_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src2_T_2 = {_src2_T_1,io_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src2 = io_isWordOp ? _src2_T_2 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 184:17]
  wire  isAdderSub = ~io_func[6]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 186:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:39]
  wire [63:0] _adderRes_T_1 = src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:33]
  wire [64:0] _adderRes_T_2 = src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [63:0] xorRes = src1 ^ src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 188:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 189:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/LSU.scala 190:28]
  wire [63:0] _res_T_1 = src1 & src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 196:32]
  wire [63:0] _res_T_2 = src1 | src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 197:32]
  wire [63:0] _res_T_4 = slt ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 198:29]
  wire [63:0] _res_T_6 = slt ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 199:29]
  wire [63:0] _res_T_8 = sltu ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 200:29]
  wire [63:0] _res_T_10 = sltu ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 201:29]
  wire [64:0] _res_T_12 = 6'h22 == io_func[5:0] ? {{1'd0}, src2} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 6'h25 == io_func[5:0] ? {{1'd0}, _res_T_1} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 6'h26 == io_func[5:0] ? {{1'd0}, _res_T_2} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 6'h37 == io_func[5:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 6'h30 == io_func[5:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 6'h31 == io_func[5:0] ? {{1'd0}, _res_T_8} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  assign io_result = res[63:0]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 204:13]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src2, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [31:0] io__instr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        setLr_0,
  input         lr_0,
  output        scInflight_0,
  output        amoReq_0,
  input  [63:0] lr_addr,
  input  [55:0] dtlb_paddr,
  input         _T_12_0,
  input         scIsSuccess_0,
  output        setLrVal_0,
  input         vmEnable,
  input         DTLBFINISH,
  input         lsuMMIO_0,
  input         _T_13_1,
  output [63:0] setLrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__vaddr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_ISAMO2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBFINISH; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] atomALU_io_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [6:0] atomALU_io_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  atomALU_io_isWordOp; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  isAtomic = io__in_bits_func[5]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 54:38]
  wire  _isAmo_T_1 = io__in_bits_func == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _isAmo_T_4 = io__in_bits_func == 7'h21; // @[src/main/scala/nutcore/backend/fu/LSU.scala 58:37]
  wire  isAmo = isAtomic & ~_isAmo_T_1 & ~_isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/LSU.scala 59:61]
  wire [63:0] _in_vaddr_T_1 = io__in_bits_src1 + io__in_bits_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:43]
  wire [63:0] in_vaddr = isAtomic ? io__in_bits_src1 : _in_vaddr_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
  wire [1:0] _in_func_T_1 = io__instr[12] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:34]
  wire [1:0] in_func = isAtomic ? _in_func_T_1 : io__in_bits_func[1:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:20]
  wire  _addrAligned_T_1 = ~in_vaddr[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 69:29]
  wire  _addrAligned_T_3 = in_vaddr[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 70:32]
  wire  _addrAligned_T_5 = in_vaddr[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 71:32]
  wire  _addrAligned_T_6 = 2'h0 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_7 = 2'h1 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_8 = 2'h2 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_9 = 2'h3 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  addrAligned = _addrAligned_T_6 | _addrAligned_T_7 & _addrAligned_T_1 | _addrAligned_T_8 & _addrAligned_T_3 |
    _addrAligned_T_9 & _addrAligned_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  hasAddrMisaligned = io__in_valid & ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 73:36]
  wire  _io_loadAddrMisaligned_T_4 = ~io__in_bits_func[3] & ~isAtomic; // @[src/main/scala/nutcore/backend/fu/LSU.scala 56:49]
  wire  _hasScAccessFault_T_1 = ~vmEnable; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:46]
  wire  _hasScAccessFault_T_6 = |(in_vaddr >= 64'h80000000 & in_vaddr < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  hasScAccessFault = io__in_valid & _isAmo_T_4 & ~vmEnable & ~_hasScAccessFault_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:58]
  wire  valid = io__in_valid & addrAligned & ~hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 86:39]
  wire  _io_vaddr_T_2 = hasAddrMisaligned | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 91:44]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] _GEN_0 = _io_vaddr_T_2 ? in_vaddr : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  atomReq = valid & isAtomic; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 97:23]
  wire  amoReq = valid & isAmo; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:22]
  wire  lrReq = valid & _isAmo_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 99:21]
  wire  scReq = valid & _isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 100:21]
  wire [2:0] funct3 = io__instr[14:12]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 108:24]
  wire  scInvalid = scReq & (io__in_bits_src1 != lr_addr | ~lr_0) & _hasScAccessFault_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 126:53]
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
  reg [63:0] atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
  reg [63:0] atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
  wire  _T = 3'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _lsExecUnit_io_in_valid_T = ~atomReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 184:48]
  wire [2:0] _GEN_2 = amoReq ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 192:15 195:{19,26}]
  wire [2:0] _GEN_3 = lrReq ? 3'h3 : _GEN_2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 196:{18,25}]
  wire [2:0] _state_T = scInvalid ? 3'h0 : 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:31]
  wire  _T_1 = 3'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire [2:0] _GEN_5 = io__out_valid ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22 211:{26,33}]
  wire [1:0] _lsExecUnit_io_in_bits_func_T = funct3[0] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 231:40]
  wire  _T_14 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_6 = _T_14 ? 3'h6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 235:37 236:15 132:22]
  wire [3:0] _lsExecUnit_io_in_bits_func_T_1 = funct3[0] ? 4'hb : 4'ha; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 262:40]
  wire [2:0] _GEN_7 = _T_14 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 266:37 267:15 132:22]
  wire  _io_out_valid_T_5 = ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 293:63]
  wire  _io_out_valid_T_6 = _T_14 | ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 293:60]
  wire [2:0] _GEN_9 = _io_out_valid_T_6 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 294:51 295:15 132:22]
  wire  _GEN_16 = 3'h4 == state & (_T_14 | ~scIsSuccess_0); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 166:30 293:34]
  wire [2:0] _GEN_17 = 3'h4 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 132:22]
  wire  _GEN_18 = 3'h3 == state | 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 272:34]
  wire [3:0] _GEN_21 = 3'h3 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _lsExecUnit_io_in_bits_func_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 276:34]
  wire  _GEN_24 = 3'h3 == state ? _T_14 : _GEN_16; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 279:34]
  wire [2:0] _GEN_25 = 3'h3 == state ? _GEN_7 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_26 = 3'h7 == state | _GEN_18; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 258:34]
  wire [3:0] _GEN_29 = 3'h7 == state ? _lsExecUnit_io_in_bits_func_T_1 : _GEN_21; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 262:34]
  wire [63:0] _GEN_30 = 3'h7 == state ? atomMemReg : io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 263:34]
  wire  _GEN_32 = 3'h7 == state ? _T_14 : _GEN_24; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 265:34]
  wire [2:0] _GEN_33 = 3'h7 == state ? _GEN_7 : _GEN_25; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_34 = 3'h6 == state ? 1'h0 : _GEN_26; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 244:34]
  wire  _GEN_35 = 3'h6 == state ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 245:34]
  wire  _GEN_40 = 3'h6 == state ? 1'h0 : _GEN_32; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 251:34]
  wire [2:0] _GEN_41 = 3'h6 == state ? 3'h7 : _GEN_33; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 252:13]
  wire  _GEN_43 = 3'h5 == state | _GEN_34; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 227:34]
  wire  _GEN_44 = 3'h5 == state | _GEN_35; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 228:34]
  wire [3:0] _GEN_46 = 3'h5 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _GEN_29; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 231:34]
  wire  _GEN_49 = 3'h5 == state ? 1'h0 : _GEN_40; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 234:34]
  wire [2:0] _GEN_50 = 3'h5 == state ? _GEN_6 : _GEN_41; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_53 = 3'h1 == state | _GEN_43; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 202:34]
  wire  _GEN_54 = 3'h1 == state | _GEN_44; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 203:34]
  wire [6:0] _GEN_56 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_46}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 206:34]
  wire [63:0] _GEN_57 = 3'h1 == state ? io__wdata : _GEN_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 207:34]
  wire  _GEN_59 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_49; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 209:34]
  wire  _GEN_69 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_59; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 191:36]
  wire  _hasException_T_1 = lsExecUnit_io__dtlbAF | lsExecUnit_io__dtlbPF | io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 300:67]
  wire  _hasException_T_3 = _hasException_T_1 | io__storeAddrMisaligned | io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 301:53]
  wire  hasException = _hasException_T_3 | io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 302:24]
  wire [31:0] lr_paddr = dtlb_paddr[31:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 316:26]
  wire  _io_out_bits_T_1 = scInvalid | _io_out_valid_T_5; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:39]
  wire [63:0] _io_out_bits_T_3 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:59]
  reg  mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 318:24]
  wire  setLrVal = lrReq & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 319:21]
  wire [63:0] setLrAddr = vmEnable ? {{32'd0}, lr_paddr} : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 320:19]
  wire  scInflight = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 143:23]
  LSExecUnit lsExecUnit ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_ready(lsExecUnit_io__in_ready),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__dtlbAF(lsExecUnit_io__dtlbAF),
    .io__vaddr(lsExecUnit_io__vaddr),
    .io__loadAccessFault(lsExecUnit_io__loadAccessFault),
    .io__storeAccessFault(lsExecUnit_io__storeAccessFault),
    .DTLBPF(lsExecUnit_DTLBPF),
    .scIsSuccess_0(lsExecUnit_scIsSuccess_0),
    .vmEnable_0(lsExecUnit_vmEnable_0),
    .ISAMO2(lsExecUnit_ISAMO2),
    .DTLBFINISH(lsExecUnit_DTLBFINISH),
    .DTLBAF(lsExecUnit_DTLBAF)
  );
  AtomALU atomALU ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__out_valid = hasException | _GEN_69; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23 305:18]
  assign io__out_bits = scReq ? {{63'd0}, _io_out_bits_T_1} : _io_out_bits_T_3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:21]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__isMMIO = mmioReg & io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 332:24]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 94:13]
  assign io__dtlbAF = lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:13]
  assign io__vaddr = io__loadAddrMisaligned | io__storeAddrMisaligned | hasScAccessFault ? _GEN_0 : lsExecUnit_io__vaddr
    ; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 90:18]
  assign io__loadAddrMisaligned = hasAddrMisaligned & (_io_loadAddrMisaligned_T_4 | _isAmo_T_1); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 74:46]
  assign io__storeAddrMisaligned = hasAddrMisaligned & (io__in_bits_func[3] | isAmo | _isAmo_T_4); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 75:47]
  assign io__loadAccessFault = lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 334:22]
  assign io__storeAccessFault = lsExecUnit_io__storeAccessFault | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:57]
  assign setLr_0 = setLr;
  assign scInflight_0 = scInflight;
  assign amoReq_0 = amoReq;
  assign setLrVal_0 = setLrVal;
  assign setLrAddr_0 = setLrAddr;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? valid & ~atomReq : _GEN_53; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 184:36]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _in_vaddr_T_1 : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 186:36]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_56; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 188:36]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_54; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 185:36]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_57; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 189:36]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_DTLBPF = _T_12_0;
  assign lsExecUnit_scIsSuccess_0 = scIsSuccess_0;
  assign lsExecUnit_vmEnable_0 = vmEnable;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign lsExecUnit_DTLBAF = _T_13_1;
  assign atomALU_io_src1 = atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 136:19]
  assign atomALU_io_src2 = io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 137:19]
  assign atomALU_io_func = io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 138:19]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 110:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T_2) begin // @[src/main/scala/utils/Hold.scala 23:65]
      if (isAtomic) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
        io_vaddr_r <= io__in_bits_src1;
      end else begin
        io_vaddr_r <= _in_vaddr_T_1;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 304:11]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (scReq) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:18]
        state <= _state_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:25]
      end else begin
        state <= _GEN_3;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      state <= _GEN_5;
    end else begin
      state <= _GEN_50;
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 239:18]
        end else if (3'h6 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 253:18]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomRegReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 240:18]
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
    end else if (io__out_valid) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:23]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:33]
    end else if (~mmioReg) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:19]
      mmioReg <= lsuMMIO_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:29]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & _T_1 & ~reset & ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:210 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  atomMemReg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  atomRegReg = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  mmioReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~_T & _T_1 & ~reset) begin
      assert(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
    end
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output [129:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [64:0] mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [129:0] io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg [129:0] io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg [129:0] io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg  io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg  io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg  io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21 63:{31,38}]
  assign io_in_ready = ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 65:49]
  assign io_out_valid = io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 60:16]
  assign io_out_bits = io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 59:37]
  always @(posedge clock) begin
    mulRes_REG <= io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    mulRes_REG_1 <= io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    io_out_bits_REG <= $signed(mulRes_REG) * $signed(mulRes_REG_1); // @[src/main/scala/nutcore/backend/fu/MDU.scala 58:49]
    io_out_bits_REG_1 <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_bits_REG_2 <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    io_out_valid_REG <= io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    io_out_valid_REG_1 <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    io_out_valid_REG_2 <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_valid_REG_3 <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end else if (io_out_valid) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:23]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:30]
    end else begin
      busy <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  mulRes_REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  mulRes_REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  io_out_bits_REG = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  io_out_bits_REG_1 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  io_out_bits_REG_2 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_sign, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output [127:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  _newReq_T_1 = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  newReq = state == 3'h0 & _newReq_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 81:18]
  reg [128:0] shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_1 = 64'h0 - io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_1 : io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_3 = 64'h0 - io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  reg  aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  reg  qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  reg [63:0] bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire [64:0] _aValx2Reg_T = {aVal,1'h0}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:32]
  reg [64:0] aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  reg [5:0] cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [31:0] canSkipShift_hi = bReg[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo = bReg[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi = |canSkipShift_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_1 = canSkipShift_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_1 = canSkipShift_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_1 = |canSkipShift_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_2 = canSkipShift_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_2 = canSkipShift_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_2 = |canSkipShift_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_3 = canSkipShift_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_3 = canSkipShift_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_3 = |canSkipShift_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_3 = canSkipShift_hi_3[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_4 = canSkipShift_hi_3[3] ? 2'h3 : _canSkipShift_T_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_8 = canSkipShift_lo_3[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_9 = canSkipShift_lo_3[3] ? 2'h3 : _canSkipShift_T_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_10 = canSkipShift_useHi_3 ? _canSkipShift_T_4 : _canSkipShift_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_11 = {canSkipShift_useHi_3,_canSkipShift_T_10}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_4 = canSkipShift_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_4 = canSkipShift_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_4 = |canSkipShift_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_15 = canSkipShift_hi_4[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_16 = canSkipShift_hi_4[3] ? 2'h3 : _canSkipShift_T_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_20 = canSkipShift_lo_4[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_21 = canSkipShift_lo_4[3] ? 2'h3 : _canSkipShift_T_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_22 = canSkipShift_useHi_4 ? _canSkipShift_T_16 : _canSkipShift_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_23 = {canSkipShift_useHi_4,_canSkipShift_T_22}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_24 = canSkipShift_useHi_2 ? _canSkipShift_T_11 : _canSkipShift_T_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_25 = {canSkipShift_useHi_2,_canSkipShift_T_24}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_5 = canSkipShift_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_5 = canSkipShift_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_5 = |canSkipShift_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_6 = canSkipShift_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_6 = canSkipShift_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_6 = |canSkipShift_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_29 = canSkipShift_hi_6[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_30 = canSkipShift_hi_6[3] ? 2'h3 : _canSkipShift_T_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_34 = canSkipShift_lo_6[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_35 = canSkipShift_lo_6[3] ? 2'h3 : _canSkipShift_T_34; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_36 = canSkipShift_useHi_6 ? _canSkipShift_T_30 : _canSkipShift_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_37 = {canSkipShift_useHi_6,_canSkipShift_T_36}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_7 = canSkipShift_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_7 = canSkipShift_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_7 = |canSkipShift_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_41 = canSkipShift_hi_7[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_42 = canSkipShift_hi_7[3] ? 2'h3 : _canSkipShift_T_41; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_46 = canSkipShift_lo_7[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_47 = canSkipShift_lo_7[3] ? 2'h3 : _canSkipShift_T_46; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_48 = canSkipShift_useHi_7 ? _canSkipShift_T_42 : _canSkipShift_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_49 = {canSkipShift_useHi_7,_canSkipShift_T_48}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_50 = canSkipShift_useHi_5 ? _canSkipShift_T_37 : _canSkipShift_T_49; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_51 = {canSkipShift_useHi_5,_canSkipShift_T_50}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_52 = canSkipShift_useHi_1 ? _canSkipShift_T_25 : _canSkipShift_T_51; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_53 = {canSkipShift_useHi_1,_canSkipShift_T_52}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_8 = canSkipShift_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_8 = canSkipShift_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_8 = |canSkipShift_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_9 = canSkipShift_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_9 = canSkipShift_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_9 = |canSkipShift_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_10 = canSkipShift_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_10 = canSkipShift_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_10 = |canSkipShift_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_57 = canSkipShift_hi_10[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_58 = canSkipShift_hi_10[3] ? 2'h3 : _canSkipShift_T_57; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_62 = canSkipShift_lo_10[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_63 = canSkipShift_lo_10[3] ? 2'h3 : _canSkipShift_T_62; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_64 = canSkipShift_useHi_10 ? _canSkipShift_T_58 : _canSkipShift_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_65 = {canSkipShift_useHi_10,_canSkipShift_T_64}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_11 = canSkipShift_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_11 = canSkipShift_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_11 = |canSkipShift_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_69 = canSkipShift_hi_11[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_70 = canSkipShift_hi_11[3] ? 2'h3 : _canSkipShift_T_69; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_74 = canSkipShift_lo_11[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_75 = canSkipShift_lo_11[3] ? 2'h3 : _canSkipShift_T_74; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_76 = canSkipShift_useHi_11 ? _canSkipShift_T_70 : _canSkipShift_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_77 = {canSkipShift_useHi_11,_canSkipShift_T_76}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_78 = canSkipShift_useHi_9 ? _canSkipShift_T_65 : _canSkipShift_T_77; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_79 = {canSkipShift_useHi_9,_canSkipShift_T_78}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_12 = canSkipShift_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_12 = canSkipShift_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_12 = |canSkipShift_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_13 = canSkipShift_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_13 = canSkipShift_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_13 = |canSkipShift_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_83 = canSkipShift_hi_13[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_84 = canSkipShift_hi_13[3] ? 2'h3 : _canSkipShift_T_83; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_88 = canSkipShift_lo_13[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_89 = canSkipShift_lo_13[3] ? 2'h3 : _canSkipShift_T_88; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_90 = canSkipShift_useHi_13 ? _canSkipShift_T_84 : _canSkipShift_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_91 = {canSkipShift_useHi_13,_canSkipShift_T_90}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_14 = canSkipShift_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_14 = canSkipShift_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_14 = |canSkipShift_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_95 = canSkipShift_hi_14[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_96 = canSkipShift_hi_14[3] ? 2'h3 : _canSkipShift_T_95; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_100 = canSkipShift_lo_14[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_101 = canSkipShift_lo_14[3] ? 2'h3 : _canSkipShift_T_100; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_102 = canSkipShift_useHi_14 ? _canSkipShift_T_96 : _canSkipShift_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_103 = {canSkipShift_useHi_14,_canSkipShift_T_102}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_104 = canSkipShift_useHi_12 ? _canSkipShift_T_91 : _canSkipShift_T_103; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_105 = {canSkipShift_useHi_12,_canSkipShift_T_104}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_106 = canSkipShift_useHi_8 ? _canSkipShift_T_79 : _canSkipShift_T_105; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_107 = {canSkipShift_useHi_8,_canSkipShift_T_106}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_108 = canSkipShift_useHi ? _canSkipShift_T_53 : _canSkipShift_T_107; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_109 = {canSkipShift_useHi,_canSkipShift_T_108}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] _GEN_18 = {{1'd0}, _canSkipShift_T_109}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire [6:0] _canSkipShift_T_110 = 7'h40 | _GEN_18; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire  canSkipShift_hi_15 = aValx2Reg[64]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [63:0] canSkipShift_lo_15 = aValx2Reg[63:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_15 = |canSkipShift_hi_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [31:0] canSkipShift_hi_16 = canSkipShift_lo_15[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo_16 = canSkipShift_lo_15[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_16 = |canSkipShift_hi_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_17 = canSkipShift_hi_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_17 = canSkipShift_hi_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_17 = |canSkipShift_hi_17; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_18 = canSkipShift_hi_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_18 = canSkipShift_hi_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_18 = |canSkipShift_hi_18; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_19 = canSkipShift_hi_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_19 = canSkipShift_hi_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_19 = |canSkipShift_hi_19; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_114 = canSkipShift_hi_19[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_115 = canSkipShift_hi_19[3] ? 2'h3 : _canSkipShift_T_114; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_119 = canSkipShift_lo_19[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_120 = canSkipShift_lo_19[3] ? 2'h3 : _canSkipShift_T_119; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_121 = canSkipShift_useHi_19 ? _canSkipShift_T_115 : _canSkipShift_T_120; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_122 = {canSkipShift_useHi_19,_canSkipShift_T_121}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_20 = canSkipShift_lo_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_20 = canSkipShift_lo_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_20 = |canSkipShift_hi_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_126 = canSkipShift_hi_20[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_127 = canSkipShift_hi_20[3] ? 2'h3 : _canSkipShift_T_126; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_131 = canSkipShift_lo_20[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_132 = canSkipShift_lo_20[3] ? 2'h3 : _canSkipShift_T_131; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_133 = canSkipShift_useHi_20 ? _canSkipShift_T_127 : _canSkipShift_T_132; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_134 = {canSkipShift_useHi_20,_canSkipShift_T_133}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_135 = canSkipShift_useHi_18 ? _canSkipShift_T_122 : _canSkipShift_T_134; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_136 = {canSkipShift_useHi_18,_canSkipShift_T_135}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_21 = canSkipShift_lo_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_21 = canSkipShift_lo_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_21 = |canSkipShift_hi_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_22 = canSkipShift_hi_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_22 = canSkipShift_hi_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_22 = |canSkipShift_hi_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_140 = canSkipShift_hi_22[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_141 = canSkipShift_hi_22[3] ? 2'h3 : _canSkipShift_T_140; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_145 = canSkipShift_lo_22[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_146 = canSkipShift_lo_22[3] ? 2'h3 : _canSkipShift_T_145; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_147 = canSkipShift_useHi_22 ? _canSkipShift_T_141 : _canSkipShift_T_146; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_148 = {canSkipShift_useHi_22,_canSkipShift_T_147}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_23 = canSkipShift_lo_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_23 = canSkipShift_lo_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_23 = |canSkipShift_hi_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_152 = canSkipShift_hi_23[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_153 = canSkipShift_hi_23[3] ? 2'h3 : _canSkipShift_T_152; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_157 = canSkipShift_lo_23[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_158 = canSkipShift_lo_23[3] ? 2'h3 : _canSkipShift_T_157; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_159 = canSkipShift_useHi_23 ? _canSkipShift_T_153 : _canSkipShift_T_158; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_160 = {canSkipShift_useHi_23,_canSkipShift_T_159}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_161 = canSkipShift_useHi_21 ? _canSkipShift_T_148 : _canSkipShift_T_160; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_162 = {canSkipShift_useHi_21,_canSkipShift_T_161}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_163 = canSkipShift_useHi_17 ? _canSkipShift_T_136 : _canSkipShift_T_162; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_164 = {canSkipShift_useHi_17,_canSkipShift_T_163}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_24 = canSkipShift_lo_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_24 = canSkipShift_lo_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_24 = |canSkipShift_hi_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_25 = canSkipShift_hi_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_25 = canSkipShift_hi_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_25 = |canSkipShift_hi_25; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_26 = canSkipShift_hi_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_26 = canSkipShift_hi_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_26 = |canSkipShift_hi_26; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_168 = canSkipShift_hi_26[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_169 = canSkipShift_hi_26[3] ? 2'h3 : _canSkipShift_T_168; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_173 = canSkipShift_lo_26[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_174 = canSkipShift_lo_26[3] ? 2'h3 : _canSkipShift_T_173; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_175 = canSkipShift_useHi_26 ? _canSkipShift_T_169 : _canSkipShift_T_174; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_176 = {canSkipShift_useHi_26,_canSkipShift_T_175}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_27 = canSkipShift_lo_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_27 = canSkipShift_lo_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_27 = |canSkipShift_hi_27; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_180 = canSkipShift_hi_27[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_181 = canSkipShift_hi_27[3] ? 2'h3 : _canSkipShift_T_180; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_185 = canSkipShift_lo_27[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_186 = canSkipShift_lo_27[3] ? 2'h3 : _canSkipShift_T_185; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_187 = canSkipShift_useHi_27 ? _canSkipShift_T_181 : _canSkipShift_T_186; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_188 = {canSkipShift_useHi_27,_canSkipShift_T_187}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_189 = canSkipShift_useHi_25 ? _canSkipShift_T_176 : _canSkipShift_T_188; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_190 = {canSkipShift_useHi_25,_canSkipShift_T_189}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_28 = canSkipShift_lo_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_28 = canSkipShift_lo_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_28 = |canSkipShift_hi_28; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_29 = canSkipShift_hi_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_29 = canSkipShift_hi_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_29 = |canSkipShift_hi_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_194 = canSkipShift_hi_29[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_195 = canSkipShift_hi_29[3] ? 2'h3 : _canSkipShift_T_194; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_199 = canSkipShift_lo_29[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_200 = canSkipShift_lo_29[3] ? 2'h3 : _canSkipShift_T_199; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_201 = canSkipShift_useHi_29 ? _canSkipShift_T_195 : _canSkipShift_T_200; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_202 = {canSkipShift_useHi_29,_canSkipShift_T_201}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_30 = canSkipShift_lo_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_30 = canSkipShift_lo_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_30 = |canSkipShift_hi_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_206 = canSkipShift_hi_30[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_207 = canSkipShift_hi_30[3] ? 2'h3 : _canSkipShift_T_206; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_211 = canSkipShift_lo_30[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_212 = canSkipShift_lo_30[3] ? 2'h3 : _canSkipShift_T_211; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_213 = canSkipShift_useHi_30 ? _canSkipShift_T_207 : _canSkipShift_T_212; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_214 = {canSkipShift_useHi_30,_canSkipShift_T_213}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_215 = canSkipShift_useHi_28 ? _canSkipShift_T_202 : _canSkipShift_T_214; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_216 = {canSkipShift_useHi_28,_canSkipShift_T_215}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_217 = canSkipShift_useHi_24 ? _canSkipShift_T_190 : _canSkipShift_T_216; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_218 = {canSkipShift_useHi_24,_canSkipShift_T_217}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_219 = canSkipShift_useHi_16 ? _canSkipShift_T_164 : _canSkipShift_T_218; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_220 = {canSkipShift_useHi_16,_canSkipShift_T_219}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _canSkipShift_T_221 = canSkipShift_useHi_15 ? 6'h0 : _canSkipShift_T_220; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [6:0] _canSkipShift_T_222 = {canSkipShift_useHi_15,_canSkipShift_T_221}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] canSkipShift = _canSkipShift_T_110 - _canSkipShift_T_222; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:45]
  wire [6:0] _value_T_1 = canSkipShift >= 7'h3f ? 7'h3f : canSkipShift; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:21]
  wire [127:0] _GEN_22 = {{63'd0}, aValx2Reg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [127:0] _shiftReg_T = _GEN_22 << cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [64:0] _GEN_19 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire  enough = hi >= _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire [64:0] _shiftReg_T_2 = hi - _GEN_19; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_3 = enough ? _shiftReg_T_2 : hi; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:24]
  wire [128:0] _shiftReg_T_5 = {_shiftReg_T_3[63:0],lo,enough}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:20]
  wire [5:0] _value_T_4 = cnt_value + 6'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_4 = cnt_value == 6'h3f ? 3'h4 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 118:{36,44} 77:22]
  wire [2:0] _GEN_5 = state == 3'h4 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
  wire [5:0] _GEN_11 = state == 3'h2 ? cnt_value : _GEN_7; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:15 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, cnt_value} : _GEN_12; // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] r = hi[64:1]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 123:13]
  wire [63:0] _resQ_T_1 = 64'h0 - lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _resQ_T_1 : lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:17]
  wire [63:0] _resR_T_1 = 64'h0 - r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _resR_T_1 : r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:17]
  wire [6:0] _GEN_21 = reset ? 7'h0 : _GEN_16; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  assign io_in_ready = state == 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 126:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end else if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      state <= 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
      state <= 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
      state <= 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 113:11]
    end else begin
      state <= _GEN_8;
    end
    if (!(newReq)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
        if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
          shiftReg <= {{1'd0}, _shiftReg_T}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
          shiftReg <= _shiftReg_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
      aSignReg <= aSign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
      qSignReg <= (aSign ^ bSign) & ~divBy0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
      if (bSign) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
        bReg <= _T_3;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
      aValx2Reg <= _aValx2Reg_T; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    cnt_value <= _GEN_21[5:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  cnt_value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output [63:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  div_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 43:25]
  wire [64:0] _mul_io_in_bits_0_T_1 = {1'h0,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_0_signBit = io_in_bits_src1[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_0_T_2 = {mul_io_in_bits_0_signBit,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _mul_io_in_bits_0_T_5 = 2'h0 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_6 = 2'h1 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_7 = 2'h2 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_8 = 2'h3 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [64:0] _mul_io_in_bits_0_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_13 = _mul_io_in_bits_0_T_9 | _mul_io_in_bits_0_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_14 = _mul_io_in_bits_0_T_13 | _mul_io_in_bits_0_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_1 = {1'h0,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_1_signBit = io_in_bits_src2[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_1_T_2 = {mul_io_in_bits_1_signBit,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] _mul_io_in_bits_1_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_1_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_13 = _mul_io_in_bits_1_T_9 | _mul_io_in_bits_1_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_14 = _mul_io_in_bits_1_T_13 | _mul_io_in_bits_1_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  div_io_in_bits_0_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_0_T_1 = div_io_in_bits_0_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_0_T_2 = {_div_io_in_bits_0_T_1,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_0_T_4 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_0_T_5 = isDivSign ? _div_io_in_bits_0_T_2 : _div_io_in_bits_0_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire  div_io_in_bits_1_signBit = io_in_bits_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_1_T_1 = div_io_in_bits_1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_1_T_2 = {_div_io_in_bits_1_T_1,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_1_T_4 = {32'h0,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_1_T_5 = isDivSign ? _div_io_in_bits_1_T_2 : _div_io_in_bits_1_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[src/main/scala/nutcore/backend/fu/MDU.scala 178:16]
  wire  io_out_bits_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _io_out_bits_T_1 = io_out_bits_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_T_2 = {_io_out_bits_T_1,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
  wire  isDivReg = _isDivReg_T ? isDiv : isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:21]
  wire  _T = mul_io_out_ready & mul_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  Multiplier mul ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 183:22]
  assign io_out_bits = isW ? _io_out_bits_T_2 : res; // @[src/main/scala/nutcore/backend/fu/MDU.scala 179:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 173:34]
  assign mul_io_in_bits_0 = _mul_io_in_bits_0_T_14 | _mul_io_in_bits_0_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_in_bits_1 = _mul_io_in_bits_1_T_14 | _mul_io_in_bits_1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _div_io_in_bits_0_T_5 : io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _div_io_in_bits_1_T_5 : io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  always @(posedge clock) begin
    isDivReg_REG <= io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg_REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_1(
  input         clock,
  input  [63:0] io_bits_privilegeMode, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mcause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_scause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_satp, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mie, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mideleg, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_medeleg // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mcause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_scause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_satp; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mie; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mideleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_medeleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestCSRState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_privilegeMode(dpic_io_privilegeMode),
    .io_mstatus(dpic_io_mstatus),
    .io_sstatus(dpic_io_sstatus),
    .io_mepc(dpic_io_mepc),
    .io_sepc(dpic_io_sepc),
    .io_mtval(dpic_io_mtval),
    .io_stval(dpic_io_stval),
    .io_mtvec(dpic_io_mtvec),
    .io_stvec(dpic_io_stvec),
    .io_mcause(dpic_io_mcause),
    .io_scause(dpic_io_scause),
    .io_satp(dpic_io_satp),
    .io_mip(dpic_io_mip),
    .io_mie(dpic_io_mie),
    .io_mscratch(dpic_io_mscratch),
    .io_sscratch(dpic_io_sscratch),
    .io_mideleg(dpic_io_mideleg),
    .io_medeleg(dpic_io_medeleg),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_privilegeMode = io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mstatus = io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sstatus = io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mepc = io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sepc = io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtval = io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stval = io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtvec = io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stvec = io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mcause = io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_scause = io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_satp = io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mip = io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mie = io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mscratch = io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sscratch = io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mideleg = io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_medeleg = io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_2(
  input         clock,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_interrupt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exception, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_exceptionPC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exceptionInst // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_interrupt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exception; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_interrupt(dpic_io_interrupt),
    .io_exception(dpic_io_exception),
    .io_exceptionPC(dpic_io_exceptionPC),
    .io_exceptionInst(dpic_io_exceptionInst),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_interrupt = io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exception = io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionPC = io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionInst = io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module CSRDiffWrapper(
  input         clock,
  input  [63:0] io_csrState_privilegeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_sstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_sepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mtval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_stval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mtvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_stvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mcause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_scause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_satp, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mip, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mie, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_sscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_mideleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_csrState_medeleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input         io_archEvent_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [31:0] io_archEvent_interrupt, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [31:0] io_archEvent_exception, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [63:0] io_archEvent_exceptionPC, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
  input  [31:0] io_archEvent_exceptionInst // @[src/main/scala/nutcore/backend/fu/CSR.scala 1049:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftestArchEvent_module_io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] difftest_REG_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg [63:0] difftest_REG_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
  reg  difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
  reg [31:0] difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
  reg [31:0] difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
  reg [63:0] difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
  reg [31:0] difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
  reg  difftestArchEvent_REG_1_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  reg [31:0] difftestArchEvent_REG_1_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  reg [31:0] difftestArchEvent_REG_1_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  reg [63:0] difftestArchEvent_REG_1_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  reg [31:0] difftestArchEvent_REG_1_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  DummyDPICWrapper_1 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .io_bits_privilegeMode(difftest_module_io_bits_privilegeMode),
    .io_bits_mstatus(difftest_module_io_bits_mstatus),
    .io_bits_sstatus(difftest_module_io_bits_sstatus),
    .io_bits_mepc(difftest_module_io_bits_mepc),
    .io_bits_sepc(difftest_module_io_bits_sepc),
    .io_bits_mtval(difftest_module_io_bits_mtval),
    .io_bits_stval(difftest_module_io_bits_stval),
    .io_bits_mtvec(difftest_module_io_bits_mtvec),
    .io_bits_stvec(difftest_module_io_bits_stvec),
    .io_bits_mcause(difftest_module_io_bits_mcause),
    .io_bits_scause(difftest_module_io_bits_scause),
    .io_bits_satp(difftest_module_io_bits_satp),
    .io_bits_mip(difftest_module_io_bits_mip),
    .io_bits_mie(difftest_module_io_bits_mie),
    .io_bits_mscratch(difftest_module_io_bits_mscratch),
    .io_bits_sscratch(difftest_module_io_bits_sscratch),
    .io_bits_mideleg(difftest_module_io_bits_mideleg),
    .io_bits_medeleg(difftest_module_io_bits_medeleg)
  );
  DummyDPICWrapper_2 difftestArchEvent_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftestArchEvent_module_clock),
    .io_valid(difftestArchEvent_module_io_valid),
    .io_bits_valid(difftestArchEvent_module_io_bits_valid),
    .io_bits_interrupt(difftestArchEvent_module_io_bits_interrupt),
    .io_bits_exception(difftestArchEvent_module_io_bits_exception),
    .io_bits_exceptionPC(difftestArchEvent_module_io_bits_exceptionPC),
    .io_bits_exceptionInst(difftestArchEvent_module_io_bits_exceptionInst)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_io_bits_privilegeMode = difftest_REG_privilegeMode; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mstatus = difftest_REG_mstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_sstatus = difftest_REG_sstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mepc = difftest_REG_mepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_sepc = difftest_REG_sepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mtval = difftest_REG_mtval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_stval = difftest_REG_stval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mtvec = difftest_REG_mtvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_stvec = difftest_REG_stvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mcause = difftest_REG_mcause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_scause = difftest_REG_scause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_satp = difftest_REG_satp; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mip = difftest_REG_mip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mie = difftest_REG_mie; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mscratch = difftest_REG_mscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_sscratch = difftest_REG_sscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_mideleg = difftest_REG_mideleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftest_module_io_bits_medeleg = difftest_REG_medeleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1055:16]
  assign difftestArchEvent_module_clock = clock;
  assign difftestArchEvent_module_io_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  assign difftestArchEvent_module_io_bits_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  assign difftestArchEvent_module_io_bits_interrupt = difftestArchEvent_REG_1_interrupt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  assign difftestArchEvent_module_io_bits_exception = difftestArchEvent_REG_1_exception; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  assign difftestArchEvent_module_io_bits_exceptionPC = difftestArchEvent_REG_1_exceptionPC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  assign difftestArchEvent_module_io_bits_exceptionInst = difftestArchEvent_REG_1_exceptionInst; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1059:25]
  always @(posedge clock) begin
    difftest_REG_privilegeMode <= io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mstatus <= io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_sstatus <= io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mepc <= io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_sepc <= io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mtval <= io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_stval <= io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mtvec <= io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_stvec <= io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mcause <= io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_scause <= io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_satp <= io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mip <= io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mie <= io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mscratch <= io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_sscratch <= io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_mideleg <= io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftest_REG_medeleg <= io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1055:26]
    difftestArchEvent_REG_valid <= io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
    difftestArchEvent_REG_interrupt <= io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
    difftestArchEvent_REG_exception <= io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
    difftestArchEvent_REG_exceptionPC <= io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
    difftestArchEvent_REG_exceptionInst <= io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:43]
    difftestArchEvent_REG_1_valid <= difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
    difftestArchEvent_REG_1_interrupt <= difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
    difftestArchEvent_REG_1_exception <= difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
    difftestArchEvent_REG_1_exceptionPC <= difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
    difftestArchEvent_REG_1_exceptionInst <= difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1059:35]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_REG_privilegeMode = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  difftest_REG_mstatus = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_sstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  difftest_REG_mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  difftest_REG_sepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  difftest_REG_mtval = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_stval = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  difftest_REG_mtvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  difftest_REG_stvec = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  difftest_REG_mcause = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  difftest_REG_scause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  difftest_REG_satp = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  difftest_REG_mip = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  difftest_REG_mie = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  difftest_REG_mscratch = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  difftest_REG_sscratch = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  difftest_REG_mideleg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  difftest_REG_medeleg = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  difftestArchEvent_REG_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  difftestArchEvent_REG_interrupt = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  difftestArchEvent_REG_exception = _RAND_20[31:0];
  _RAND_21 = {2{`RANDOM}};
  difftestArchEvent_REG_exceptionPC = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  difftestArchEvent_REG_exceptionInst = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  difftestArchEvent_REG_1_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  difftestArchEvent_REG_1_interrupt = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exception = _RAND_25[31:0];
  _RAND_26 = {2{`RANDOM}};
  difftestArchEvent_REG_1_exceptionPC = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exceptionInst = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_12, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_13, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_15, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_3, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_9, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_11, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_crossBoundaryFault, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_instrValid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_illegalJump_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_illegalJump_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_dmemExceptionAddr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_xretIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_xretIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_xretIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_imemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_dmemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_sum, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_mxr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_loadPF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_storePF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_laf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_saf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wenFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isPerfRead, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isExit, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_vmEnable, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_rfWenReal, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         set_lr,
  output        lr_0,
  input         meip_0,
  output [63:0] lrAddr_0,
  output [63:0] satp_0,
  input         mtip_0,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [11:0] intrVecIDU_0,
  input  [63:0] set_lr_addr,
  input         msip_0,
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  wire  CSRDiffWrapper_clock; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire  CSRDiffWrapper_io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [63:0] CSRDiffWrapper_io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
  reg [1:0] priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
  reg [63:0] mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
  reg [63:0] mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
  reg [63:0] mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
  reg [63:0] mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
  reg [63:0] mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
  reg [63:0] mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
  reg [63:0] mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
  wire [11:0] _mip_T = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:22]
  wire [63:0] _GEN_85 = {{52'd0}, _mip_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire [63:0] _mip_T_1 = _GEN_85 | mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire  mip_s_u = _mip_T_1[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_s = _mip_T_1[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_h = _mip_T_1[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_m = _mip_T_1[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_u = _mip_T_1[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_s = _mip_T_1[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_h = _mip_T_1[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_m = _mip_T_1[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_u = _mip_T_1[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_s = _mip_T_1[9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_h = _mip_T_1[10]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_m = _mip_T_1[11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  reg [63:0] mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  reg [63:0] medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
  reg [63:0] mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
  reg [63:0] mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
  reg [63:0] stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 379:32]
  reg [63:0] satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
  wire [3:0] satpStruct_mode = satp[63:60]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 384:33]
  wire  _vmEnable_T_1 = priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:38]
  wire  vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  reg [63:0] sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
  reg [63:0] scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
  reg [63:0] stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
  reg [63:0] sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
  reg [63:0] scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
  reg  lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
  reg [63:0] lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
  reg [63:0] perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [5:0] lo = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] _T_25 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 507:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdata_T_29 = 12'hf12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_30 = 12'h180 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_59 = _rdata_T_30 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_31 = 12'h140 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_60 = _rdata_T_31 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_88 = _rdata_T_59 | _rdata_T_60; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_32 = 12'h306 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_61 = _rdata_T_32 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_89 = _rdata_T_88 | _rdata_T_61; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_33 = 12'hf11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_34 = 12'h104 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_5 = mie & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_63 = _rdata_T_34 ? _rdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_91 = _rdata_T_89 | _rdata_T_63; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_35 = 12'h144 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _GEN_86 = {{52'd0}, _T_25}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_6 = _GEN_86 & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_64 = _rdata_T_35 ? _rdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_92 = _rdata_T_91 | _rdata_T_64; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_36 = 12'h100 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_7 = mstatus & 64'h80000003000d8122; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_65 = _rdata_T_36 ? _rdata_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_93 = _rdata_T_92 | _rdata_T_65; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_37 = 12'h305 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_66 = _rdata_T_37 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_94 = _rdata_T_93 | _rdata_T_66; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_38 = 12'h300 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_9 = mstatus & 64'h8000000f007ff9aa; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_67 = _rdata_T_38 ? _rdata_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_95 = _rdata_T_94 | _rdata_T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_39 = 12'hf13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_40 = 12'h340 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_69 = _rdata_T_40 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_97 = _rdata_T_95 | _rdata_T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_41 = 12'h142 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_70 = _rdata_T_41 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_98 = _rdata_T_97 | _rdata_T_70; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_42 = 12'h302 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_71 = _rdata_T_42 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_99 = _rdata_T_98 | _rdata_T_71; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_43 = 12'h105 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_72 = _rdata_T_43 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_100 = _rdata_T_99 | _rdata_T_72; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_44 = 12'h141 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_73 = _rdata_T_44 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_101 = _rdata_T_100 | _rdata_T_73; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_45 = 12'h342 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_74 = _rdata_T_45 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_102 = _rdata_T_101 | _rdata_T_74; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_46 = 12'h304 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_75 = _rdata_T_46 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_103 = _rdata_T_102 | _rdata_T_75; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_47 = 12'hb01 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_76 = _rdata_T_47 ? perfCnts_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_104 = _rdata_T_103 | _rdata_T_76; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_48 = 12'h143 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_77 = _rdata_T_48 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_105 = _rdata_T_104 | _rdata_T_77; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_49 = 12'h301 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_78 = _rdata_T_49 ? 64'h8000000000141105 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_106 = _rdata_T_105 | _rdata_T_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_50 = 12'hb00 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_79 = _rdata_T_50 ? perfCnts_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_107 = _rdata_T_106 | _rdata_T_79; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_51 = 12'h344 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_80 = _rdata_T_51 ? _GEN_86 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_108 = _rdata_T_107 | _rdata_T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_52 = 12'hb02 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_81 = _rdata_T_52 ? perfCnts_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_109 = _rdata_T_108 | _rdata_T_81; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_53 = 12'h303 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_82 = _rdata_T_53 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_110 = _rdata_T_109 | _rdata_T_82; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_54 = 12'hf14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_55 = 12'h341 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_84 = _rdata_T_55 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_112 = _rdata_T_110 | _rdata_T_84; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_56 = 12'h343 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_85 = _rdata_T_56 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_85; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_57 = 12'h106 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_86 = _rdata_T_57 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 512:30]
  wire [63:0] _wdata_T_1 = ~io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:33]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:30]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 515:30]
  wire [63:0] _wdata_T_4 = ~csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:33]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:30]
  wire  _wdata_T_6 = 7'h1 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_7 = 7'h2 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_8 = 7'h3 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_9 = 7'h5 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_10 = 7'h6 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_11 = 7'h7 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_in_bits_src1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 522:69]
  wire [7:0] wen_lo = {io_cfIn_exceptionVec_7,io_cfIn_exceptionVec_6,io_cfIn_exceptionVec_5,io_cfIn_exceptionVec_4,1'h0,
    io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire [15:0] _wen_T = {io_cfIn_exceptionVec_15,1'h0,io_cfIn_exceptionVec_13,io_cfIn_exceptionVec_12,4'h0,wen_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire  _wen_T_2 = ~(|_wen_T); // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:23]
  wire  _wen_T_4 = io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:64]
  wire  wen = io_in_valid & ~(|_wen_T) & io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:56]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 526:39]
  wire  isCSRRS = io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 531:40]
  wire  isCSRRC = io_in_bits_func == 7'h3 | io_in_bits_func == 7'h7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 532:40]
  wire  noWriteSideEffect = (isCSRRS | isCSRRC) & io_cfIn_instr[19:15] == 5'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 533:48]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~noWriteSideEffect; // @[src/main/scala/nutcore/backend/fu/CSR.scala 535:58]
  wire  _tvm_T_1 = priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:57]
  wire  tvm = mstatusStruct_tvm & priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:39]
  wire  _io_sfence_vma_invalid_T = priviledgeMode == 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:43]
  wire  _isIllegalTVM_T_1 = addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:42]
  wire  isIllegalTVM = tvm & wen & addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:34]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite | isIllegalTVM; // @[src/main/scala/nutcore/backend/fu/CSR.scala 544:57]
  wire  _canWriteCSR_T = ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:28]
  wire  _canWriteCSR_T_1 = wen & ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:25]
  wire  canWriteCSR = wen & ~isIllegalAccess & (addr != 12'h180 | satpLegalMode); // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:45]
  wire [63:0] _satp_T = wdata & 64'h8ffff000000fffff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _satp_T_2 = satp & 64'h70000ffffff00000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _satp_T_3 = _satp_T | _satp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mie_T = wdata & sieMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_1 = ~sieMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _mie_T_2 = mie & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mstatus_T = wdata & 64'hc0122; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_2 = mstatus & 64'hfffffffffff3fedd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_3 = _mstatus_T | _mstatus_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_mpp = _mstatus_T_3[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_3[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix = mstatus_mstatusOld_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_3[62:13],mstatus_mppFix,_mstatus_T_3[10:0]}
    ; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_6 = canWriteCSR & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mtvec_T = wdata & 64'hfffffffffffffffc; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mtvec_T_2 = mtvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtvec_T_3 = _mtvec_T | _mtvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mstatus_T_4 = wdata & 64'h80000000007e19aa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_6 = mstatus & 64'h7fffffffff81e655; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_7 = _mstatus_T_4 | _mstatus_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_1_mpp = _mstatus_T_7[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_1_fs = _mstatus_T_7[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix_1 = mstatus_mstatusOld_1_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_1_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew_1 = {mstatus_mstatusOld_1_fs == 2'h3,_mstatus_T_7[62:13],mstatus_mppFix_1,_mstatus_T_7[
    10:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_8 = canWriteCSR & addr == 12'h300 ? mstatus_mstatusNew_1 : _GEN_6; // @[src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_10 = canWriteCSR & addr == 12'h142 ? wdata : scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_65 = addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _medeleg_T = wdata & 64'hb3ff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'hffffffffffff4c00; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _stvec_T_2 = stvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _stvec_T_3 = _mtvec_T | _stvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _sepc_T = wdata & 64'hfffffffffffffffe; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _sepc_T_2 = sepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _sepc_T_3 = _sepc_T | _sepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_13 = canWriteCSR & addr == 12'h141 ? _sepc_T_3 : sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_14 = canWriteCSR & addr == 12'h342 ? wdata : mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mie_T_4 = wdata & 64'haaa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_6 = mie & 64'hfffffffffffff555; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_7 = _mie_T_4 | _mie_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_17 = canWriteCSR & addr == 12'h143 ? wdata : stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_79 = addr == 12'hb00; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_81 = addr == 12'hb02; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'hfffffffffffffddd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mepc_T_2 = mepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mepc_T_3 = _sepc_T | _mepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_21 = canWriteCSR & addr == 12'h341 ? _mepc_T_3 : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_22 = canWriteCSR & addr == 12'h343 ? wdata : mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _isIllegalAddr_illegalAddr_T_1 = _rdata_T_29 ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_3 = _rdata_T_30 ? 1'h0 : _isIllegalAddr_illegalAddr_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_5 = _rdata_T_31 ? 1'h0 : _isIllegalAddr_illegalAddr_T_3; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_7 = _rdata_T_32 ? 1'h0 : _isIllegalAddr_illegalAddr_T_5; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_9 = _rdata_T_33 ? 1'h0 : _isIllegalAddr_illegalAddr_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_11 = _rdata_T_34 ? 1'h0 : _isIllegalAddr_illegalAddr_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_13 = _rdata_T_35 ? 1'h0 : _isIllegalAddr_illegalAddr_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_15 = _rdata_T_36 ? 1'h0 : _isIllegalAddr_illegalAddr_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_17 = _rdata_T_37 ? 1'h0 : _isIllegalAddr_illegalAddr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_19 = _rdata_T_38 ? 1'h0 : _isIllegalAddr_illegalAddr_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_21 = _rdata_T_39 ? 1'h0 : _isIllegalAddr_illegalAddr_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_23 = _rdata_T_40 ? 1'h0 : _isIllegalAddr_illegalAddr_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_25 = _rdata_T_41 ? 1'h0 : _isIllegalAddr_illegalAddr_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_27 = _rdata_T_42 ? 1'h0 : _isIllegalAddr_illegalAddr_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_29 = _rdata_T_43 ? 1'h0 : _isIllegalAddr_illegalAddr_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_31 = _rdata_T_44 ? 1'h0 : _isIllegalAddr_illegalAddr_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_33 = _rdata_T_45 ? 1'h0 : _isIllegalAddr_illegalAddr_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_35 = _rdata_T_46 ? 1'h0 : _isIllegalAddr_illegalAddr_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_37 = _rdata_T_47 ? 1'h0 : _isIllegalAddr_illegalAddr_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_39 = _rdata_T_48 ? 1'h0 : _isIllegalAddr_illegalAddr_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_41 = _rdata_T_49 ? 1'h0 : _isIllegalAddr_illegalAddr_T_39; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_43 = _rdata_T_50 ? 1'h0 : _isIllegalAddr_illegalAddr_T_41; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_45 = _rdata_T_51 ? 1'h0 : _isIllegalAddr_illegalAddr_T_43; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_47 = _rdata_T_52 ? 1'h0 : _isIllegalAddr_illegalAddr_T_45; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_49 = _rdata_T_53 ? 1'h0 : _isIllegalAddr_illegalAddr_T_47; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_51 = _rdata_T_54 ? 1'h0 : _isIllegalAddr_illegalAddr_T_49; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_53 = _rdata_T_55 ? 1'h0 : _isIllegalAddr_illegalAddr_T_51; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_55 = _rdata_T_56 ? 1'h0 : _isIllegalAddr_illegalAddr_T_53; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  isIllegalAddr = _rdata_T_57 ? 1'h0 : _isIllegalAddr_illegalAddr_T_55; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  resetSatp = _isIllegalTVM_T_1 & wen & _canWriteCSR_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 552:42]
  wire  _io_isExit_T = addr == 12'h344; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:38]
  wire  _io_isExit_T_1 = addr == 12'h144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:56]
  wire  _io_isExit_T_9 = _canWriteCSR_T_1 | ~wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:30]
  wire  _io_isExit_T_10 = io_out_valid & (addr == 12'h344 | addr == 12'h144) & _wen_T_4 & _io_isExit_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:93]
  wire [63:0] _mipReg_T = wdata & 64'h77f; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mipReg_T_2 = mipReg & 64'hfffffffffffff880; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_3 = _mipReg_T | _mipReg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mipReg_T_6 = mipReg & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_7 = _mie_T | _mipReg_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _isEbreak_T_1 = io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:90]
  wire  isEcall = addr == 12'h0 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 569:88]
  wire  isMret = _T_65 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 570:88]
  wire  isSret = addr == 12'h102 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 571:88]
  wire  isUret = addr == 12'h2 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 572:88]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 639:63]
  wire  hasInstrAccessFault = io_cfIn_exceptionVec_1 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 640:67]
  wire  hasLoadPageFault = io_dmemMMU_loadPF | io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 641:43]
  wire  hasStorePageFault = io_dmemMMU_storePF | io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 642:45]
  wire  hasLoadAccessFault = io_dmemMMU_laf | io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:42]
  wire  hasStoreAccessFault = io_dmemMMU_saf | io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 644:43]
  wire [38:0] _imemExceptionAddr_T_1 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 651:42]
  wire  imemExceptionAddr_signBit = _imemExceptionAddr_T_1[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_2 = imemExceptionAddr_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_3 = {_imemExceptionAddr_T_2,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_6 = {25'h0,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_7 = vmEnable ? _imemExceptionAddr_T_3 : _imemExceptionAddr_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 651:12]
  wire  imemExceptionAddr_signBit_1 = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_8 = imemExceptionAddr_signBit_1 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_9 = {_imemExceptionAddr_T_8,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_10 = {25'h0,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_11 = vmEnable ? _imemExceptionAddr_T_9 : _imemExceptionAddr_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 652:12]
  wire [63:0] _imemExceptionAddr_T_12 = io_cfIn_crossBoundaryFault ? _imemExceptionAddr_T_7 : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 650:10]
  wire [63:0] imemExceptionAddr = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_12; // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:29]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 679:31]
  wire [11:0] _ideleg_T = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:41]
  wire [63:0] _GEN_87 = {{52'd0}, _ideleg_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:26]
  wire [63:0] ideleg = mideleg & _GEN_87; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:26]
  wire  _intrVecEnable_0_T_2 = priviledgeMode < 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:125]
  wire  _intrVecEnable_0_T_4 = priviledgeMode == 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 683:53]
  wire  _intrVecEnable_0_T_7 = priviledgeMode == 2'h3 & mstatusStruct_ie_m | _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 683:87]
  wire  intrVecEnable_0 = ideleg[0] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_1 = ideleg[1] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_2 = ideleg[2] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_3 = ideleg[3] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_4 = ideleg[4] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_5 = ideleg[5] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_6 = ideleg[6] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_7 = ideleg[7] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_8 = ideleg[8] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_9 = ideleg[9] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_10 = ideleg[10] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire  intrVecEnable_11 = ideleg[11] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 682:51]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _ideleg_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:27]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:65]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:65]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:49]
  wire [5:0] intrVecIDU_lo = {intrVec[5],1'h0,intrVec[3],1'h0,intrVec[1],1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 688:100]
  wire [11:0] intrVecIDU = {intrVec[11],1'h0,intrVec[9],1'h0,intrVec[7],1'h0,intrVecIDU_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 688:100]
  wire [2:0] _intrNO_T = io_cfIn_intrVec_5 ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [3:0] _intrNO_T_1 = io_cfIn_intrVec_9 ? 4'h9 : {{1'd0}, _intrNO_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [3:0] _intrNO_T_2 = io_cfIn_intrVec_1 ? 4'h1 : _intrNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [3:0] _intrNO_T_3 = io_cfIn_intrVec_7 ? 4'h7 : _intrNO_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [3:0] _intrNO_T_4 = io_cfIn_intrVec_11 ? 4'hb : _intrNO_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _intrNO_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:69]
  wire [5:0] _raiseIntr_T = {io_cfIn_intrVec_5,io_cfIn_intrVec_9,io_cfIn_intrVec_1,io_cfIn_intrVec_7,io_cfIn_intrVec_11,
    io_cfIn_intrVec_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:69]
  wire  raiseIntr = |_raiseIntr_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 694:76]
  wire  _illegalMret_T = io_in_valid & isMret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:33]
  wire  illegalMret = io_in_valid & isMret & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 697:43]
  wire  _illegalSret_T = io_in_valid & isSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:33]
  wire  illegalSret = io_in_valid & isSret & _intrVecEnable_0_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:43]
  wire  illegalSModeSret = _illegalSret_T & _tvm_T_1 & mstatusStruct_tsr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 699:76]
  wire  isIllegalPrivOp = illegalMret | illegalSret | illegalSModeSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 700:52]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[src/main/scala/nutcore/backend/fu/CSR.scala 705:46]
  wire  csrExceptionVec_11 = _intrVecEnable_0_T_4 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 706:70]
  wire  csrExceptionVec_9 = _tvm_T_1 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 707:70]
  wire  csrExceptionVec_8 = _io_sfence_vma_invalid_T & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 708:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen | isIllegalPrivOp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:79]
  wire [7:0] raiseExceptionVec_lo = {hasStoreAccessFault,1'h0,hasLoadAccessFault,1'h0,csrExceptionVec_3,
    csrExceptionVec_2,hasInstrAccessFault,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 716:43]
  wire [15:0] _raiseExceptionVec_T = {hasStorePageFault,1'h0,hasLoadPageFault,1'h0,csrExceptionVec_11,1'h0,
    csrExceptionVec_9,csrExceptionVec_8,raiseExceptionVec_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 716:43]
  wire [15:0] raiseExceptionVec = _raiseExceptionVec_T | _wen_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 716:50]
  wire  raiseException = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:42]
  wire [2:0] _exceptionNO_T_1 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [2:0] _exceptionNO_T_3 = raiseExceptionVec[7] ? 3'h7 : _exceptionNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_5 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _exceptionNO_T_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_7 = raiseExceptionVec[15] ? 4'hf : _exceptionNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_9 = raiseExceptionVec[4] ? 4'h4 : _exceptionNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_11 = raiseExceptionVec[6] ? 4'h6 : _exceptionNO_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_13 = raiseExceptionVec[8] ? 4'h8 : _exceptionNO_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_15 = raiseExceptionVec[9] ? 4'h9 : _exceptionNO_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_17 = raiseExceptionVec[11] ? 4'hb : _exceptionNO_T_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_19 = raiseExceptionVec[0] ? 4'h0 : _exceptionNO_T_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_21 = raiseExceptionVec[2] ? 4'h2 : _exceptionNO_T_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_23 = raiseExceptionVec[1] ? 4'h1 : _exceptionNO_T_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] _exceptionNO_T_25 = raiseExceptionVec[12] ? 4'hc : _exceptionNO_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _exceptionNO_T_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 718:74]
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:28]
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:53]
  wire [63:0] _GEN_88 = {{60'd0}, _causeNO_T_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:48]
  wire [63:0] causeNO = _causeNO_T | _GEN_88; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:48]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 724:58]
  wire [63:0] _redirectTarget_T_3 = _imemExceptionAddr_T_9 + 64'h4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 728:31]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 765:18]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 767:21]
  wire  delegS = _delegS_T_1[0] & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 767:36]
  wire [63:0] trapTarget = delegS ? stvec : mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 773:20]
  wire [63:0] _GEN_52 = _illegalSret_T & ~illegalSret & ~illegalSModeSret ? sepc : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 820:63 833:15]
  wire [63:0] retTarget = io_in_valid & isUret ? 64'h0 : _GEN_52; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:26 844:15]
  wire [63:0] _redirectTarget_T_4 = raiseExceptionIntr ? trapTarget : retTarget; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:8]
  wire [63:0] redirectTarget = resetSatp ? _redirectTarget_T_3 : _redirectTarget_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 727:27]
  reg [63:0] redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 740:36]
  wire  addrNotLegal_signBit = redirectTargetReg[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,redirectTargetReg[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _addrNotLegal_T_3 = redirectTargetReg != _addrNotLegal_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 742:23]
  wire  _addrNotLegal_T_5 = |redirectTargetReg[63:39]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 743:44]
  wire  addrNotLegal = vmEnable ? _addrNotLegal_T_3 : _addrNotLegal_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 741:25]
  reg  hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 745:31]
  reg  isIllegalXRET_REG; // @[src/main/scala/nutcore/backend/fu/CSR.scala 746:30]
  wire  isIllegalXRET = isIllegalXRET_REG & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/CSR.scala 746:50]
  wire  _T_162 = io_xretIsIllegal_ready & io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_27 = _T_162 ? 1'h0 : hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 749:38 750:20 745:31]
  wire  _GEN_28 = isIllegalXRET | _GEN_27; // @[src/main/scala/nutcore/backend/fu/CSR.scala 747:24 748:20]
  wire  isPageFault = hasInstrPageFault | hasLoadPageFault | hasStorePageFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 768:59]
  wire  isAddrMisAligned = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 769:48]
  wire  isAccessFault = hasInstrAccessFault | hasLoadAccessFault | hasStoreAccessFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 770:65]
  wire [63:0] _GEN_29 = delegS ? io_dmemExceptionAddr : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:21 779:15]
  wire [63:0] _GEN_30 = delegS ? _GEN_22 : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:21 781:15]
  wire [63:0] tval = hasInstrPageFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 786:21]
  wire [63:0] _GEN_31 = delegS ? tval : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:21 788:15]
  wire [63:0] _GEN_32 = delegS ? _GEN_22 : tval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:21 790:15]
  wire [63:0] tval_1 = hasInstrAccessFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 795:21]
  wire [63:0] _GEN_33 = delegS ? tval_1 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 796:21 797:15]
  wire [63:0] _GEN_34 = delegS ? _GEN_22 : tval_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 796:21 799:15]
  wire [63:0] _GEN_35 = isAccessFault ? _GEN_33 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 794:83]
  wire [63:0] _GEN_36 = isAccessFault ? _GEN_34 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/CSR.scala 794:83]
  wire [63:0] _GEN_37 = isPageFault ? _GEN_31 : _GEN_35; // @[src/main/scala/nutcore/backend/fu/CSR.scala 785:77]
  wire [63:0] _GEN_38 = isPageFault ? _GEN_32 : _GEN_36; // @[src/main/scala/nutcore/backend/fu/CSR.scala 785:77]
  wire [63:0] _GEN_39 = isAddrMisAligned ? _GEN_29 : _GEN_37; // @[src/main/scala/nutcore/backend/fu/CSR.scala 777:60]
  wire [63:0] _GEN_40 = isAddrMisAligned ? _GEN_30 : _GEN_38; // @[src/main/scala/nutcore/backend/fu/CSR.scala 777:60]
  wire [63:0] _GEN_41 = io_instrValid ? _GEN_39 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 776:24]
  wire [63:0] _GEN_42 = io_instrValid ? _GEN_40 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/CSR.scala 776:24]
  wire  mstatusOld_pie_m = mstatus[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 805:47]
  wire  mstatusNew_ie_u = mstatus[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_ie_h = mstatus[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_pie_u = mstatus[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_pie_s = mstatus[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_pie_h = mstatus[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_spp = mstatus[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [1:0] mstatusNew_hpp = mstatus[10:9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [1:0] mstatusNew_fs = mstatus[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [1:0] mstatusNew_xs = mstatus[16:15]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [8:0] mstatusNew_pad0 = mstatus[31:23]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [1:0] mstatusNew_uxl = mstatus[33:32]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [1:0] mstatusNew_sxl = mstatus[35:34]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire [26:0] mstatusNew_pad1 = mstatus[62:36]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_sd = mstatus[63]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 806:47]
  wire  mstatusNew_mprv = mstatusStruct_mpp != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 810:37 811:23 806:30]
  wire [5:0] mstatus_lo_lo = {mstatusNew_pie_s,mstatusNew_pie_u,mstatusOld_pie_m,mstatusNew_ie_h,mstatusStruct_ie_s,
    mstatusNew_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 815:27]
  wire [14:0] mstatus_lo = {mstatusNew_fs,2'h0,mstatusNew_hpp,mstatusNew_spp,1'h1,mstatusNew_pie_h,mstatus_lo_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 815:27]
  wire [6:0] mstatus_hi_lo = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_mprv,
    mstatusNew_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 815:27]
  wire [63:0] _mstatus_T_8 = {mstatusNew_sd,mstatusNew_pad1,mstatusNew_sxl,mstatusNew_uxl,mstatusNew_pad0,
    mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 815:27]
  wire [1:0] _GEN_44 = _illegalMret_T & ~illegalMret ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 804:42 809:20 262:31]
  wire [63:0] _GEN_45 = _illegalMret_T & ~illegalMret ? _mstatus_T_8 : _GEN_8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 804:42 815:13]
  wire [1:0] _priviledgeMode_T = {1'h0,mstatusNew_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 825:26]
  wire [1:0] _GEN_89 = {{1'd0}, mstatusNew_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 826:26]
  wire  mstatusNew_1_mprv = _GEN_89 != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 826:37 827:23 822:30]
  wire [5:0] mstatus_lo_lo_1 = {1'h1,mstatusNew_pie_u,mstatusStruct_ie_m,mstatusNew_ie_h,mstatusNew_pie_s,
    mstatusNew_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 831:27]
  wire [14:0] mstatus_lo_1 = {mstatusNew_fs,mstatusStruct_mpp,mstatusNew_hpp,1'h0,mstatusOld_pie_m,mstatusNew_pie_h,
    mstatus_lo_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 831:27]
  wire [6:0] mstatus_hi_lo_1 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_1_mprv
    ,mstatusNew_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 831:27]
  wire [63:0] _mstatus_T_9 = {mstatusNew_sd,mstatusNew_pad1,mstatusNew_sxl,mstatusNew_uxl,mstatusNew_pad0,
    mstatusStruct_tsr,mstatus_hi_lo_1,mstatus_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 831:27]
  wire [5:0] mstatus_lo_lo_2 = {mstatusNew_pie_s,1'h1,mstatusStruct_ie_m,mstatusNew_ie_h,mstatusStruct_ie_s,
    mstatusNew_pie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:27]
  wire [14:0] mstatus_lo_2 = {mstatusNew_fs,mstatusStruct_mpp,mstatusNew_hpp,mstatusNew_spp,mstatusOld_pie_m,
    mstatusNew_pie_h,mstatus_lo_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:27]
  wire [6:0] mstatus_hi_lo_2 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,
    mstatusStruct_mprv,mstatusNew_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:27]
  wire [63:0] _mstatus_T_10 = {mstatusNew_sd,mstatusNew_pad1,mstatusNew_sxl,mstatusNew_uxl,mstatusNew_pad0,
    mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:27]
  wire  tvalZeroWen = ~(isPageFault | isAddrMisAligned | isAccessFault) | raiseIntr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 847:73]
  wire [1:0] _GEN_60 = delegS ? priviledgeMode : {{1'd0}, mstatusNew_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 855:22 850:30]
  wire  mstatusNew_3_pie_s = delegS ? mstatusStruct_ie_s : mstatusNew_pie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 856:24 850:30]
  wire  mstatusNew_3_ie_s = delegS ? 1'h0 : mstatusStruct_ie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 857:23 850:30]
  wire [1:0] mstatusNew_3_mpp = delegS ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 850:30 867:22]
  wire  mstatusNew_3_pie_m = delegS ? mstatusOld_pie_m : mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 850:30 868:24]
  wire  mstatusNew_3_ie_m = delegS & mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19 850:30 869:23]
  wire [5:0] mstatus_lo_lo_3 = {mstatusNew_3_pie_s,mstatusNew_pie_u,mstatusNew_3_ie_m,mstatusNew_ie_h,mstatusNew_3_ie_s,
    mstatusNew_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 883:27]
  wire  mstatusNew_3_spp = _GEN_60[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 850:30]
  wire [14:0] mstatus_lo_3 = {mstatusNew_fs,mstatusNew_3_mpp,mstatusNew_hpp,mstatusNew_3_spp,mstatusNew_3_pie_m,
    mstatusNew_pie_h,mstatus_lo_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 883:27]
  wire [63:0] _mstatus_T_11 = {mstatusNew_sd,mstatusNew_pad1,mstatusNew_sxl,mstatusNew_uxl,mstatusNew_pad0,
    mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 883:27]
  wire  perfCntCondDisable_0 = wen & _T_79 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1017:42]
  wire  _WIRE = 1'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1008:{33,33}]
  wire [63:0] _perfCnts_0_T_5 = perfCnts_0 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:105]
  wire  perfCntCondDisable_2 = wen & _T_81 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1017:42]
  wire [63:0] _perfCnts_2_T_5 = perfCnts_2 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:105]
  wire [63:0] _perfCnts_2_T_7 = perfCnts_2 + 64'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1001:86]
  wire [3:0] _T_198 = raiseIntr & io_instrValid ? intrNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1094:43]
  wire [3:0] _T_200 = raiseException & io_instrValid ? exceptionNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1095:43]
  CSRDiffWrapper CSRDiffWrapper ( // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:29]
    .clock(CSRDiffWrapper_clock),
    .io_csrState_privilegeMode(CSRDiffWrapper_io_csrState_privilegeMode),
    .io_csrState_mstatus(CSRDiffWrapper_io_csrState_mstatus),
    .io_csrState_sstatus(CSRDiffWrapper_io_csrState_sstatus),
    .io_csrState_mepc(CSRDiffWrapper_io_csrState_mepc),
    .io_csrState_sepc(CSRDiffWrapper_io_csrState_sepc),
    .io_csrState_mtval(CSRDiffWrapper_io_csrState_mtval),
    .io_csrState_stval(CSRDiffWrapper_io_csrState_stval),
    .io_csrState_mtvec(CSRDiffWrapper_io_csrState_mtvec),
    .io_csrState_stvec(CSRDiffWrapper_io_csrState_stvec),
    .io_csrState_mcause(CSRDiffWrapper_io_csrState_mcause),
    .io_csrState_scause(CSRDiffWrapper_io_csrState_scause),
    .io_csrState_satp(CSRDiffWrapper_io_csrState_satp),
    .io_csrState_mip(CSRDiffWrapper_io_csrState_mip),
    .io_csrState_mie(CSRDiffWrapper_io_csrState_mie),
    .io_csrState_mscratch(CSRDiffWrapper_io_csrState_mscratch),
    .io_csrState_sscratch(CSRDiffWrapper_io_csrState_sscratch),
    .io_csrState_mideleg(CSRDiffWrapper_io_csrState_mideleg),
    .io_csrState_medeleg(CSRDiffWrapper_io_csrState_medeleg),
    .io_archEvent_valid(CSRDiffWrapper_io_archEvent_valid),
    .io_archEvent_interrupt(CSRDiffWrapper_io_archEvent_interrupt),
    .io_archEvent_exception(CSRDiffWrapper_io_archEvent_exception),
    .io_archEvent_exceptionPC(CSRDiffWrapper_io_archEvent_exceptionPC),
    .io_archEvent_exceptionInst(CSRDiffWrapper_io_archEvent_exceptionInst)
  );
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 887:16]
  assign io_out_bits = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_redirect_target = redirectTarget[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 736:22]
  assign io_redirect_valid = io_in_valid & _isEbreak_T_1 | raiseExceptionIntr | resetSatp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 734:80]
  assign io_xretIsIllegal_valid = hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 752:26]
  assign io_xretIsIllegal_bits = redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 753:25]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 610:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 611:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_wenFix = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:42]
  assign io_isPerfRead = io_out_valid & addr >= 12'hb00 & addr < 12'hb03; // @[src/main/scala/nutcore/backend/fu/CSR.scala 554:52]
  assign io_isExit = _io_isExit_T_10 & io_rfWenReal & rdata != 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:55]
  assign io_vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  assign io_sfence_vma_invalid = priviledgeMode == 2'h0 | tvm; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:53]
  assign io_wfi_invalid = priviledgeMode != 2'h3 & mstatusStruct_tw; // @[src/main/scala/nutcore/backend/fu/CSR.scala 546:46]
  assign lr_0 = lr;
  assign lrAddr_0 = lrAddr;
  assign satp_0 = satp;
  assign intrVecIDU_0 = intrVecIDU;
  assign CSRDiffWrapper_clock = clock;
  assign CSRDiffWrapper_io_csrState_privilegeMode = {{62'd0}, priviledgeMode}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1073:28]
  assign CSRDiffWrapper_io_csrState_mstatus = mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1074:22]
  assign CSRDiffWrapper_io_csrState_sstatus = mstatus & 64'h80000003000d8122; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1075:33]
  assign CSRDiffWrapper_io_csrState_mepc = mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1076:19]
  assign CSRDiffWrapper_io_csrState_sepc = sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1077:19]
  assign CSRDiffWrapper_io_csrState_mtval = mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1078:19]
  assign CSRDiffWrapper_io_csrState_stval = stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1079:19]
  assign CSRDiffWrapper_io_csrState_mtvec = mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1080:20]
  assign CSRDiffWrapper_io_csrState_stvec = stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1081:20]
  assign CSRDiffWrapper_io_csrState_mcause = mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1082:21]
  assign CSRDiffWrapper_io_csrState_scause = scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1083:21]
  assign CSRDiffWrapper_io_csrState_satp = satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1084:19]
  assign CSRDiffWrapper_io_csrState_mip = mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1085:18]
  assign CSRDiffWrapper_io_csrState_mie = mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1086:18]
  assign CSRDiffWrapper_io_csrState_mscratch = mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1087:23]
  assign CSRDiffWrapper_io_csrState_sscratch = sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1088:23]
  assign CSRDiffWrapper_io_csrState_mideleg = mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1089:22]
  assign CSRDiffWrapper_io_csrState_medeleg = medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1090:22]
  assign CSRDiffWrapper_io_archEvent_valid = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 724:58]
  assign CSRDiffWrapper_io_archEvent_interrupt = {{28'd0}, _T_198}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1094:37]
  assign CSRDiffWrapper_io_archEvent_exception = {{28'd0}, _T_200}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1095:37]
  assign CSRDiffWrapper_io_archEvent_exceptionPC = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 655:23]
  assign CSRDiffWrapper_io_archEvent_exceptionInst = io_cfIn_instr[31:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1097:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
      priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        priviledgeMode <= 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 858:22]
      end else begin
        priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 870:22]
      end
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:26]
      priviledgeMode <= 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:20]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 820:63]
      priviledgeMode <= _priviledgeMode_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 825:20]
    end else begin
      priviledgeMode <= _GEN_44;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
      mtvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end else if (canWriteCSR & addr == 12'h305) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mtvec <= _mtvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
      mcounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end else if (canWriteCSR & addr == 12'h306) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mcounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
      mcause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        mcause <= _GEN_14;
      end else begin
        mcause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 865:14]
      end
    end else begin
      mcause <= _GEN_14;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
      mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        mtval <= _GEN_42;
      end else if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 871:26]
        mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 872:15]
      end else begin
        mtval <= _GEN_42;
      end
    end else begin
      mtval <= _GEN_42;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
      mepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        mepc <= _GEN_21;
      end else if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 655:23]
        mepc <= io_illegalJump_bits;
      end else begin
        mepc <= _imemExceptionAddr_T_11;
      end
    end else begin
      mepc <= _GEN_21;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
      mie <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end else if (canWriteCSR & addr == 12'h304) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (canWriteCSR & addr == 12'h104) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
      mipReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end else if (_canWriteCSR_T_1 & _io_isExit_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_canWriteCSR_T_1 & _io_isExit_T) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
      mstatus <= 64'ha00001800; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      mstatus <= _mstatus_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 883:13]
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:26]
      mstatus <= _mstatus_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:13]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 820:63]
      mstatus <= _mstatus_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 831:13]
    end else begin
      mstatus <= _GEN_45;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
      medeleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end else if (canWriteCSR & addr == 12'h302) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      medeleg <= _medeleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
      mideleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end else if (canWriteCSR & addr == 12'h303) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mideleg <= _mideleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
      mscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end else if (canWriteCSR & addr == 12'h340) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
      stvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end else if (canWriteCSR & addr == 12'h105) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      stvec <= _stvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
      satp <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end else if (canWriteCSR & _isIllegalTVM_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      satp <= _satp_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
      sepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 655:23]
          sepc <= io_illegalJump_bits;
        end else begin
          sepc <= _imemExceptionAddr_T_11;
        end
      end else begin
        sepc <= _GEN_13;
      end
    end else begin
      sepc <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
      scause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        scause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 853:14]
      end else begin
        scause <= _GEN_10;
      end
    end else begin
      scause <= _GEN_10;
    end
    if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 848:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:19]
        if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 859:26]
          stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 860:15]
        end else begin
          stval <= _GEN_41;
        end
      end else begin
        stval <= _GEN_41;
      end
    end else begin
      stval <= _GEN_41;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
      sscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end else if (canWriteCSR & addr == 12'h140) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      sscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
      scounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end else if (canWriteCSR & addr == 12'h106) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      scounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 820:63]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 832:8]
    end else if (_illegalMret_T & ~illegalMret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 804:42]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 816:8]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lr <= set_lr_val; // @[src/main/scala/nutcore/backend/fu/CSR.scala 416:8]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
      lrAddr <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lrAddr <= set_lr_addr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 417:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (~perfCntCondDisable_0) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:96]
      perfCnts_0 <= _perfCnts_0_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:100]
    end else if (canWriteCSR & addr == 12'hb00) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (canWriteCSR & addr == 12'hb01) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 1001:35]
      perfCnts_2 <= _perfCnts_2_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1001:60]
    end else if (perfCntCondMinstret & ~perfCntCondDisable_2) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:96]
      perfCnts_2 <= _perfCnts_2_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 993:100]
    end else if (canWriteCSR & addr == 12'hb02) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (io_redirect_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 740:36]
      if (resetSatp) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 727:27]
        redirectTargetReg <= _redirectTarget_T_3;
      end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:8]
        if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 773:20]
          redirectTargetReg <= stvec;
        end else begin
          redirectTargetReg <= mtvec;
        end
      end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:26]
        redirectTargetReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 844:15]
      end else begin
        redirectTargetReg <= _GEN_52;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 745:31]
      hasIllegalXRET <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 745:31]
    end else begin
      hasIllegalXRET <= _GEN_28;
    end
    isIllegalXRET_REG <= io_redirect_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 746:30]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priviledgeMode = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcounteren = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtval = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mepc = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mipReg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  stvec = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  satp = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  sepc = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  scause = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  stval = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  sscratch = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  scounteren = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  lr = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  lrAddr = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  perfCnts_0 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  perfCnts_1 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  perfCnts_2 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  redirectTargetReg = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  hasIllegalXRET = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  isIllegalXRET_REG = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MOU(
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module DummyDPICWrapper_3(
  input         clock,
  input         io_bits_hasTrap, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_cycleCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_instrCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_code, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasTrap; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_instrCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasWFI; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_code; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestTrapEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_hasTrap(dpic_io_hasTrap),
    .io_cycleCnt(dpic_io_cycleCnt),
    .io_instrCnt(dpic_io_instrCnt),
    .io_hasWFI(dpic_io_hasWFI),
    .io_code(dpic_io_code),
    .io_pc(dpic_io_pc),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_hasTrap = io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_cycleCnt = io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instrCnt = io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_hasWFI = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_code = io_bits_code; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module EXUDiffWrapper(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [38:0] io_in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [63:0] io_in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_code; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] cycleCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
  wire [63:0] _cycleCnt_T_1 = cycleCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:24]
  reg [63:0] instrCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
  wire [63:0] _instrCnt_T_1 = instrCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:26]
  wire  nutcoretrap = io_in_bits_ctrl_isNutCoreTrap & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 194:66]
  DummyDPICWrapper_3 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .io_bits_hasTrap(difftest_module_io_bits_hasTrap),
    .io_bits_cycleCnt(difftest_module_io_bits_cycleCnt),
    .io_bits_instrCnt(difftest_module_io_bits_instrCnt),
    .io_bits_code(difftest_module_io_bits_code),
    .io_bits_pc(difftest_module_io_bits_pc)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_io_bits_hasTrap = nutcoretrap; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 199:21]
  assign difftest_module_io_bits_cycleCnt = cycleCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 202:21]
  assign difftest_module_io_bits_instrCnt = instrCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 203:21]
  assign difftest_module_io_bits_code = io_in_bits_data_src1[31:0]; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 200:21]
  assign difftest_module_io_bits_pc = {{25'd0}, io_in_bits_cf_pc}; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 201:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
      cycleCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
    end else begin
      cycleCnt <= _cycleCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
      instrCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
    end else if (perfCntCondMinstret) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 189:22]
      instrCnt <= _instrCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cycleCnt = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  instrCnt = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [3:0]  io__in_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [2:0]  io__in_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [6:0]  io__in_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [4:0]  io__in_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__out_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__out_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isExit, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__forward_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__sfence_vma_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__wfi_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12_0,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         falseWire,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_1,
  input         io_extra_msip,
  input         io_in_valid
);
  wire  alu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_offset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_iVmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_jumpIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isMissPredict; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_actualTarget; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_REG_0_fuOpType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [1:0] alu_REG_0_btbType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isRVC; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  lsu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [6:0] lsu_io__in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [31:0] lsu_io__instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbAF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scInflight_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_amoReq_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [55:0] lsu_dtlb_paddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_12_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scIsSuccess_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLrVal_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_DTLBFINISH; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lsuMMIO_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_13_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_setLrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  mdu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [6:0] mdu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  csr_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [6:0] csr_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_instrValid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_illegalJump_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wenFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isPerfRead; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_rfWenReal; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_meip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_lrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_satp_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_mtip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMultiCommit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr_val; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [11:0] csr_intrVecIDU_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_set_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_msip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  mou_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [6:0] mou_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushICache_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushTLB_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  diffMod_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [38:0] diffMod_io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [63:0] diffMod_io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  _fuValids_0_T_2 = ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:84]
  wire [15:0] _fuValids_0_T_4 = {2'h0,1'h0,io__in_bits_cf_exceptionVec_12,4'h0,4'h0,1'h0,io__in_bits_cf_exceptionVec_2,
    io__in_bits_cf_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:125]
  wire  _csr_io_cfIn_exceptionVec_13_T = lsu_io__in_valid & lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:62]
  wire  _csr_io_cfIn_exceptionVec_13_T_2 = io__in_bits_ctrl_fuOpType == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _csr_io_cfIn_exceptionVec_13_T_6 = io__in_bits_ctrl_fuOpType[5] & ~_csr_io_cfIn_exceptionVec_13_T_2 |
    io__in_bits_ctrl_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 64:69]
  wire  _csr_io_cfIn_exceptionVec_13_T_7 = ~_csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/fu/LSU.scala 65:40]
  wire  _T = alu_io_jumpIsIllegal_ready & alu_io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = csr_io_xretIsIllegal_ready & csr_io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_0 = csr_io_vmEnable | io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 104:48 73:15]
  wire  _GEN_1 = csr_io_vmEnable ? io__in_bits_cf_exceptionVec_1 : 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 73:15 106:50]
  wire  fuValids_1 = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4
    ); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  fuValids_3 = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 53:12 src/main/scala/nutcore/backend/seq/EXU.scala 58:26]
  wire  _hasException_T_1 = lsuTlbPF | lsu_io__dtlbAF | lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 123:50]
  wire  _hasException_T_3 = _hasException_T_1 | lsu_io__storeAddrMisaligned | lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 124:63]
  wire  hasException = _hasException_T_3 | lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 125:30]
  wire [38:0] _io_out_bits_decode_cf_redirect_T_target = csr_io_redirect_valid ? csr_io_redirect_target :
    alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_bits_decode_cf_redirect_T_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_valid_T_1 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_3 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _io_out_valid_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_4 = _io_out_valid_T_3 | csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 146:6]
  wire  _io_forward_wb_rfData_T = alu_io_out_ready & alu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _T_10 = _io_forward_wb_rfData_T & ~isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 163:43]
  wire  _T_12 = _io_forward_wb_rfData_T & isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 164:43]
  wire  _T_13 = lsu_io__out_ready & lsu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_14 = mdu_io_out_ready & mdu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = csr_io_out_ready & csr_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  ALU alu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    .io_iVmEnable(alu_io_iVmEnable),
    .io_jumpIsIllegal_ready(alu_io_jumpIsIllegal_ready),
    .io_jumpIsIllegal_valid(alu_io_jumpIsIllegal_valid),
    .io_jumpIsIllegal_bits(alu_io_jumpIsIllegal_bits),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC)
  );
  UnpipelinedLSU lsu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsu_io__isMMIO),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__dtlbAF(lsu_io__dtlbAF),
    .io__vaddr(lsu_io__vaddr),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .io__loadAccessFault(lsu_io__loadAccessFault),
    .io__storeAccessFault(lsu_io__storeAccessFault),
    .setLr_0(lsu_setLr_0),
    .lr_0(lsu_lr_0),
    .scInflight_0(lsu_scInflight_0),
    .amoReq_0(lsu_amoReq_0),
    .lr_addr(lsu_lr_addr),
    .dtlb_paddr(lsu_dtlb_paddr),
    ._T_12_0(lsu__T_12_0),
    .scIsSuccess_0(lsu_scIsSuccess_0),
    .setLrVal_0(lsu_setLrVal_0),
    .vmEnable(lsu_vmEnable),
    .DTLBFINISH(lsu_DTLBFINISH),
    .lsuMMIO_0(lsu_lsuMMIO_0),
    ._T_13_1(lsu__T_13_1),
    .setLrAddr_0(lsu_setLrAddr_0)
  );
  MDU mdu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_5(csr_io_cfIn_exceptionVec_5),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_7(csr_io_cfIn_exceptionVec_7),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_exceptionVec_13(csr_io_cfIn_exceptionVec_13),
    .io_cfIn_exceptionVec_15(csr_io_cfIn_exceptionVec_15),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossBoundaryFault(csr_io_cfIn_crossBoundaryFault),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_illegalJump_valid(csr_io_illegalJump_valid),
    .io_illegalJump_bits(csr_io_illegalJump_bits),
    .io_dmemExceptionAddr(csr_io_dmemExceptionAddr),
    .io_xretIsIllegal_ready(csr_io_xretIsIllegal_ready),
    .io_xretIsIllegal_valid(csr_io_xretIsIllegal_valid),
    .io_xretIsIllegal_bits(csr_io_xretIsIllegal_bits),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_laf(csr_io_dmemMMU_laf),
    .io_dmemMMU_saf(csr_io_dmemMMU_saf),
    .io_wenFix(csr_io_wenFix),
    .io_isPerfRead(csr_io_isPerfRead),
    .io_isExit(csr_io_isExit),
    .io_vmEnable(csr_io_vmEnable),
    .io_rfWenReal(csr_io_rfWenReal),
    .io_sfence_vma_invalid(csr_io_sfence_vma_invalid),
    .io_wfi_invalid(csr_io_wfi_invalid),
    .set_lr(csr_set_lr),
    .lr_0(csr_lr_0),
    .meip_0(csr_meip_0),
    .lrAddr_0(csr_lrAddr_0),
    .satp_0(csr_satp_0),
    .mtip_0(csr_mtip_0),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .intrVecIDU_0(csr_intrVecIDU_0),
    .set_lr_addr(csr_set_lr_addr),
    .msip_0(csr_msip_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret)
  );
  MOU mou ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  EXUDiffWrapper diffMod ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
    .clock(diffMod_clock),
    .reset(diffMod_reset),
    .io_in_valid(diffMod_io_in_valid),
    .io_in_bits_cf_pc(diffMod_io_in_bits_cf_pc),
    .io_in_bits_ctrl_isNutCoreTrap(diffMod_io_in_bits_ctrl_isNutCoreTrap),
    .io_in_bits_data_src1(diffMod_io_in_bits_data_src1),
    .io_flush(diffMod_io_flush),
    .perfCntCondMinstret(diffMod_perfCntCondMinstret)
  );
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 154:31]
  assign io__out_valid = io__in_valid & _io_out_valid_T_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 143:31]
  assign io__out_bits_decode_cf_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 131:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 130:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target :
    _io_out_bits_decode_cf_redirect_T_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid :
    _io_out_bits_decode_cf_redirect_T_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 128:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~hasException | ~fuValids_1) & ~(csr_io_wenFix &
    fuValids_3); // @[src/main/scala/nutcore/backend/seq/EXU.scala 126:68]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 127:14]
  assign io__out_bits_isMMIO = io__out_bits_decode_ctrl_rfWen & csr_io_isPerfRead | lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:61 112:24 62:22]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 148:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 149:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 151:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 150:35]
  assign io__out_bits_isExit = csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 134:22]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__forward_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 156:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/EXU.scala 157:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 158:24]
  assign io__forward_wb_rfData = _io_forward_wb_rfData_T ? alu_io_out_bits : lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 159:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 160:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 89:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__sfence_vma_invalid = csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 86:25]
  assign io__wfi_invalid = csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 87:18]
  assign lr = csr_lr_0;
  assign scInflight = lsu_scInflight_0;
  assign REG_valid = alu_REG_0_valid;
  assign REG_pc = alu_REG_0_pc;
  assign REG_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_actualTarget = alu_REG_0_actualTarget;
  assign REG_fuOpType = alu_REG_0_fuOpType;
  assign REG_btbType = alu_REG_0_btbType;
  assign REG_isRVC = alu_REG_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign lrAddr = csr_lrAddr_0;
  assign satp = csr_satp_0;
  assign flushICache = mou_flushICache_0;
  assign flushTLB = mou_flushTLB_0;
  assign intrVecIDU = csr_intrVecIDU_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 85:15]
  assign alu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 53:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/EXU.scala 52:17]
  assign alu_io_iVmEnable = csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 90:20]
  assign alu_io_jumpIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:45]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 51:21]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 52:21]
  assign lsu_io__out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 64:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/EXU.scala 61:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_lr_0 = lr;
  assign lsu_lr_addr = lrAddr;
  assign lsu_dtlb_paddr = paddr;
  assign lsu__T_12_0 = _T_12_0;
  assign lsu_scIsSuccess_0 = scIsSuccess;
  assign lsu_vmEnable = vmEnable;
  assign lsu_DTLBFINISH = tlbFinish;
  assign lsu_lsuMMIO_0 = ismmio;
  assign lsu__T_13_1 = _T_13_1;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4)
    ; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/CSR.scala 207:15]
  assign csr_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 84:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_1 = _T | _T_1 ? _GEN_1 : io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 74:48]
  assign csr_io_cfIn_exceptionVec_5 = lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 76:45]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:49]
  assign csr_io_cfIn_exceptionVec_7 = lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 77:46]
  assign csr_io_cfIn_exceptionVec_12 = _T | _T_1 ? _GEN_0 : io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_13 = lsu_io__in_valid & lsu_io__dtlbPF & _csr_io_cfIn_exceptionVec_13_T_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:79]
  assign csr_io_cfIn_exceptionVec_15 = _csr_io_cfIn_exceptionVec_13_T & _csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 79:80]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_crossBoundaryFault = io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_instrValid = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:36]
  assign csr_io_illegalJump_valid = alu_io_jumpIsIllegal_valid | csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 95:60]
  assign csr_io_illegalJump_bits = alu_io_jumpIsIllegal_valid ? alu_io_jumpIsIllegal_bits : csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 96:36]
  assign csr_io_dmemExceptionAddr = lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:28]
  assign csr_io_xretIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 98:45]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_laf = io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_saf = io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_rfWenReal = io__in_bits_ctrl_rfWen & io__in_bits_ctrl_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 85:45]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_msip_0 = io_extra_msip;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign mou_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 118:15]
  assign diffMod_clock = clock;
  assign diffMod_reset = reset;
  assign diffMod_io_in_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 171:25]
  assign diffMod_io_in_bits_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_ctrl_isNutCoreTrap = io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_data_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_flush = io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 173:22]
  assign diffMod_perfCntCondMinstret = io_in_valid;
endmodule
module DummyDPICWrapper_4(
  input         clock,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_skip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_isRVC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_rfwen, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_wpdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_wdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_instr, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_special // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_skip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isRVC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_rfwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_fpwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_vecwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_wpdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_wdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_instr; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [9:0] dpic_io_robIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_lqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_sqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isLoad; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isStore; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_nFused; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_special; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestInstrCommit dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_skip(dpic_io_skip),
    .io_isRVC(dpic_io_isRVC),
    .io_rfwen(dpic_io_rfwen),
    .io_fpwen(dpic_io_fpwen),
    .io_vecwen(dpic_io_vecwen),
    .io_wpdest(dpic_io_wpdest),
    .io_wdest(dpic_io_wdest),
    .io_pc(dpic_io_pc),
    .io_instr(dpic_io_instr),
    .io_robIdx(dpic_io_robIdx),
    .io_lqIdx(dpic_io_lqIdx),
    .io_sqIdx(dpic_io_sqIdx),
    .io_isLoad(dpic_io_isLoad),
    .io_isStore(dpic_io_isStore),
    .io_nFused(dpic_io_nFused),
    .io_special(dpic_io_special),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_skip = io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isRVC = io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_rfwen = io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_fpwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_vecwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wpdest = io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wdest = io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instr = io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_robIdx = 10'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_lqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isLoad = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isStore = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_nFused = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_special = io_bits_special; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DiffInstrCommitWrapper(
  input         clock,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_skip, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_isRVC, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_rfwen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [4:0]  io_wpdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [7:0]  io_wdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [63:0] io_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [31:0] io_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [7:0]  io_special // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_special; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [4:0] difftest_REG_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [7:0] difftest_REG_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [63:0] difftest_REG_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [31:0] difftest_REG_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [7:0] difftest_REG_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  DummyDPICWrapper_4 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_skip(difftest_module_io_bits_skip),
    .io_bits_isRVC(difftest_module_io_bits_isRVC),
    .io_bits_rfwen(difftest_module_io_bits_rfwen),
    .io_bits_wpdest(difftest_module_io_bits_wpdest),
    .io_bits_wdest(difftest_module_io_bits_wdest),
    .io_bits_pc(difftest_module_io_bits_pc),
    .io_bits_instr(difftest_module_io_bits_instr),
    .io_bits_special(difftest_module_io_bits_special)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_skip = difftest_REG_skip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_isRVC = difftest_REG_isRVC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_rfwen = difftest_REG_rfwen; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_wpdest = difftest_REG_wpdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_wdest = difftest_REG_wdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_pc = difftest_REG_pc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_instr = difftest_REG_instr; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_special = difftest_REG_special; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_skip <= io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_isRVC <= io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_rfwen <= io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_wpdest <= io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_wdest <= io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_pc <= io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_instr <= io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_special <= io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_skip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  difftest_REG_isRVC = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  difftest_REG_rfwen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  difftest_REG_wpdest = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  difftest_REG_wdest = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_pc = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  difftest_REG_instr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  difftest_REG_special = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_5(
  input         clock,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_address, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_address; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestIntWriteback dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_address(dpic_io_address),
    .io_data(dpic_io_data),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_address = io_bits_address; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DiffIntWbWrapper(
  input         clock,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
  input  [4:0]  io_address, // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
  input  [63:0] io_data // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_address; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  reg [4:0] difftest_REG_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  reg [63:0] difftest_REG_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  DummyDPICWrapper_5 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_address(difftest_module_io_bits_address),
    .io_bits_data(difftest_module_io_bits_data)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_address = difftest_REG_address; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_data = difftest_REG_data; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
    difftest_REG_address <= io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
    difftest_REG_data <= io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_address = _RAND_1[4:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_data = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [2:0]  io__in_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isExit, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__wb_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [4:0]  io__wb_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [63:0] io__wb_rfData, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [38:0] io__redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        falseWire_0,
  output        io_in_valid
);
  wire  DiffInstrCommitWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [4:0] DiffInstrCommitWrapper_io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [7:0] DiffInstrCommitWrapper_io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [63:0] DiffInstrCommitWrapper_io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [31:0] DiffInstrCommitWrapper_io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [7:0] DiffInstrCommitWrapper_io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffIntWbWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire  DiffIntWbWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [4:0] DiffIntWbWrapper_io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [63:0] DiffIntWbWrapper_io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  signBit = io__in_bits_decode_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _T = signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire  _T_4 = io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 89:51]
  wire [1:0] _T_6 = {io__in_bits_isExit,1'h0}; // @[difftest/src/main/scala/Bundles.scala 81:19]
  wire  falseWire = 1'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 62:{27,27}]
  DiffInstrCommitWrapper DiffInstrCommitWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
    .clock(DiffInstrCommitWrapper_clock),
    .io_valid(DiffInstrCommitWrapper_io_valid),
    .io_skip(DiffInstrCommitWrapper_io_skip),
    .io_isRVC(DiffInstrCommitWrapper_io_isRVC),
    .io_rfwen(DiffInstrCommitWrapper_io_rfwen),
    .io_wpdest(DiffInstrCommitWrapper_io_wpdest),
    .io_wdest(DiffInstrCommitWrapper_io_wdest),
    .io_pc(DiffInstrCommitWrapper_io_pc),
    .io_instr(DiffInstrCommitWrapper_io_instr),
    .io_special(DiffInstrCommitWrapper_io_special)
  );
  DiffIntWbWrapper DiffIntWbWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
    .clock(DiffIntWbWrapper_clock),
    .io_valid(DiffIntWbWrapper_io_valid),
    .io_address(DiffIntWbWrapper_io_address),
    .io_data(DiffIntWbWrapper_io_data)
  );
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 35:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 36:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/seq/WBU.scala 41:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 42:60]
  assign falseWire_0 = falseWire;
  assign io_in_valid = io__in_valid;
  assign DiffInstrCommitWrapper_clock = clock;
  assign DiffInstrCommitWrapper_io_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 84:20]
  assign DiffInstrCommitWrapper_io_skip = io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/seq/WBU.scala 87:19]
  assign DiffInstrCommitWrapper_io_isRVC = io__in_bits_decode_cf_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 88:56]
  assign DiffInstrCommitWrapper_io_rfwen = io__wb_rfWen & io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 89:35]
  assign DiffInstrCommitWrapper_io_wpdest = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 91:21]
  assign DiffInstrCommitWrapper_io_wdest = {{3'd0}, io__wb_rfDest}; // @[src/main/scala/nutcore/backend/seq/WBU.scala 90:20]
  assign DiffInstrCommitWrapper_io_pc = {_T,io__in_bits_decode_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  assign DiffInstrCommitWrapper_io_instr = io__in_bits_decode_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/WBU.scala 86:20]
  assign DiffInstrCommitWrapper_io_special = {{6'd0}, _T_6}; // @[difftest/src/main/scala/Bundles.scala 81:13]
  assign DiffIntWbWrapper_clock = clock;
  assign DiffIntWbWrapper_io_valid = io__wb_rfWen & _T_4; // @[src/main/scala/nutcore/backend/seq/WBU.scala 116:35]
  assign DiffIntWbWrapper_io_address = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 117:22]
  assign DiffIntWbWrapper_io_data = io__wb_rfData; // @[src/main/scala/nutcore/backend/seq/WBU.scala 118:19]
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_0,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_lr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_meip_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scInflight; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isMissPredict; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_actualTarget; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_REG_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_REG_btbType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isRVC; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_amoReq; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_lrAddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [55:0] exu_paddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_satp; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_12_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scIsSuccess; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_mtip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushICache; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_falseWire; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_vmEnable; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushTLB; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [11:0] exu_intrVecIDU; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_tlbFinish; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_ismmio; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_13_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_msip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_falseWire_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io__in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _T_4 = exu_io__out_valid; // @[src/main/scala/utils/Pipeline.scala 26:22]
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  ISU isu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(isu_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(isu_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(isu_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(isu_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossBoundaryFault(exu_io__in_bits_cf_crossBoundaryFault),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_isNutCoreTrap(exu_io__in_bits_ctrl_isNutCoreTrap),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_instr(exu_io__out_bits_decode_cf_instr),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_isMMIO(exu_io__out_bits_isMMIO),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__out_bits_isExit(exu_io__out_bits_isExit),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_laf(exu_io__memMMU_dmem_laf),
    .io__memMMU_dmem_saf(exu_io__memMMU_dmem_saf),
    .io__sfence_vma_invalid(exu_io__sfence_vma_invalid),
    .io__wfi_invalid(exu_io__wfi_invalid),
    .lr(exu_lr),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .scInflight(exu_scInflight),
    .REG_valid(exu_REG_valid),
    .REG_pc(exu_REG_pc),
    .REG_isMissPredict(exu_REG_isMissPredict),
    .REG_actualTarget(exu_REG_actualTarget),
    .REG_fuOpType(exu_REG_fuOpType),
    .REG_btbType(exu_REG_btbType),
    .REG_isRVC(exu_REG_isRVC),
    .amoReq(exu_amoReq),
    .lrAddr(exu_lrAddr),
    .paddr(exu_paddr),
    .satp(exu_satp),
    ._T_12_0(exu__T_12_0),
    .scIsSuccess(exu_scIsSuccess),
    .io_extra_mtip(exu_io_extra_mtip),
    .flushICache(exu_flushICache),
    .falseWire(exu_falseWire),
    .vmEnable(exu_vmEnable),
    .flushTLB(exu_flushTLB),
    .intrVecIDU(exu_intrVecIDU),
    .tlbFinish(exu_tlbFinish),
    .ismmio(exu_ismmio),
    ._T_13_1(exu__T_13_1),
    .io_extra_msip(exu_io_extra_msip),
    .io_in_valid(exu_io_in_valid)
  );
  WBU wbu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
    .clock(wbu_clock),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_isMMIO(wbu_io__in_bits_isMMIO),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_isExit(wbu_io__in_bits_isExit),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .falseWire_0(wbu_falseWire_0),
    .io_in_valid(wbu_io_in_valid)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 698:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_sfence_vma_invalid = exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:25]
  assign io_wfi_invalid = exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign lr = exu_lr;
  assign scInflight = exu_scInflight;
  assign REG_valid = exu_REG_valid;
  assign REG_pc = exu_REG_pc;
  assign REG_isMissPredict = exu_REG_isMissPredict;
  assign REG_actualTarget = exu_REG_actualTarget;
  assign REG_fuOpType = exu_REG_fuOpType;
  assign REG_btbType = exu_REG_btbType;
  assign REG_isRVC = exu_REG_isRVC;
  assign amoReq = exu_amoReq;
  assign lrAddr = exu_lrAddr;
  assign satp = exu_satp;
  assign flushICache = exu_flushICache;
  assign flushTLB = exu_flushTLB;
  assign intrVecIDU = exu_intrVecIDU;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_flush = io_flush[0]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 688:27]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossBoundaryFault = exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_isNutCoreTrap = exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 689:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_laf = io_memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_saf = io_memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_paddr = paddr;
  assign exu__T_12_0 = _T_12;
  assign exu_scIsSuccess = scIsSuccess;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_falseWire = wbu_falseWire_0;
  assign exu_vmEnable = vmEnable;
  assign exu_tlbFinish = tlbFinish;
  assign exu_ismmio = ismmio;
  assign exu__T_13_1 = _T_13_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign wbu_clock = clock;
  assign wbu_io__in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isMMIO = wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isExit = wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_instr <= isu_io_out_bits_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pc <= isu_io_out_bits_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_crossBoundaryFault <= isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_isNutCoreTrap <= isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src1 <= isu_io_out_bits_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src2 <= isu_io_out_bits_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_imm <= isu_io_out_bits_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _T_4;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_instr <= exu_io__out_bits_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isMMIO <= exu_io__out_bits_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_0 <= exu_io__out_bits_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_1 <= exu_io__out_bits_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_2 <= exu_io__out_bits_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_3 <= exu_io__out_bits_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isExit <= exu_io__out_bits_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_crossBoundaryFault = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_isNutCoreTrap = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  valid_1 = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc = _RAND_25[38:0];
  _RAND_26 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  wbu_io_in_bits_r_isMMIO = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3 = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  wbu_io_in_bits_r_isExit = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_0_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_1_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
  end
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_2_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_2_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_2_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [1:0]  io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire [31:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [31:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_5; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_9 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_10 = 2'h2 == io_chosen ? 3'h3 : _GEN_9; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_17 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_18 = 2'h2 == io_chosen ? 8'hff : _GEN_17; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_21; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire [1:0] io_chosen_choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire  _T_4 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = 2'h3 == io_chosen ? 1'h0 : _GEN_2; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? 32'h0 : _GEN_6; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? 3'h0 : _GEN_10; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? 4'h0 : _GEN_14; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? 8'h0 : _GEN_18; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? 64'h0 : _GEN_22; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_0_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [1:0] inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_13 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  LockingArbiter_1 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
  end
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [86:0]  io_in_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [86:0]  io_out_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:20]
  wire  hitExec = hitCheck & ~hitADCheck & hitFlag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:41]
  wire  hitinstrPF = ~hitExec & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 290:52]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
  wire  isFlush = needFlush | io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 314:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26 315:{40,52}]
  wire  _GEN_4 = _alreadyOutFire_T & needFlush ? 1'h0 : _GEN_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 316:{37,49}]
  reg  missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  _T_5 = ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 324:13]
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = raddrCancel ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:29]
  wire  _GEN_16 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire [2:0] _GEN_17 = _T_10 ? 3'h2 : _GEN_15; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38 342:15]
  wire  _GEN_18 = _T_10 ? missPTEAF : _GEN_16; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26 341:38]
  wire  _GEN_20 = isFlush ? 1'h0 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22 340:19]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire [2:0] _GEN_22 = is_reserved ? 3'h4 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 372:21]
  wire  _GEN_23 = is_reserved | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 371:32 374:25]
  wire [2:0] _GEN_24 = ~missflag_v | ~missflag_r & missflag_w ? 3'h4 : _GEN_22; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:43]
  wire  _GEN_25 = ~missflag_v | ~missflag_r & missflag_w | _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 358:45]
  wire [55:0] _GEN_26 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_117 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_117; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:24]
  wire  permExec = permCheck & ~_T_21 & ~permAD & ~misaligned & missflag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:75]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = 8'h40 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | 64'h40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire  _GEN_27 = ~permExec | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 396:{30,40}]
  wire  _GEN_29 = ~permExec ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 396:30 304:32 399:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_30 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_31 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire  _GEN_32 = level != 2'h0 ? _GEN_27 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 383:36]
  wire [2:0] _GEN_33 = level != 2'h0 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_34 = level != 2'h0 & _GEN_29; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_35 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_43 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_51 = isFlush ? 18'h3ffff : _GEN_43; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 302:26]
  wire [17:0] _GEN_60 = _T_12 ? _GEN_51 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_87 = 3'h2 == state ? _GEN_60 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_100 = 3'h1 == state ? 18'h3ffff : _GEN_87; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_100; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_36 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_37 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_24 : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_38 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_25 : _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_39 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_26 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_40 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_30; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_41 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_31; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_42 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_44 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [2:0] _GEN_45 = isFlush ? 3'h0 : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 353:17]
  wire  _GEN_46 = isFlush ? missIPF : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 352:24]
  wire [55:0] _GEN_47 = isFlush ? raddr : _GEN_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 352:24]
  wire [7:0] _GEN_48 = isFlush ? 8'h0 : _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 305:32]
  wire [63:0] _GEN_49 = isFlush ? memRespStore : _GEN_41; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 301:25]
  wire  _GEN_50 = isFlush ? 1'h0 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 304:32]
  wire [17:0] _GEN_52 = isFlush ? missMaskStore : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 303:26]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_53 = _T_12 ? _GEN_45 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_54 = _T_12 ? _GEN_20 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
  wire  _GEN_55 = _T_12 ? _GEN_46 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 351:33]
  wire  _GEN_59 = _T_12 & _GEN_50; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_62 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire [2:0] _GEN_63 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire [2:0] _GEN_64 = isFlush ? 3'h0 : _GEN_63; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 420:22 421:15]
  wire [2:0] _GEN_65 = io_isFinish | io_flush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_66 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 428:15 318:24]
  wire  _GEN_67 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_68 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire [2:0] _GEN_69 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_70 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_71 = 3'h4 == state ? _GEN_65 : _GEN_69; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_72 = 3'h4 == state ? _GEN_66 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_73 = 3'h4 == state ? _GEN_67 : _GEN_70; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_74 = 3'h4 == state ? _GEN_68 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_75 = 3'h3 == state ? _GEN_64 : _GEN_71; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_76 = 3'h3 == state ? _GEN_20 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_77 = 3'h3 == state ? missIPF : _GEN_72; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_78 = 3'h3 == state ? missPTEAF : _GEN_73; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_79 = 3'h3 == state ? _GEN_2 : _GEN_74; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_99 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_59; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_99; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _io_mem_req_valid_T_3 = ~isFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:76]
  wire  _T_34 = missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:50]
  wire  _T_35 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire  out_req_valid = io_in_valid & (hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _instrAF_T_2 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _instrAF_T_5 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _instrAF_T_6 = {_instrAF_T_5,_instrAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _instrAF_T_7 = |_instrAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  hasException = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  assign io_in_ready = io_out_ready & _T_35 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:75]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_user = io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 500:16]
  assign io_iaf = out_req_valid & (~_instrAF_T_7 | missPTEAF); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 486:30]
  assign io_isFinish = _alreadyOutFire_T | hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:32]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 339:15]
      end else begin
        state <= _GEN_17;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_53;
    end else begin
      state <= _GEN_75;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_62;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_49;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_52;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_47;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_79;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 332:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 340:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      needFlush <= _GEN_54;
    end else begin
      needFlush <= _GEN_76;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
      missIPF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          missIPF <= _GEN_55;
        end else begin
          missIPF <= _GEN_77;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(isFlush)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
          missPTEAF <= _GEN_18;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_78;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else begin
      REG <= missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_51;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_48;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= _T_34 & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  memRespStore = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  missMaskStore = _RAND_4[17:0];
  _RAND_5 = {2{`RANDOM}};
  raddr = _RAND_5[55:0];
  _RAND_6 = {1{`RANDOM}};
  alreadyOutFire = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  needFlush = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  missIPF = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missPTEAF = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_2 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  REG_3 = _RAND_12[26:0];
  _RAND_13 = {1{`RANDOM}};
  REG_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  REG_5 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  REG_6 = _RAND_15[7:0];
  _RAND_16 = {2{`RANDOM}};
  REG_7 = _RAND_16[43:0];
  _RAND_17 = {2{`RANDOM}};
  REG_8 = _RAND_17[55:0];
  _RAND_18 = {1{`RANDOM}};
  blockRefill = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_out_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_out_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  wire  _reqIsLegalInstr_T_2 = io_in_req_bits_addr >= 39'h40000000 & io_in_req_bits_addr < 39'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _reqIsLegalInstr_T_5 = io_in_req_bits_addr >= 39'h80000000 & io_in_req_bits_addr < 39'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _reqIsLegalInstr_T_6 = {_reqIsLegalInstr_T_5,_reqIsLegalInstr_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _reqIsLegalInstr_T_7 = |_reqIsLegalInstr_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  reqIsLegalInstr = vmEnable | _reqIsLegalInstr_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 119:34]
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
  wire  _lastReqAddr_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _lastReqAddr_T_2 = _lastReqAddr_T & ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:67]
  reg [38:0] lastReqAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
  wire  _T_1 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_5 = _T_1 & io_in_resp_bits_user[38:0] == lastReqAddr ? 1'h0 : hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 127:96 128:19 120:28]
  wire  _GEN_6 = _lastReqAddr_T | _GEN_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 125:33 126:19]
  reg  hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
  wire  _hasIllegalInflight_T = ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:27]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  _GEN_10 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _GEN_11 = mdUpdate & vmEnable | _GEN_10; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [86:0] tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  _GEN_19 = io_in_req_valid & _hasIllegalInflight_T ? ~hasInflight : io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:23 158:50 159:25]
  wire  _GEN_20 = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 170:23]
  wire  _GEN_21 = ~vmEnable ? io_in_req_valid & reqIsLegalInstr : tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 156:24 170:23]
  reg [86:0] userBits; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
  EmbeddedTLBExec tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_ipf(tlbExec_io_ipf),
    .io_iaf(tlbExec_io_iaf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBMD mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? _GEN_19 : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19]
  assign io_in_resp_valid = hasIllegalInflight & io_iaf | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 202:24]
  assign io_in_resp_bits_rdata = hasIllegalInflight & io_iaf ? 64'h0 : io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 203:29]
  assign io_in_resp_bits_user = hasIllegalInflight & io_iaf ? userBits : io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 206:34]
  assign io_out_req_valid = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_21; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 191:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 170:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 167:32 170:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_iaf = vmEnable ? tlbExec_io_iaf : hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 212:16]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_user = tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_20; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 190:28]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_flush = io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:20]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 123:21]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 124:19]
    end else begin
      hasInflight <= _GEN_6;
    end
    if (_lastReqAddr_T & ~io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
      lastReqAddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
    end else if (_T_1 | io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 132:38]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 133:24]
    end else if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 134:44]
      hasIllegalInflight <= ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:24]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:20]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:28]
    end else begin
      valid <= _GEN_11;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_user <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
      userBits <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  hasInflight = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  hasIllegalInflight = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_8[38:0];
  _RAND_9 = {3{`RANDOM}};
  tlbExec_io_in_bits_r_user = _RAND_9[86:0];
  _RAND_10 = {3{`RANDOM}};
  userBits = _RAND_10[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PTERequestFilter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_u // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  isLegal = |(io_in_req_bits_addr >= 32'h80000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasInflight_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [7:0] _io_in_resp_bits_rdata_T = {3'h7,io_u,4'hf}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 570:33]
  assign io_in_req_ready = isLegal ? io_out_req_ready : ~hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 562:25]
  assign io_in_resp_valid = ~io_out_resp_valid & hasInflight | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 567:22]
  assign io_in_resp_bits_rdata = ~io_out_resp_valid & hasInflight ? {{56'd0}, _io_in_resp_bits_rdata_T} :
    io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 570:27]
  assign io_out_req_valid = io_in_req_valid & isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 561:39]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end else if (~io_out_resp_valid & hasInflight) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:44]
      hasInflight <= 1'h0;
    end else begin
      hasInflight <= _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasInflight = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_fake(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [95:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  reg  needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  _GEN_1 = io_flush[0] & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26 567:{44,56}]
  wire  _alreadyOutFire_T = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire [2:0] _GEN_9 = _alreadyOutFire_T | needFlush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [86:0] memuser; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5 & ~needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 601:47]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_in_resp_bits_user = memuser; // @[src/main/scala/nutcore/mem/Cache.scala 612:93]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T & ~io_flush[0]) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    end else if (state == 3'h0 & needFlush) begin // @[src/main/scala/nutcore/mem/Cache.scala 568:40]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 568:52]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
      memuser <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  needFlush = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alreadyOutFire = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reqaddr = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  mmiordata = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  memrdata = _RAND_6[63:0];
  _RAND_7 = {3{`RANDOM}};
  memuser = _RAND_7[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [2:0]   io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [3:0]   io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [7:0]   io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [2:0]   io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [7:0]   io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_out_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          lr_0,
  input          scInflight_0,
  input          ISAMO,
  input  [63:0]  lr_addr,
  output [55:0]  paddr_0,
  output         scIsSuccess_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_r = hitMeta_flag[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire [7:0] _hitRefillFlag_T_1 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 269:26]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  _hitCheck_T_7 = ~io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:31]
  wire  _hitLoad_T_1 = hitCheck & ~hitADCheck; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 276:26]
  wire  hitLoad = hitCheck & ~hitADCheck & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 276:41]
  wire  hitStore = _hitLoad_T_1 & hitFlag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:42]
  reg  io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
  reg  io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
  reg  io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
  reg  io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
  wire  _loadPF_T_5 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _loadPF_T_7 = ~hitLoad & _loadPF_T_5 & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:40]
  wire  _loadPF_T_8 = ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:50]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = raddrCancel ? 3'h5 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:59]
  wire  _GEN_16 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire  _loadPF_T_16 = _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:38]
  wire  _storePF_T_15 = io_in_bits_cmd[0] | ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 361:40]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire [2:0] _GEN_22 = is_reserved ? 3'h5 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 377:23]
  wire  _GEN_23 = is_reserved ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 371:32 378:24]
  wire  _GEN_24 = is_reserved ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 371:32 379:25]
  wire [2:0] _GEN_25 = ~missflag_v | ~missflag_r & missflag_w ? 3'h5 : _GEN_22; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:73]
  wire  _GEN_26 = ~missflag_v | ~missflag_r & missflag_w ? _loadPF_T_5 & _loadPF_T_8 : _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 360:22]
  wire  _GEN_27 = ~missflag_v | ~missflag_r & missflag_w ? io_in_bits_cmd[0] | ISAMO : _GEN_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 361:23]
  wire [55:0] _GEN_28 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_73 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_73; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u & _hitCheck_T_7); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a | ~missflag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:36]
  wire  _permLoad_T_5 = permCheck & ~_T_21 & ~permAD & ~misaligned; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 390:60]
  wire  permLoad = permCheck & ~_T_21 & ~permAD & ~misaligned & (missflag_r | io_pf_status_mxr & missflag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 390:75]
  wire  permStore = _permLoad_T_5 & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 391:76]
  wire [63:0] updateData = {56'h0,io_in_bits_cmd[0],7'h40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 392:31]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = _hitRefillFlag_T_1 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | updateData; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire [2:0] _GEN_29 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 3'h5 : 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 403:80 404:21 408:21]
  wire  _GEN_30 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit
     & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 403:80 405:22]
  wire  _GEN_31 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[
    0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 403:80 406:23]
  wire  _GEN_32 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 403:80 409:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_33 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_34 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire [2:0] _GEN_35 = level != 2'h0 ? _GEN_29 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_36 = level != 2'h0 ? _GEN_30 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 383:36]
  wire  _GEN_37 = level != 2'h0 ? _GEN_31 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 383:36]
  wire  _GEN_38 = level != 2'h0 & _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_39 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_48 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_67 = _T_12 ? _GEN_48 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_95 = 3'h2 == state ? _GEN_67 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_110 = 3'h1 == state ? 18'h3ffff : _GEN_95; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_110; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_40 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_41 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_25 : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_42 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_26 : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_43 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_27 : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_44 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_28 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_45 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_46 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_47 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_49 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_59 = _T_12 ? _GEN_41 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_61 = _T_12 ? _GEN_42 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 351:33]
  wire  _GEN_62 = _T_12 ? _GEN_43 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 351:33]
  wire  _GEN_66 = _T_12 & _GEN_47; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_69 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire [2:0] _GEN_70 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire [2:0] _GEN_72 = io_isFinish | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_74 = io_isFinish | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_75 = io_isFinish | alreadyOutFire ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire [2:0] _GEN_76 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_77 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_78 = 3'h4 == state ? _GEN_72 : _GEN_76; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_80 = 3'h4 == state ? _GEN_74 : _GEN_77; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_81 = 3'h4 == state ? _GEN_75 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_82 = 3'h3 == state ? _GEN_70 : _GEN_78; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_85 = 3'h3 == state ? missPTEAF : _GEN_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_86 = 3'h3 == state ? _GEN_2 : _GEN_81; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_89 = 3'h2 == state ? _GEN_61 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_90 = 3'h2 == state ? _GEN_62 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_104 = 3'h1 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_89; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_105 = 3'h1 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_90; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_109 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_66; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  loadPF = 3'h0 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_104; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  storePF = 3'h0 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_105; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_109; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _T_45 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_59 = ~scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:12]
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire [63:0] _GEN_79 = {{8'd0}, paddr}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:49]
  wire  _scIsSuccess_T_7 = hit | state == 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:81]
  wire  out_req_valid = io_in_valid & _scIsSuccess_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _ldReqAF_T_2 = paddr >= 56'h38000000 & paddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_5 = paddr >= 56'h3c000000 & paddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_8 = paddr >= 56'h40600000 & paddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_11 = paddr >= 56'h50000000 & paddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_14 = paddr >= 56'h40001000 & paddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_17 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_20 = paddr >= 56'h40002000 & paddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_23 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _ldReqAF_T_24 = {_ldReqAF_T_23,_ldReqAF_T_20,_ldReqAF_T_17,_ldReqAF_T_14,_ldReqAF_T_11,_ldReqAF_T_8,
    _ldReqAF_T_5,_ldReqAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _ldReqAF_T_25 = |_ldReqAF_T_24; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  ldReqAF = out_req_valid & ~_ldReqAF_T_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 489:34]
  wire  loadAF = (ldReqAF | missPTEAF) & _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 491:54]
  wire  storeAF = ldReqAF & io_in_bits_cmd[0] | ldReqAF & _loadPF_T_5 & ISAMO | missPTEAF & _storePF_T_15; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 492:79]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _hasException_T_2 = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  hasException = _hasException_T_2 | loadPF | storePF | loadAF | storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 494:72]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  wire  scIsSuccess = _T_59 | lr_0 & lr_addr == _GEN_79 | ~(hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:60]
  assign io_in_ready = io_out_ready & _T_45 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException & scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:92]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_windex = REG_1; // @[src/main/scala/nutcore/mem/TLB.scala 218:17]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_isFinish = _alreadyOutFire_T | _hasException_T_2 | ~scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:54]
  assign paddr_0 = paddr;
  assign scIsSuccess_0 = scIsSuccess;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
      io_pf_loadPF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= _GEN_61;
    end else begin
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
      io_pf_storePF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= _GEN_62;
    end else begin
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
      io_pf_laf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end else begin
      io_pf_laf_REG <= loadAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
      io_pf_saf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end else begin
      io_pf_saf_REG <= storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 342:15]
      end else begin
        state <= _GEN_15;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_59;
    end else begin
      state <= _GEN_82;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_69;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_46;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_49;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_44;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_86;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(_T_10)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
          missPTEAF <= _GEN_16;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_85;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else begin
      REG <= 3'h2 == state & _GEN_66;
    end
    REG_1 <= io_in_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_48;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_45;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= missMetaRefill & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed: SC is inflight but TLB receives a read request\n    at EmbeddedTLB.scala:476 assert(!scInflight || !io.in.valid || req.isWrite(), \"SC is inflight but TLB receives a read request\")\n"
            ); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  io_pf_loadPF_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_pf_storePF_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_pf_laf_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_pf_saf_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  level = _RAND_6[1:0];
  _RAND_7 = {2{`RANDOM}};
  memRespStore = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  missMaskStore = _RAND_8[17:0];
  _RAND_9 = {2{`RANDOM}};
  raddr = _RAND_9[55:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  missPTEAF = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_1 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  REG_2 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  REG_3 = _RAND_15[26:0];
  _RAND_16 = {1{`RANDOM}};
  REG_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  REG_5 = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  REG_6 = _RAND_18[7:0];
  _RAND_19 = {2{`RANDOM}};
  REG_7 = _RAND_19[43:0];
  _RAND_20 = {2{`RANDOM}};
  REG_8 = _RAND_20[55:0];
  _RAND_21 = {1{`RANDOM}};
  blockRefill = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
    end
  end
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [63:0] io_out_bits_wdata // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_rindex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  reg [3:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 4'hf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         lr,
  input         scInflight,
  input         amoReq,
  input  [63:0] lrAddr,
  output [55:0] paddr,
  input  [63:0] CSRSATP,
  output        _T_12_0,
  output        scIsSuccess_0,
  output        vmEnable_0,
  input         MOUFlushTLB,
  output        tlbFinish_0,
  output        _T_13_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_lr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_lr_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [55:0] tlbExec_paddr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_rindex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  _GEN_7 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _GEN_8 = mdUpdate & vmEnable | _GEN_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [2:0] tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [3:0] tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [7:0] tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [63:0] tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  _T_7 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_15 = _T_7 ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_8 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_16 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_15; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
  wire  _GEN_36 = tlbExec_io_out_valid & ~tlbExec_io_out_ready | alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:{37,37,37}]
  wire  _T_10 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _tlbFinish_T_2 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _tlbFinish_T_3 = tlbExec_io_pf_laf | tlbExec_io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _tlbFinish_T_4 = _tlbFinish_T_2 | _tlbFinish_T_3; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  tlbFinish = tlbExec_io_out_valid & ~alreadyOutFinish | _tlbFinish_T_4 | ~scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 180:95]
  wire  _T_12 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _T_13 = io_csrMMU_laf | io_csrMMU_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  EmbeddedTLBExec_1 tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_isFinish(tlbExec_io_isFinish),
    .lr_0(tlbExec_lr_0),
    .scInflight_0(tlbExec_scInflight_0),
    .ISAMO(tlbExec_ISAMO),
    .lr_addr(tlbExec_lr_addr),
    .paddr_0(tlbExec_paddr_0),
    .scIsSuccess_0(tlbExec_scIsSuccess_0)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19 149:23]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 148:24 169:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 169:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 163:26 169:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 164:25 169:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 165:27 169:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 166:27 169:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_csrMMU_loadPF = ~vmEnable ? 1'h0 : tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 150:24 95:17]
  assign io_csrMMU_storePF = ~vmEnable ? 1'h0 : tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 151:25 95:17]
  assign io_csrMMU_laf = ~vmEnable ? 1'h0 : tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 152:21 95:17]
  assign io_csrMMU_saf = ~vmEnable ? 1'h0 : tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 153:21 95:17]
  assign paddr = tlbExec_paddr_0;
  assign _T_12_0 = _T_12;
  assign scIsSuccess_0 = tlbExec_scIsSuccess_0;
  assign vmEnable_0 = vmEnable;
  assign tlbFinish_0 = tlbFinish;
  assign _T_13_1 = _T_13;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_size = tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_cmd = tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wmask = tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wdata = tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 src/main/scala/utils/Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_lr_0 = lr;
  assign tlbExec_scInflight_0 = scInflight;
  assign tlbExec_ISAMO = amoReq;
  assign tlbExec_lr_addr = lrAddr;
  assign tlbEmpty_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 147:29 169:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else begin
      valid <= _GEN_8;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_16;
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_addr <= tlbExec_io_out_bits_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_size <= tlbExec_io_out_bits_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_cmd <= tlbExec_io_out_bits_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wmask <= tlbExec_io_out_bits_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wdata <= tlbExec_io_out_bits_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
    end else if (alreadyOutFinish & _T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:53]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:72]
    end else begin
      alreadyOutFinish <= _GEN_36;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  valid_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  tlbEmpty_io_in_bits_r_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  alreadyOutFinish = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_fake_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_out_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_out_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_mmio_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        ismmio_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = io_in_resp_valid | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire [2:0] _GEN_9 = _GEN_3 ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [3:0] cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  reg [2:0] size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  reg [63:0] wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  reg [7:0] wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [3:0] mmiocmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [3:0] memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5; // @[src/main/scala/nutcore/mem/Cache.scala 601:30]
  assign io_in_resp_bits_cmd = ismmioRec ? mmiocmd : memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 609:29]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_out_mem_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_out_mem_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_out_mem_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_mmio_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mmio_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mmio_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  assign ismmio_0 = ismmio;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
      cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
      size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
      wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
      wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
      mmiocmd <= io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
      memcmd <= io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  alreadyOutFire = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reqaddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cmd = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  size = _RAND_5[2:0];
  _RAND_6 = {2{`RANDOM}};
  wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wmask = _RAND_7[7:0];
  _RAND_8 = {2{`RANDOM}};
  mmiordata = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  mmiocmd = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  memrdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  memcmd = _RAND_11[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_imem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_imem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_imem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_imem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_dmem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_dmem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [2:0]  io_dmem_mem_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_dmem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_dmem_mem_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_dmem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_dmem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_dmem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_extra_meip_0,
  output        isWFI,
  input         io_extra_mtip,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_reset; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_flushVec; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [1:0] frontend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_isWFI; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [11:0] frontend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  backend_clock; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_reset; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_flush; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_laf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_saf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_lr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_meip_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scInflight; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_amoReq; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_lrAddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [55:0] backend_paddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_satp; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scIsSuccess; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_mtip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_vmEnable; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [11:0] backend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_tlbFinish; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_ismmio; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_13_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_msip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  mmioXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_0_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [2:0] mmioXbar_io_in_1_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [2:0] mmioXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  dmemXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_2_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_2_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  itlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] itlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_imem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [1:0] io_imem_cache_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  dtlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] dtlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_lr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_amoReq; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_lrAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [55:0] dtlb_paddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_12_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_vmEnable_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_tlbFinish_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_13_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_1_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_dmem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_ismmio_0; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  reg [63:0] dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [1:0] ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  reg [1:0] ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] _ringBufferAllowin_T_1 = ringBufferHead + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire [1:0] _ringBufferAllowin_T_4 = ringBufferHead + 2'h2; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire  ringBufferAllowin = _ringBufferAllowin_T_1 != ringBufferTail & _ringBufferAllowin_T_4 != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 33:124]
  wire  needEnqueue_0 = frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 36:27 37:20]
  wire [1:0] enqueueSize = {{1'd0}, needEnqueue_0}; // @[src/main/scala/utils/PipelineVector.scala 40:44]
  wire  enqueueFire_0 = enqueueSize >= 2'h1; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  enqueueFire_1 = enqueueSize >= 2'h2; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  wen = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _T_1 = {{1'd0}, ringBufferHead}; // @[src/main/scala/utils/PipelineVector.scala 45:45]
  wire [63:0] _dataBuffer_T_cf_instr = needEnqueue_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pnpc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [3:0] _dataBuffer_T_cf_brIdx = needEnqueue_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [2:0] _dataBuffer_T_ctrl_fuType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [6:0] _dataBuffer_T_ctrl_fuOpType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc1 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc2 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfDest = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _dataBuffer_T_data_imm = needEnqueue_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _GEN_0 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_2 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_3 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_4 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_5 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_6 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_7 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_8 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_9 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_10 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_11 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_28 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_29 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_30 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_31 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_32 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_33 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_34 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_35 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_72 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_73 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_74 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_75 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_92 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_93 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_94 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_95 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_100 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_101 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_102 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_103 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_108 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_109 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_110 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_111 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_116 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_117 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_118 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_119 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_132 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_133 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_1_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_134 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_2_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_135 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_3_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_136 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_137 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_138 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_139 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_144 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_145 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_146 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_147 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_160 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_0_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_161 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_1_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_162 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_2_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_163 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_3_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_164 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_0_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_165 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_1_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_166 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_2_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_167 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_3_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_168 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_169 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_170 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_171 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_172 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_173 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_174 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_175 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_176 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_177 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_178 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_179 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_180 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_181 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_182 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_183 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_184 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_185 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_186 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_187 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_188 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_189 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_190 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_191 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_192 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_193 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_194 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_195 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_220 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_221 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_222 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_223 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_224 = enqueueFire_0 ? _GEN_0 : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_225 = enqueueFire_0 ? _GEN_1 : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_226 = enqueueFire_0 ? _GEN_2 : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_227 = enqueueFire_0 ? _GEN_3 : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_228 = enqueueFire_0 ? _GEN_4 : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_229 = enqueueFire_0 ? _GEN_5 : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_230 = enqueueFire_0 ? _GEN_6 : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_231 = enqueueFire_0 ? _GEN_7 : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_232 = enqueueFire_0 ? _GEN_8 : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_233 = enqueueFire_0 ? _GEN_9 : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_234 = enqueueFire_0 ? _GEN_10 : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_235 = enqueueFire_0 ? _GEN_11 : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_252 = enqueueFire_0 ? _GEN_28 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_253 = enqueueFire_0 ? _GEN_29 : dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_254 = enqueueFire_0 ? _GEN_30 : dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_255 = enqueueFire_0 ? _GEN_31 : dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_256 = enqueueFire_0 ? _GEN_32 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_257 = enqueueFire_0 ? _GEN_33 : dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_258 = enqueueFire_0 ? _GEN_34 : dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_259 = enqueueFire_0 ? _GEN_35 : dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_296 = enqueueFire_0 ? _GEN_72 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_297 = enqueueFire_0 ? _GEN_73 : dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_298 = enqueueFire_0 ? _GEN_74 : dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_299 = enqueueFire_0 ? _GEN_75 : dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_316 = enqueueFire_0 ? _GEN_92 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_317 = enqueueFire_0 ? _GEN_93 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_318 = enqueueFire_0 ? _GEN_94 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_319 = enqueueFire_0 ? _GEN_95 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_324 = enqueueFire_0 ? _GEN_100 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_325 = enqueueFire_0 ? _GEN_101 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_326 = enqueueFire_0 ? _GEN_102 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_327 = enqueueFire_0 ? _GEN_103 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_332 = enqueueFire_0 ? _GEN_108 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_333 = enqueueFire_0 ? _GEN_109 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_334 = enqueueFire_0 ? _GEN_110 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_335 = enqueueFire_0 ? _GEN_111 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_340 = enqueueFire_0 ? _GEN_116 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_341 = enqueueFire_0 ? _GEN_117 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_342 = enqueueFire_0 ? _GEN_118 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_343 = enqueueFire_0 ? _GEN_119 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_348 = enqueueFire_0 ? _GEN_124 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_349 = enqueueFire_0 ? _GEN_125 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_350 = enqueueFire_0 ? _GEN_126 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_351 = enqueueFire_0 ? _GEN_127 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_356 = enqueueFire_0 ? _GEN_132 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_357 = enqueueFire_0 ? _GEN_133 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_358 = enqueueFire_0 ? _GEN_134 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_359 = enqueueFire_0 ? _GEN_135 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_360 = enqueueFire_0 ? _GEN_136 : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_361 = enqueueFire_0 ? _GEN_137 : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_362 = enqueueFire_0 ? _GEN_138 : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_363 = enqueueFire_0 ? _GEN_139 : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_368 = enqueueFire_0 ? _GEN_144 : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_369 = enqueueFire_0 ? _GEN_145 : dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_370 = enqueueFire_0 ? _GEN_146 : dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_371 = enqueueFire_0 ? _GEN_147 : dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_384 = enqueueFire_0 ? _GEN_160 : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_385 = enqueueFire_0 ? _GEN_161 : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_386 = enqueueFire_0 ? _GEN_162 : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_387 = enqueueFire_0 ? _GEN_163 : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_388 = enqueueFire_0 ? _GEN_164 : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_389 = enqueueFire_0 ? _GEN_165 : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_390 = enqueueFire_0 ? _GEN_166 : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_391 = enqueueFire_0 ? _GEN_167 : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_392 = enqueueFire_0 ? _GEN_168 : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_393 = enqueueFire_0 ? _GEN_169 : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_394 = enqueueFire_0 ? _GEN_170 : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_395 = enqueueFire_0 ? _GEN_171 : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_396 = enqueueFire_0 ? _GEN_172 : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_397 = enqueueFire_0 ? _GEN_173 : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_398 = enqueueFire_0 ? _GEN_174 : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_399 = enqueueFire_0 ? _GEN_175 : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_400 = enqueueFire_0 ? _GEN_176 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_401 = enqueueFire_0 ? _GEN_177 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_402 = enqueueFire_0 ? _GEN_178 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_403 = enqueueFire_0 ? _GEN_179 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_404 = enqueueFire_0 ? _GEN_180 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_405 = enqueueFire_0 ? _GEN_181 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_406 = enqueueFire_0 ? _GEN_182 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_407 = enqueueFire_0 ? _GEN_183 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_408 = enqueueFire_0 ? _GEN_184 : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_409 = enqueueFire_0 ? _GEN_185 : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_410 = enqueueFire_0 ? _GEN_186 : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_411 = enqueueFire_0 ? _GEN_187 : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_412 = enqueueFire_0 ? _GEN_188 : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_413 = enqueueFire_0 ? _GEN_189 : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_414 = enqueueFire_0 ? _GEN_190 : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_415 = enqueueFire_0 ? _GEN_191 : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_416 = enqueueFire_0 ? _GEN_192 : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_417 = enqueueFire_0 ? _GEN_193 : dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_418 = enqueueFire_0 ? _GEN_194 : dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_419 = enqueueFire_0 ? _GEN_195 : dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_444 = enqueueFire_0 ? _GEN_220 : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_445 = enqueueFire_0 ? _GEN_221 : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_446 = enqueueFire_0 ? _GEN_222 : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_447 = enqueueFire_0 ? _GEN_223 : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [1:0] _T_4 = 2'h1 + ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 46:45]
  wire [1:0] _ringBufferHead_T_1 = ringBufferHead + enqueueSize; // @[src/main/scala/utils/PipelineVector.scala 47:42]
  wire [63:0] _GEN_1122 = 2'h1 == ringBufferTail ? dataBuffer_1_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1123 = 2'h2 == ringBufferTail ? dataBuffer_2_data_imm : _GEN_1122; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1150 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_isNutCoreTrap : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1151 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_isNutCoreTrap : _GEN_1150; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1154 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1155 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfDest : _GEN_1154; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1158 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1159 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfWen : _GEN_1158; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1162 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1163 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc2 : _GEN_1162; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1166 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1167 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc1 : _GEN_1166; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1170 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1171 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuOpType : _GEN_1170; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1174 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1175 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuType : _GEN_1174; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1178 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1179 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src2Type : _GEN_1178; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1182 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1183 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src1Type : _GEN_1182; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1198 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_crossBoundaryFault : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1199 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_crossBoundaryFault : _GEN_1198; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1206 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1207 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_brIdx : _GEN_1206; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1214 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1215 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_1 : _GEN_1214; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1222 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1223 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_3 : _GEN_1222; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1230 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1231 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_5 : _GEN_1230; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1238 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1239 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_7 : _GEN_1238; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1246 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1247 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_9 : _GEN_1246; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1254 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1255 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_11 : _GEN_1254; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1262 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_1 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1263 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_1 : _GEN_1262; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1266 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_2 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1267 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_2 : _GEN_1266; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1306 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_12 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1307 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_12 : _GEN_1306; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1334 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1335 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pnpc : _GEN_1334; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1338 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1339 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pc : _GEN_1338; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1342 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1343 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_instr : _GEN_1342; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _dequeueSize_T = backend_io_in_0_ready & backend_io_in_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] dequeueSize = {{1'd0}, _dequeueSize_T}; // @[src/main/scala/utils/PipelineVector.scala 64:42]
  wire  dequeueFire = dequeueSize > 2'h0; // @[src/main/scala/utils/PipelineVector.scala 65:35]
  wire [1:0] _ringBufferTail_T_1 = ringBufferTail + dequeueSize; // @[src/main/scala/utils/PipelineVector.scala 67:42]
  Frontend_inorder frontend ( // @[src/main/scala/nutcore/NutCore.scala 131:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(frontend_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(frontend_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_iaf(frontend_io_iaf),
    .io_sfence_vma_invalid(frontend_io_sfence_vma_invalid),
    .io_wfi_invalid(frontend_io_wfi_invalid),
    .REG_valid(frontend_REG_valid),
    .REG_pc(frontend_REG_pc),
    .REG_isMissPredict(frontend_REG_isMissPredict),
    .REG_actualTarget(frontend_REG_actualTarget),
    .REG_fuOpType(frontend_REG_fuOpType),
    .REG_btbType(frontend_REG_btbType),
    .REG_isRVC(frontend_REG_isRVC),
    .isWFI(frontend_isWFI),
    .flushICache(frontend_flushICache),
    .flushTLB(frontend_flushTLB),
    .intrVecIDU(frontend_intrVecIDU)
  );
  Backend_inorder backend ( // @[src/main/scala/nutcore/NutCore.scala 174:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(backend_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(backend_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(backend_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(backend_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(backend_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(backend_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(backend_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(backend_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(backend_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_laf(backend_io_memMMU_dmem_laf),
    .io_memMMU_dmem_saf(backend_io_memMMU_dmem_saf),
    .io_sfence_vma_invalid(backend_io_sfence_vma_invalid),
    .io_wfi_invalid(backend_io_wfi_invalid),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    .lr(backend_lr),
    .io_extra_meip_0(backend_io_extra_meip_0),
    .scInflight(backend_scInflight),
    .REG_valid(backend_REG_valid),
    .REG_pc(backend_REG_pc),
    .REG_isMissPredict(backend_REG_isMissPredict),
    .REG_actualTarget(backend_REG_actualTarget),
    .REG_fuOpType(backend_REG_fuOpType),
    .REG_btbType(backend_REG_btbType),
    .REG_isRVC(backend_REG_isRVC),
    .amoReq(backend_amoReq),
    .lrAddr(backend_lrAddr),
    .paddr(backend_paddr),
    .satp(backend_satp),
    ._T_12(backend__T_12),
    .scIsSuccess(backend_scIsSuccess),
    .io_extra_mtip(backend_io_extra_mtip),
    .flushICache(backend_flushICache),
    .vmEnable(backend_vmEnable),
    .flushTLB(backend_flushTLB),
    .intrVecIDU(backend_intrVecIDU),
    .tlbFinish(backend_tlbFinish),
    .ismmio(backend_ismmio),
    ._T_13_0(backend__T_13_0),
    .io_extra_msip(backend_io_extra_msip)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[src/main/scala/nutcore/NutCore.scala 178:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(mmioXbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(mmioXbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(mmioXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[src/main/scala/nutcore/NutCore.scala 179:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(dmemXbar_io_in_1_req_ready),
    .io_in_1_req_valid(dmemXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(dmemXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(dmemXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(dmemXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(dmemXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(dmemXbar_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(dmemXbar_io_in_2_req_ready),
    .io_in_2_req_valid(dmemXbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(dmemXbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(dmemXbar_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(dmemXbar_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(dmemXbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(dmemXbar_io_in_2_resp_bits_rdata),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  EmbeddedTLB itlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user),
    .io_mem_req_ready(itlb_io_mem_req_ready),
    .io_mem_req_valid(itlb_io_mem_req_valid),
    .io_mem_req_bits_addr(itlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(itlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(itlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(itlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(itlb_io_mem_resp_bits_rdata),
    .io_flush(itlb_io_flush),
    .io_csrMMU_priviledgeMode(itlb_io_csrMMU_priviledgeMode),
    .io_iaf(itlb_io_iaf),
    .CSRSATP(itlb_CSRSATP),
    .MOUFlushTLB(itlb_MOUFlushTLB)
  );
  PTERequestFilter filter ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_in_req_ready(filter_io_in_req_ready),
    .io_in_req_valid(filter_io_in_req_valid),
    .io_in_req_bits_addr(filter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_io_out_req_ready),
    .io_out_req_valid(filter_io_out_req_valid),
    .io_out_req_bits_addr(filter_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_io_out_resp_bits_rdata),
    .io_u(filter_io_u)
  );
  Cache_fake io_imem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_imem_cache_clock),
    .reset(io_imem_cache_reset),
    .io_in_req_ready(io_imem_cache_io_in_req_ready),
    .io_in_req_valid(io_imem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_imem_cache_io_in_req_bits_addr),
    .io_in_req_bits_user(io_imem_cache_io_in_req_bits_user),
    .io_in_resp_ready(io_imem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_imem_cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(io_imem_cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(io_imem_cache_io_in_resp_bits_user),
    .io_flush(io_imem_cache_io_flush),
    .io_out_mem_req_ready(io_imem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_imem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_imem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(io_imem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_imem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_rdata(io_imem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_imem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_imem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_imem_cache_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(io_imem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_imem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_imem_cache_io_mmio_resp_bits_rdata)
  );
  EmbeddedTLB_1 dtlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(dtlb_clock),
    .reset(dtlb_reset),
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata),
    .io_mem_req_ready(dtlb_io_mem_req_ready),
    .io_mem_req_valid(dtlb_io_mem_req_valid),
    .io_mem_req_bits_addr(dtlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(dtlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(dtlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(dtlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(dtlb_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(dtlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(dtlb_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(dtlb_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(dtlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(dtlb_io_csrMMU_storePF),
    .io_csrMMU_laf(dtlb_io_csrMMU_laf),
    .io_csrMMU_saf(dtlb_io_csrMMU_saf),
    .lr(dtlb_lr),
    .scInflight(dtlb_scInflight),
    .amoReq(dtlb_amoReq),
    .lrAddr(dtlb_lrAddr),
    .paddr(dtlb_paddr),
    .CSRSATP(dtlb_CSRSATP),
    ._T_12_0(dtlb__T_12_0),
    .scIsSuccess_0(dtlb_scIsSuccess_0),
    .vmEnable_0(dtlb_vmEnable_0),
    .MOUFlushTLB(dtlb_MOUFlushTLB),
    .tlbFinish_0(dtlb_tlbFinish_0),
    ._T_13_1(dtlb__T_13_1)
  );
  PTERequestFilter filter_1 ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_1_clock),
    .reset(filter_1_reset),
    .io_in_req_ready(filter_1_io_in_req_ready),
    .io_in_req_valid(filter_1_io_in_req_valid),
    .io_in_req_bits_addr(filter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_1_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_1_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_1_io_out_req_ready),
    .io_out_req_valid(filter_1_io_out_req_valid),
    .io_out_req_bits_addr(filter_1_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_1_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_1_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_1_io_out_resp_bits_rdata),
    .io_u(filter_1_io_u)
  );
  Cache_fake_1 io_dmem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_dmem_cache_clock),
    .reset(io_dmem_cache_reset),
    .io_in_req_ready(io_dmem_cache_io_in_req_ready),
    .io_in_req_valid(io_dmem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_dmem_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(io_dmem_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_dmem_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_dmem_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_dmem_cache_io_in_req_bits_wdata),
    .io_in_resp_valid(io_dmem_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_dmem_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_dmem_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(io_dmem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_dmem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_dmem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_size(io_dmem_cache_io_out_mem_req_bits_size),
    .io_out_mem_req_bits_cmd(io_dmem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wmask(io_dmem_cache_io_out_mem_req_bits_wmask),
    .io_out_mem_req_bits_wdata(io_dmem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(io_dmem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_dmem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_dmem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_dmem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_dmem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_dmem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_dmem_cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(io_dmem_cache_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(io_dmem_cache_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(io_dmem_cache_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(io_dmem_cache_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(io_dmem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_dmem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(io_dmem_cache_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(io_dmem_cache_io_mmio_resp_bits_rdata),
    .ismmio_0(io_dmem_cache_ismmio_0)
  );
  assign io_imem_mem_req_valid = io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_mem_req_bits_addr = io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_dmem_mem_req_valid = io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_addr = io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_size = io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_cmd = io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wmask = io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wdata = io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign isWFI = frontend_isWFI;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_out_0_ready = ringBufferAllowin | ~frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_iaf = itlb_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 189:21]
  assign frontend_io_sfence_vma_invalid = backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 215:36]
  assign frontend_io_wfi_invalid = backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 216:29]
  assign frontend_REG_valid = backend_REG_valid;
  assign frontend_REG_pc = backend_REG_pc;
  assign frontend_REG_isMissPredict = backend_REG_isMissPredict;
  assign frontend_REG_actualTarget = backend_REG_actualTarget;
  assign frontend_REG_fuOpType = backend_REG_fuOpType;
  assign frontend_REG_btbType = backend_REG_btbType;
  assign frontend_REG_isRVC = backend_REG_isRVC;
  assign frontend_flushICache = backend_flushICache;
  assign frontend_flushTLB = backend_flushTLB;
  assign frontend_intrVecIDU = backend_intrVecIDU;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = ringBufferHead != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 2'h3 == ringBufferTail ? dataBuffer_3_cf_instr : _GEN_1343; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pc : _GEN_1339; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pnpc : _GEN_1335; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_1 : _GEN_1263; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_2 : _GEN_1267; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_12 : _GEN_1307; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_1 : _GEN_1215; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_3 : _GEN_1223; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_5 : _GEN_1231; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_7 : _GEN_1239; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_9 : _GEN_1247; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_11 : _GEN_1255; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 2'h3 == ringBufferTail ? dataBuffer_3_cf_brIdx : _GEN_1207; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_crossBoundaryFault = 2'h3 == ringBufferTail ? dataBuffer_3_cf_crossBoundaryFault :
    _GEN_1199; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src1Type : _GEN_1183; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src2Type : _GEN_1179; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuType : _GEN_1175; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuOpType : _GEN_1171; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc1 : _GEN_1167; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc2 : _GEN_1163; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfWen : _GEN_1159; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfDest : _GEN_1155; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_isNutCoreTrap = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_isNutCoreTrap : _GEN_1151; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 2'h3 == ringBufferTail ? dataBuffer_3_data_imm : _GEN_1123; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[src/main/scala/nutcore/NutCore.scala 219:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_memMMU_dmem_loadPF = dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_storePF = dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_laf = dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_saf = dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_extra_meip_0 = io_extra_meip_0;
  assign backend_paddr = dtlb_paddr;
  assign backend__T_12 = dtlb__T_12_0;
  assign backend_scIsSuccess = dtlb_scIsSuccess_0;
  assign backend_io_extra_mtip = io_extra_mtip;
  assign backend_vmEnable = dtlb_vmEnable_0;
  assign backend_tlbFinish = dtlb_tlbFinish_0;
  assign backend_ismmio = io_dmem_cache_ismmio_0;
  assign backend__T_13_0 = dtlb__T_13_1;
  assign backend_io_extra_msip = io_extra_msip;
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_0_req_bits_addr = io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_valid = io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_addr = io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_size = io_dmem_cache_io_mmio_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_cmd = io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wmask = io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wdata = io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_1_req_valid = filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_addr = filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_cmd = filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_wdata = filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_valid = filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_addr = filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_cmd = filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_wdata = filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_out_req_ready = io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_valid = io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_cmd = io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_rdata = io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_out_req_ready = io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_valid = io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_rdata = io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_user = io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_mem_req_ready = filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_valid = filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_bits_rdata = filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_flush = frontend_io_flushVec[0]; // @[src/main/scala/nutcore/NutCore.scala 184:35]
  assign itlb_io_csrMMU_priviledgeMode = backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign itlb_CSRSATP = backend_satp;
  assign itlb_MOUFlushTLB = backend_flushTLB;
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_in_req_valid = itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_addr = itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_cmd = itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_wdata = itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_out_req_ready = dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_valid = dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_bits_rdata = dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_u = backend_io_memMMU_imem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_imem_cache_clock = clock;
  assign io_imem_cache_reset = reset;
  assign io_imem_cache_io_in_req_valid = itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/NutCore.scala 193:19]
  assign io_imem_cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign dtlb_clock = clock;
  assign dtlb_reset = reset;
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_mem_req_ready = filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_valid = filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_bits_rdata = filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_csrMMU_priviledgeMode = backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_sum = backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_mxr = backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_lr = backend_lr;
  assign dtlb_scInflight = backend_scInflight;
  assign dtlb_amoReq = backend_amoReq;
  assign dtlb_lrAddr = backend_lrAddr;
  assign dtlb_CSRSATP = backend_satp;
  assign dtlb_MOUFlushTLB = backend_flushTLB;
  assign filter_1_clock = clock;
  assign filter_1_reset = reset;
  assign filter_1_io_in_req_valid = dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_addr = dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_cmd = dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_wdata = dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_out_req_ready = dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_valid = dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_bits_rdata = dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_u = backend_io_memMMU_dmem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_dmem_cache_clock = clock;
  assign io_dmem_cache_reset = reset;
  assign io_dmem_cache_io_in_req_valid = dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_cmd = mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_instr <= _GEN_224;
        end
      end else begin
        dataBuffer_0_cf_instr <= _GEN_224;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pc <= _GEN_228;
        end
      end else begin
        dataBuffer_0_cf_pc <= _GEN_228;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pnpc <= _GEN_232;
        end
      end else begin
        dataBuffer_0_cf_pnpc <= _GEN_232;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_1 <= _GEN_252;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_1 <= _GEN_252;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_2 <= _GEN_256;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_2 <= _GEN_256;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_12 <= _GEN_296;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_12 <= _GEN_296;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_1 <= _GEN_316;
        end
      end else begin
        dataBuffer_0_cf_intrVec_1 <= _GEN_316;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_3 <= _GEN_324;
        end
      end else begin
        dataBuffer_0_cf_intrVec_3 <= _GEN_324;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_5 <= _GEN_332;
        end
      end else begin
        dataBuffer_0_cf_intrVec_5 <= _GEN_332;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_7 <= _GEN_340;
        end
      end else begin
        dataBuffer_0_cf_intrVec_7 <= _GEN_340;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_9 <= _GEN_348;
        end
      end else begin
        dataBuffer_0_cf_intrVec_9 <= _GEN_348;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_11 <= _GEN_356;
        end
      end else begin
        dataBuffer_0_cf_intrVec_11 <= _GEN_356;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_brIdx <= _GEN_360;
        end
      end else begin
        dataBuffer_0_cf_brIdx <= _GEN_360;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_crossBoundaryFault <= _GEN_368;
        end
      end else begin
        dataBuffer_0_cf_crossBoundaryFault <= _GEN_368;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src1Type <= _GEN_384;
        end
      end else begin
        dataBuffer_0_ctrl_src1Type <= _GEN_384;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src2Type <= _GEN_388;
        end
      end else begin
        dataBuffer_0_ctrl_src2Type <= _GEN_388;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuType <= _GEN_392;
        end
      end else begin
        dataBuffer_0_ctrl_fuType <= _GEN_392;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuOpType <= _GEN_396;
        end
      end else begin
        dataBuffer_0_ctrl_fuOpType <= _GEN_396;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc1 <= _GEN_400;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc1 <= _GEN_400;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc2 <= _GEN_404;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc2 <= _GEN_404;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfWen <= _GEN_408;
        end
      end else begin
        dataBuffer_0_ctrl_rfWen <= _GEN_408;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfDest <= _GEN_412;
        end
      end else begin
        dataBuffer_0_ctrl_rfDest <= _GEN_412;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_416;
        end
      end else begin
        dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_416;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_data_imm <= _GEN_444;
        end
      end else begin
        dataBuffer_0_data_imm <= _GEN_444;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_instr <= _GEN_225;
        end
      end else begin
        dataBuffer_1_cf_instr <= _GEN_225;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pc <= _GEN_229;
        end
      end else begin
        dataBuffer_1_cf_pc <= _GEN_229;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pnpc <= _GEN_233;
        end
      end else begin
        dataBuffer_1_cf_pnpc <= _GEN_233;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_1 <= _GEN_253;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_1 <= _GEN_253;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_2 <= _GEN_257;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_2 <= _GEN_257;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_12 <= _GEN_297;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_12 <= _GEN_297;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_1 <= _GEN_317;
        end
      end else begin
        dataBuffer_1_cf_intrVec_1 <= _GEN_317;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_3 <= _GEN_325;
        end
      end else begin
        dataBuffer_1_cf_intrVec_3 <= _GEN_325;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_5 <= _GEN_333;
        end
      end else begin
        dataBuffer_1_cf_intrVec_5 <= _GEN_333;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_7 <= _GEN_341;
        end
      end else begin
        dataBuffer_1_cf_intrVec_7 <= _GEN_341;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_9 <= _GEN_349;
        end
      end else begin
        dataBuffer_1_cf_intrVec_9 <= _GEN_349;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_11 <= _GEN_357;
        end
      end else begin
        dataBuffer_1_cf_intrVec_11 <= _GEN_357;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_brIdx <= _GEN_361;
        end
      end else begin
        dataBuffer_1_cf_brIdx <= _GEN_361;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_crossBoundaryFault <= _GEN_369;
        end
      end else begin
        dataBuffer_1_cf_crossBoundaryFault <= _GEN_369;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src1Type <= _GEN_385;
        end
      end else begin
        dataBuffer_1_ctrl_src1Type <= _GEN_385;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src2Type <= _GEN_389;
        end
      end else begin
        dataBuffer_1_ctrl_src2Type <= _GEN_389;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuType <= _GEN_393;
        end
      end else begin
        dataBuffer_1_ctrl_fuType <= _GEN_393;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuOpType <= _GEN_397;
        end
      end else begin
        dataBuffer_1_ctrl_fuOpType <= _GEN_397;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc1 <= _GEN_401;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc1 <= _GEN_401;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc2 <= _GEN_405;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc2 <= _GEN_405;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfWen <= _GEN_409;
        end
      end else begin
        dataBuffer_1_ctrl_rfWen <= _GEN_409;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfDest <= _GEN_413;
        end
      end else begin
        dataBuffer_1_ctrl_rfDest <= _GEN_413;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_417;
        end
      end else begin
        dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_417;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_data_imm <= _GEN_445;
        end
      end else begin
        dataBuffer_1_data_imm <= _GEN_445;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_instr <= _GEN_226;
        end
      end else begin
        dataBuffer_2_cf_instr <= _GEN_226;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pc <= _GEN_230;
        end
      end else begin
        dataBuffer_2_cf_pc <= _GEN_230;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pnpc <= _GEN_234;
        end
      end else begin
        dataBuffer_2_cf_pnpc <= _GEN_234;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_1 <= _GEN_254;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_1 <= _GEN_254;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_2 <= _GEN_258;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_2 <= _GEN_258;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_12 <= _GEN_298;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_12 <= _GEN_298;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_1 <= _GEN_318;
        end
      end else begin
        dataBuffer_2_cf_intrVec_1 <= _GEN_318;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_3 <= _GEN_326;
        end
      end else begin
        dataBuffer_2_cf_intrVec_3 <= _GEN_326;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_5 <= _GEN_334;
        end
      end else begin
        dataBuffer_2_cf_intrVec_5 <= _GEN_334;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_7 <= _GEN_342;
        end
      end else begin
        dataBuffer_2_cf_intrVec_7 <= _GEN_342;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_9 <= _GEN_350;
        end
      end else begin
        dataBuffer_2_cf_intrVec_9 <= _GEN_350;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_11 <= _GEN_358;
        end
      end else begin
        dataBuffer_2_cf_intrVec_11 <= _GEN_358;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_brIdx <= _GEN_362;
        end
      end else begin
        dataBuffer_2_cf_brIdx <= _GEN_362;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_crossBoundaryFault <= _GEN_370;
        end
      end else begin
        dataBuffer_2_cf_crossBoundaryFault <= _GEN_370;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src1Type <= _GEN_386;
        end
      end else begin
        dataBuffer_2_ctrl_src1Type <= _GEN_386;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src2Type <= _GEN_390;
        end
      end else begin
        dataBuffer_2_ctrl_src2Type <= _GEN_390;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuType <= _GEN_394;
        end
      end else begin
        dataBuffer_2_ctrl_fuType <= _GEN_394;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuOpType <= _GEN_398;
        end
      end else begin
        dataBuffer_2_ctrl_fuOpType <= _GEN_398;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc1 <= _GEN_402;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc1 <= _GEN_402;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc2 <= _GEN_406;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc2 <= _GEN_406;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfWen <= _GEN_410;
        end
      end else begin
        dataBuffer_2_ctrl_rfWen <= _GEN_410;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfDest <= _GEN_414;
        end
      end else begin
        dataBuffer_2_ctrl_rfDest <= _GEN_414;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_418;
        end
      end else begin
        dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_418;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_data_imm <= _GEN_446;
        end
      end else begin
        dataBuffer_2_data_imm <= _GEN_446;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_instr <= _GEN_227;
        end
      end else begin
        dataBuffer_3_cf_instr <= _GEN_227;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pc <= _GEN_231;
        end
      end else begin
        dataBuffer_3_cf_pc <= _GEN_231;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pnpc <= _GEN_235;
        end
      end else begin
        dataBuffer_3_cf_pnpc <= _GEN_235;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_1 <= _GEN_255;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_1 <= _GEN_255;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_2 <= _GEN_259;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_2 <= _GEN_259;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_12 <= _GEN_299;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_12 <= _GEN_299;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_1 <= _GEN_319;
        end
      end else begin
        dataBuffer_3_cf_intrVec_1 <= _GEN_319;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_3 <= _GEN_327;
        end
      end else begin
        dataBuffer_3_cf_intrVec_3 <= _GEN_327;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_5 <= _GEN_335;
        end
      end else begin
        dataBuffer_3_cf_intrVec_5 <= _GEN_335;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_7 <= _GEN_343;
        end
      end else begin
        dataBuffer_3_cf_intrVec_7 <= _GEN_343;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_9 <= _GEN_351;
        end
      end else begin
        dataBuffer_3_cf_intrVec_9 <= _GEN_351;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_11 <= _GEN_359;
        end
      end else begin
        dataBuffer_3_cf_intrVec_11 <= _GEN_359;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_brIdx <= _GEN_363;
        end
      end else begin
        dataBuffer_3_cf_brIdx <= _GEN_363;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_crossBoundaryFault <= _GEN_371;
        end
      end else begin
        dataBuffer_3_cf_crossBoundaryFault <= _GEN_371;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src1Type <= _GEN_387;
        end
      end else begin
        dataBuffer_3_ctrl_src1Type <= _GEN_387;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src2Type <= _GEN_391;
        end
      end else begin
        dataBuffer_3_ctrl_src2Type <= _GEN_391;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuType <= _GEN_395;
        end
      end else begin
        dataBuffer_3_ctrl_fuType <= _GEN_395;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuOpType <= _GEN_399;
        end
      end else begin
        dataBuffer_3_ctrl_fuOpType <= _GEN_399;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc1 <= _GEN_403;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc1 <= _GEN_403;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc2 <= _GEN_407;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc2 <= _GEN_407;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfWen <= _GEN_411;
        end
      end else begin
        dataBuffer_3_ctrl_rfWen <= _GEN_411;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfDest <= _GEN_415;
        end
      end else begin
        dataBuffer_3_ctrl_rfDest <= _GEN_415;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_419;
        end
      end else begin
        dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_419;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_data_imm <= _GEN_447;
        end
      end else begin
        dataBuffer_3_data_imm <= _GEN_447;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 30:33]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 72:24]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      ringBufferHead <= _ringBufferHead_T_1; // @[src/main/scala/utils/PipelineVector.scala 47:24]
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 31:33]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 73:24]
    end else if (dequeueFire) begin // @[src/main/scala/utils/PipelineVector.scala 66:22]
      ringBufferTail <= _ringBufferTail_T_1; // @[src/main/scala/utils/PipelineVector.scala 67:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataBuffer_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dataBuffer_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  dataBuffer_0_cf_crossBoundaryFault = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  dataBuffer_0_ctrl_isNutCoreTrap = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  dataBuffer_0_data_imm = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  dataBuffer_1_cf_instr = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  dataBuffer_1_cf_pc = _RAND_25[38:0];
  _RAND_26 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_12 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  dataBuffer_1_cf_crossBoundaryFault = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  dataBuffer_1_ctrl_isNutCoreTrap = _RAND_46[0:0];
  _RAND_47 = {2{`RANDOM}};
  dataBuffer_1_data_imm = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  dataBuffer_2_cf_instr = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  dataBuffer_2_cf_pc = _RAND_49[38:0];
  _RAND_50 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc = _RAND_50[38:0];
  _RAND_51 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  dataBuffer_2_cf_crossBoundaryFault = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  dataBuffer_2_ctrl_isNutCoreTrap = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  dataBuffer_2_data_imm = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  dataBuffer_3_cf_instr = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  dataBuffer_3_cf_pc = _RAND_73[38:0];
  _RAND_74 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc = _RAND_74[38:0];
  _RAND_75 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  dataBuffer_3_cf_crossBoundaryFault = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1 = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  dataBuffer_3_ctrl_isNutCoreTrap = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  dataBuffer_3_data_imm = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  ringBufferHead = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  ringBufferTail = _RAND_97[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_in_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_in_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_out_mem_resp_bits_rdata // @[src/main/scala/system/Coherence.scala 31:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/system/Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[src/main/scala/system/Coherence.scala 46:24]
  wire  _reqLatch_T = ~inflight; // @[src/main/scala/system/Coherence.scala 52:42]
  reg [31:0] reqLatch_addr; // @[src/main/scala/system/Coherence.scala 52:27]
  wire  _io_out_mem_req_valid_T_1 = io_in_req_valid & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 65:43]
  wire  _T_20 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_31 = io_in_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_31 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 89:{60,68}]
  wire  _T_34 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = _T_34 ? 3'h4 : state; // @[src/main/scala/system/Coherence.scala 45:22 94:{36,44}]
  wire  _T_36 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_37 = io_out_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [2:0] _GEN_16 = _T_36 & _T_37 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 96:101 45:22 96:93]
  wire [2:0] _GEN_17 = _T_36 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 97:{57,65}]
  wire [2:0] _GEN_18 = 3'h5 == state ? _GEN_17 : state; // @[src/main/scala/system/Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_16 : _GEN_18; // @[src/main/scala/system/Coherence.scala 74:18]
  wire [31:0] _GEN_20 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_25 = 3'h3 == state | _io_out_mem_req_valid_T_1; // @[src/main/scala/system/Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_26 = 3'h3 == state ? _GEN_15 : _GEN_19; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_28 = 3'h2 == state ? 1'h0 : io_out_mem_resp_valid; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_29 = 3'h2 == state ? 4'h0 : io_out_mem_resp_bits_cmd; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_30 = 3'h2 == state ? 64'h0 : io_out_mem_resp_bits_rdata; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [31:0] _GEN_32 = 3'h2 == state ? io_in_req_bits_addr : _GEN_20; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_37 = 3'h2 == state ? _io_out_mem_req_valid_T_1 : _GEN_25; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_40 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_28; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_41 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_29; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_42 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_30; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [31:0] _GEN_43 = 3'h1 == state ? io_in_req_bits_addr : _GEN_32; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_48 = 3'h1 == state ? _io_out_mem_req_valid_T_1 : _GEN_37; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_in_req_ready = io_out_mem_req_ready & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 66:43]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_40; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_41; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_42; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _io_out_mem_req_valid_T_1 : _GEN_48; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_43; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/system/Coherence.scala 72:14]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/system/Coherence.scala 45:22]
      state <= 3'h0; // @[src/main/scala/system/Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (_T_20) begin // @[src/main/scala/system/Coherence.scala 76:29]
        state <= 3'h4;
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (3'h2 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
        state <= _GEN_14;
      end else begin
        state <= _GEN_26;
      end
    end
    if (~inflight) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_addr <= io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 52:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/system/Coherence.scala 49:9]
    end
  end
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_aw_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_aw_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [1:0]  io_out_aw_bits_burst, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [1:0]  io_out_ar_bits_burst, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _io_out_ar_bits_len_T_1 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:30]
  wire  _io_out_w_bits_last_T = io_in_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _io_out_w_bits_last_T_1 = io_in_req_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [2:0] _io_in_resp_bits_cmd_T = io_out_r_bits_last ? 3'h6 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:28]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 & io_out_w_bits_last | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _wAck_T_1 = _wSend_T_1 & io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 188:41]
  wire  _GEN_2 = _wAck_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _io_in_resp_bits_cmd_T}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_len = io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_size = io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_aw_bits_burst = io_out_ar_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_w_bits_last = _io_out_w_bits_last_T | _io_out_w_bits_last_T_1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 177:54]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_ar_bits_len = {{5'd0}, _io_out_ar_bits_len_T_1}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:24]
  assign io_out_ar_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 170:24]
  assign io_out_ar_bits_burst = 2'h2; // @[src/main/scala/bus/simplebus/ToAXI4.scala 171:24]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
  end
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_out_2_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h80000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [2:0] _outSelVec_enc_T = outMatchVec_2 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _outSelVec_enc_T_1 = outMatchVec_1 ? 3'h2 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] outSelVec_enc = outMatchVec_0 ? 3'h1 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [2:0] _reqInvalidAddr_T = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire [1:0] _GEN_5 = io_in_resp_valid ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  _io_in_req_ready_T_4 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_4 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_5 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_6 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_7 = outSelRespVec_2 ? io_out_2_resp_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_8 = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_req_ready = _io_in_req_ready_T_4 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_4 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_8 | _io_in_resp_bits_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_3 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
  end
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_mtip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_msip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         isWFI_0,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  reg [63:0] freq_reg; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire [15:0] freq = freq_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 38:22]
  reg [63:0] inc_reg; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire [15:0] inc = inc_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 40:20]
  reg [15:0] cnt; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[src/main/scala/device/AXI4CLINT.scala 43:21]
  wire  tick = nextCnt == freq; // @[src/main/scala/device/AXI4CLINT.scala 45:23]
  wire [63:0] _GEN_15 = {{48'd0}, inc}; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_1 = mtime + _GEN_15; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_3 = mtime + 64'h186a0; // @[src/main/scala/device/AXI4CLINT.scala 51:35]
  wire [7:0] _T_11 = io__in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_12 = io__in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_13 = io__in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_14 = io__in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_15 = io__in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_16 = io__in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_17 = io__in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_18 = io__in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_19 = {_T_18,_T_17,_T_16,_T_15,_T_14,_T_13,_T_12,_T_11}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _io_in_r_bits_data_T = 16'h0 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 16'h8000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 16'hbff8 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 16'h8008 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_4 = 16'h4000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T ? msip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_1 ? freq_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_2 ? mtime : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_8 = _io_in_r_bits_data_T_3 ? inc_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_4 ? mtimecmp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_5 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_11 = _io_in_r_bits_data_T_10 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_12 = _io_in_r_bits_data_T_11 | _io_in_r_bits_data_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _msip_T = io__in_w_bits_data & _T_19; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _msip_T_1 = ~_T_19; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _msip_T_2 = msip & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _msip_T_3 = _msip_T | _msip_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _freq_reg_T_2 = freq_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _freq_reg_T_3 = _msip_T | _freq_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtime_T_6 = mtime & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtime_T_7 = _msip_T | _mtime_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _inc_reg_T_2 = inc_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _inc_reg_T_3 = _msip_T | _inc_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtimecmp_T_2 = mtimecmp & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtimecmp_T_3 = _msip_T | _mtimecmp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  reg  io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = _io_in_r_bits_data_T_12 | _io_in_r_bits_data_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__extra_mtip = io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:21]
  assign io__extra_msip = io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'hbff8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtime <= _mtime_T_7; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (isWFI_0) begin // @[src/main/scala/device/AXI4CLINT.scala 51:18]
      mtime <= _mtime_T_3; // @[src/main/scala/device/AXI4CLINT.scala 51:26]
    end else if (tick) begin // @[src/main/scala/device/AXI4CLINT.scala 46:15]
      mtime <= _mtime_T_1; // @[src/main/scala/device/AXI4CLINT.scala 46:23]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h4000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtimecmp <= _mtimecmp_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      msip <= _msip_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 37:25]
      freq_reg <= 64'h2710; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      freq_reg <= _freq_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 39:24]
      inc_reg <= 64'h1; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8008) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      inc_reg <= _inc_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 42:20]
      cnt <= 16'h0; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end else if (nextCnt < freq) begin // @[src/main/scala/device/AXI4CLINT.scala 44:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    io_extra_mtip_REG <= mtime >= mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 66:38]
    io_extra_msip_REG <= msip != 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 67:37]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  freq_reg = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inc_reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  io_extra_mtip_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_extra_msip_REG = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
  end
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_meip_0, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  reg [31:0] enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  wire [7:0] _T_12 = io__in_w_bits_strb >> io__in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4PLIC.scala 89:85]
  wire [7:0] _T_21 = _T_12[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_22 = _T_12[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_23 = _T_12[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_24 = _T_12[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_25 = _T_12[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_26 = _T_12[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_27 = _T_12[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_28 = _T_12[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_29 = {_T_28,_T_27,_T_26,_T_25,_T_24,_T_23,_T_22,_T_21}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T_1 = 26'h2000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 26'h4 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 26'h200000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_6 = _rdata_T_1 ? enable_0_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_8 = _rdata_T_3 ? priority_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_9 = _rdata_T_4 ? threshold_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_6 | _rdata_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] rdata = _rdata_T_12 | _rdata_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _enable_0_0_T = io__in_w_bits_data[31:0] & _T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _enable_0_0_T_1 = ~_T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _enable_0_0_T_2 = enable_0_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _enable_0_0_T_3 = _enable_0_0_T | _enable_0_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _priority_0_T_2 = priority_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _priority_0_T_3 = _enable_0_0_T | _priority_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _threshold_0_T_2 = threshold_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _threshold_0_T_3 = _enable_0_0_T | _threshold_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = {rdata,rdata}; // @[src/main/scala/device/AXI4PLIC.scala 91:25]
  assign io__extra_meip_0 = 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      priority_0 <= _priority_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h2000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      enable_0_0 <= _enable_0_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      threshold_0 <= _threshold_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  enable_0_0 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  threshold_0 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_aw_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_aw_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_aw_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_aw_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mem_aw_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  output [1:0]  io_mem_aw_bits_burst, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_w_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mem_w_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_w_bits_strb, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_b_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_ar_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_ar_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_ar_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_ar_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mem_ar_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mem_r_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_req_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_req_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_resp_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_resp_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/system/NutShell.scala 45:14]
);
  wire  nutcore_clock; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_reset; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [2:0] nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_isWFI; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  cohMg_clock; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_reset; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  xbar_clock; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_reset; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_in_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  io_mem_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_aw_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_aw_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [1:0] io_mem_bridge_io_out_aw_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [1:0] io_mem_bridge_io_out_ar_bits_burst; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  clint_clock; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_reset; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [7:0] clint_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_isWFI_0; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] clint_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_clock; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_reset; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [7:0] plic_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] plic_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  NutCore nutcore ( // @[src/main/scala/system/NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_size(nutcore_io_dmem_mem_req_bits_size),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wmask(nutcore_io_dmem_mem_req_bits_wmask),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .isWFI(nutcore_isWFI),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_msip(nutcore_io_extra_msip)
  );
  CoherenceManager cohMg ( // @[src/main/scala/system/NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[src/main/scala/system/NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  SimpleBusAddressMapper memAddrMap ( // @[src/main/scala/system/NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_size(memAddrMap_io_in_req_bits_size),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(memAddrMap_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_size(memAddrMap_io_out_req_bits_size),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(memAddrMap_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter io_mem_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(io_mem_bridge_clock),
    .reset(io_mem_bridge_reset),
    .io_in_req_ready(io_mem_bridge_io_in_req_ready),
    .io_in_req_valid(io_mem_bridge_io_in_req_valid),
    .io_in_req_bits_addr(io_mem_bridge_io_in_req_bits_addr),
    .io_in_req_bits_size(io_mem_bridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_mem_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_mem_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_mem_bridge_io_in_req_bits_wdata),
    .io_in_resp_valid(io_mem_bridge_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_mem_bridge_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_mem_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(io_mem_bridge_io_out_aw_ready),
    .io_out_aw_valid(io_mem_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(io_mem_bridge_io_out_aw_bits_addr),
    .io_out_aw_bits_len(io_mem_bridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(io_mem_bridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(io_mem_bridge_io_out_aw_bits_burst),
    .io_out_w_ready(io_mem_bridge_io_out_w_ready),
    .io_out_w_valid(io_mem_bridge_io_out_w_valid),
    .io_out_w_bits_data(io_mem_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(io_mem_bridge_io_out_w_bits_strb),
    .io_out_w_bits_last(io_mem_bridge_io_out_w_bits_last),
    .io_out_b_valid(io_mem_bridge_io_out_b_valid),
    .io_out_ar_ready(io_mem_bridge_io_out_ar_ready),
    .io_out_ar_valid(io_mem_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(io_mem_bridge_io_out_ar_bits_addr),
    .io_out_ar_bits_len(io_mem_bridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(io_mem_bridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(io_mem_bridge_io_out_ar_bits_burst),
    .io_out_r_valid(io_mem_bridge_io_out_r_valid),
    .io_out_r_bits_data(io_mem_bridge_io_out_r_bits_data),
    .io_out_r_bits_last(io_mem_bridge_io_out_r_bits_last)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[src/main/scala/system/NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_cmd(mmioXbar_io_out_2_resp_bits_cmd),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  AXI4CLINT clint ( // @[src/main/scala/system/NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_aw_ready(clint_io__in_aw_ready),
    .io__in_aw_valid(clint_io__in_aw_valid),
    .io__in_aw_bits_addr(clint_io__in_aw_bits_addr),
    .io__in_w_ready(clint_io__in_w_ready),
    .io__in_w_valid(clint_io__in_w_valid),
    .io__in_w_bits_data(clint_io__in_w_bits_data),
    .io__in_w_bits_strb(clint_io__in_w_bits_strb),
    .io__in_b_ready(clint_io__in_b_ready),
    .io__in_b_valid(clint_io__in_b_valid),
    .io__in_ar_ready(clint_io__in_ar_ready),
    .io__in_ar_valid(clint_io__in_ar_valid),
    .io__in_ar_bits_addr(clint_io__in_ar_bits_addr),
    .io__in_r_ready(clint_io__in_r_ready),
    .io__in_r_valid(clint_io__in_r_valid),
    .io__in_r_bits_data(clint_io__in_r_bits_data),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .isWFI_0(clint_isWFI_0),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_1 clint_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(clint_io_in_bridge_clock),
    .reset(clint_io_in_bridge_reset),
    .io_in_req_ready(clint_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(clint_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(clint_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(clint_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(clint_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(clint_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(clint_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(clint_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(clint_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(clint_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(clint_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(clint_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(clint_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(clint_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(clint_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(clint_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(clint_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(clint_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(clint_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(clint_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(clint_io_in_bridge_io_out_r_bits_data)
  );
  AXI4PLIC plic ( // @[src/main/scala/system/NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_aw_ready(plic_io__in_aw_ready),
    .io__in_aw_valid(plic_io__in_aw_valid),
    .io__in_aw_bits_addr(plic_io__in_aw_bits_addr),
    .io__in_w_ready(plic_io__in_w_ready),
    .io__in_w_valid(plic_io__in_w_valid),
    .io__in_w_bits_data(plic_io__in_w_bits_data),
    .io__in_w_bits_strb(plic_io__in_w_bits_strb),
    .io__in_b_ready(plic_io__in_b_ready),
    .io__in_b_valid(plic_io__in_b_valid),
    .io__in_ar_ready(plic_io__in_ar_ready),
    .io__in_ar_valid(plic_io__in_ar_valid),
    .io__in_ar_bits_addr(plic_io__in_ar_bits_addr),
    .io__in_r_ready(plic_io__in_r_ready),
    .io__in_r_valid(plic_io__in_r_valid),
    .io__in_r_bits_data(plic_io__in_r_bits_data),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_1 plic_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(plic_io_in_bridge_clock),
    .reset(plic_io_in_bridge_reset),
    .io_in_req_ready(plic_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(plic_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(plic_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(plic_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(plic_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(plic_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(plic_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(plic_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(plic_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(plic_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(plic_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(plic_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(plic_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(plic_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(plic_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(plic_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(plic_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(plic_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(plic_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(plic_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(plic_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(plic_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(plic_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(plic_io_in_bridge_io_out_r_bits_data)
  );
  assign io_mem_aw_valid = io_mem_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_addr = io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_len = io_mem_bridge_io_out_aw_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_size = io_mem_bridge_io_out_aw_bits_size; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_burst = io_mem_bridge_io_out_aw_bits_burst; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_valid = io_mem_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_data = io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_strb = io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_last = io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_valid = io_mem_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_addr = io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_len = io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_size = io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mmio_req_valid = mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_resp_ready = mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_out_req_ready = memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_valid = memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_valid = xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_addr = xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_size = xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_cmd = xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wmask = xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wdata = xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_out_req_ready = io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_clock = clock;
  assign io_mem_bridge_reset = reset;
  assign io_mem_bridge_io_in_req_valid = memAddrMap_io_out_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_size = memAddrMap_io_out_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wmask = memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_out_aw_ready = io_mem_aw_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_w_ready = io_mem_w_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_b_valid = io_mem_b_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_ar_ready = io_mem_ar_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_valid = io_mem_r_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_data = io_mem_r_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_last = io_mem_r_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_valid = io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_aw_valid = clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_aw_bits_addr = clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_valid = clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_data = clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_strb = clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_b_ready = clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_valid = clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_bits_addr = clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_r_ready = clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_isWFI_0 = nutcore_isWFI;
  assign clint_io_in_bridge_clock = clock;
  assign clint_io_in_bridge_reset = reset;
  assign clint_io_in_bridge_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_out_aw_ready = clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_w_ready = clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_b_valid = clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_ar_ready = clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_valid = clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_bits_data = clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_aw_valid = plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_aw_bits_addr = plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_valid = plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_data = plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_strb = plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_b_ready = plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_valid = plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_bits_addr = plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_r_ready = plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_clock = clock;
  assign plic_io_in_bridge_reset = reset;
  assign plic_io_in_bridge_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_out_aw_ready = plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_w_ready = plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_b_valid = plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_ar_ready = plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_valid = plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_bits_data = plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
endmodule
module DifftestMem1P(
  input         clock,
  input         reset,
  input         read_valid, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input  [63:0] read_index, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  output [63:0] read_data_0, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input         write_valid, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_index, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_data_0, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_mask_0 // @[difftest/src/main/scala/common/Mem.scala 204:17]
);
  wire  helper_0_r_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_w_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_mask; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_clock; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  _T_1 = ~reset; // @[difftest/src/main/scala/common/Mem.scala 214:16]
  wire [64:0] _T_3 = read_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 215:26]
  wire [65:0] _T_4 = {{1'd0}, _T_3}; // @[difftest/src/main/scala/common/Mem.scala 215:39]
  wire [64:0] _T_9 = write_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 223:27]
  wire [65:0] _T_10 = {{1'd0}, _T_9}; // @[difftest/src/main/scala/common/Mem.scala 223:40]
  MemRWHelper helper_0 ( // @[difftest/src/main/scala/common/Mem.scala 197:49]
    .r_enable(helper_0_r_enable),
    .r_index(helper_0_r_index),
    .r_data(helper_0_r_data),
    .w_enable(helper_0_w_enable),
    .w_index(helper_0_w_index),
    .w_data(helper_0_w_data),
    .w_mask(helper_0_w_mask),
    .clock(helper_0_clock)
  );
  assign read_data_0 = helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 211:13]
  assign helper_0_r_enable = ~reset & read_valid; // @[difftest/src/main/scala/common/Mem.scala 214:30]
  assign helper_0_r_index = _T_4[63:0]; // @[difftest/src/main/scala/common/Mem.scala 102:13]
  assign helper_0_w_enable = _T_1 & write_valid; // @[difftest/src/main/scala/common/Mem.scala 222:30]
  assign helper_0_w_index = _T_10[63:0]; // @[difftest/src/main/scala/common/Mem.scala 150:13]
  assign helper_0_w_data = write_data_0; // @[difftest/src/main/scala/common/Mem.scala 151:12]
  assign helper_0_w_mask = write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 152:12]
  assign helper_0_clock = clock; // @[difftest/src/main/scala/common/Mem.scala 220:13]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~(~read_valid | ~write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed: read and write come at the same cycle\n    at Mem.scala:263 assert(!read.valid || !write.valid, \"read and write come at the same cycle\")\n"
            ); // @[difftest/src/main/scala/common/Mem.scala 263:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (_T_1) begin
      assert(~read_valid | ~write_valid); // @[difftest/src/main/scala/common/Mem.scala 263:9]
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_bits_last, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [1:0]  io_in_ar_bits_burst, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_bits_last // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  rdata_mem_clock; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_reset; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_read_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_write_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  reg [7:0] c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [7:0] readBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _len_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [7:0] len_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [7:0] _GEN_0 = _len_T ? io_in_ar_bits_len : len_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg [1:0] burst_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [1:0] _GEN_1 = _len_T ? io_in_ar_bits_burst : burst_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [31:0] _wrapAddr_WIRE = {{24'd0}, io_in_ar_bits_len}; // @[src/main/scala/device/AXI4Slave.scala 45:{69,69}]
  wire [38:0] _GEN_32 = {{7'd0}, _wrapAddr_WIRE}; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T = _GEN_32 << io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T_1 = ~_wrapAddr_T; // @[src/main/scala/device/AXI4Slave.scala 45:42]
  wire [38:0] _GEN_19 = {{7'd0}, io_in_ar_bits_addr}; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  wire [38:0] wrapAddr = _GEN_19 & _wrapAddr_T_1; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  reg [38:0] raddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [38:0] _GEN_2 = _len_T ? wrapAddr : raddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [7:0] _value_T_1 = readBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [7:0] _GEN_3 = _GEN_1 == 2'h2 & readBeatCnt == _GEN_0 ? 8'h0 : _value_T_1; // @[src/main/scala/device/AXI4Slave.scala 50:{77,93} src/main/scala/chisel3/util/Counter.scala 77:15]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  wire [7:0] _GEN_4 = ren ? _GEN_3 : readBeatCnt; // @[src/main/scala/device/AXI4Slave.scala 48:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] _value_T_3 = c_value + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [31:0] _value_T_4 = io_in_ar_bits_addr >> io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 57:45]
  wire [31:0] _value_T_5 = _value_T_4 & _wrapAddr_WIRE; // @[src/main/scala/device/AXI4Slave.scala 57:67]
  wire  _T_7 = io_in_ar_bits_len != 8'h0 & io_in_ar_bits_burst == 2'h2; // @[src/main/scala/device/AXI4Slave.scala 58:40]
  wire  _T_11 = io_in_ar_bits_len == 8'h7; // @[src/main/scala/device/AXI4Slave.scala 60:30]
  wire  _T_12 = io_in_ar_bits_len == 8'h1 | io_in_ar_bits_len == 8'h3 | _T_11; // @[src/main/scala/device/AXI4Slave.scala 59:71]
  wire  _T_14 = _T_12 | io_in_ar_bits_len == 8'hf; // @[src/main/scala/device/AXI4Slave.scala 60:38]
  wire [31:0] _GEN_7 = _len_T ? _value_T_5 : {{24'd0}, _GEN_4}; // @[src/main/scala/device/AXI4Slave.scala 56:29 57:23]
  wire  _r_busy_T_2 = io_in_r_valid & io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 70:56]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_8 = _r_busy_T_2 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_9 = _len_T | _GEN_8; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_valid_T_2 = ren & (_len_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_10 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_11 = _io_in_r_valid_T_2 | _GEN_10; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [7:0] writeBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _waddr_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [31:0] waddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [31:0] _GEN_12 = _waddr_T ? io_in_aw_bits_addr : waddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  _T_18 = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [7:0] _value_T_7 = writeBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_15 = io_in_b_valid ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_16 = _waddr_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T_1 = _T_18 & io_in_w_bits_last; // @[src/main/scala/device/AXI4Slave.scala 97:43]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_17 = io_in_b_valid ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_18 = _io_in_b_valid_T_1 | _GEN_17; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = _GEN_12 & 32'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [28:0] _GEN_21 = {{21'd0}, writeBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T[31:3] + _GEN_21; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [38:0] _rIdx_T = _GEN_2 & 39'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [35:0] _GEN_22 = {{28'd0}, readBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [35:0] rIdx = _rIdx_T[38:3] + _GEN_22; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'h10000000; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire [31:0] rdata_lo = {io_in_w_bits_data[31:24],io_in_w_bits_data[23:16],io_in_w_bits_data[15:8],io_in_w_bits_data[7:
    0]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [31:0] rdata_hi = {io_in_w_bits_data[63:56],io_in_w_bits_data[55:48],io_in_w_bits_data[47:40],io_in_w_bits_data[
    39:32]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [7:0] _rdata_T_18 = io_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_19 = io_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_20 = io_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_21 = io_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_22 = io_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_23 = io_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_24 = io_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [7:0] _rdata_T_25 = io_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[difftest/src/main/scala/common/Mem.scala 248:45]
  wire [31:0] rdata_lo_1 = {_rdata_T_21,_rdata_T_20,_rdata_T_19,_rdata_T_18}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  wire [31:0] rdata_hi_1 = {_rdata_T_25,_rdata_T_24,_rdata_T_23,_rdata_T_22}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  reg  rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  reg  rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  reg [63:0] rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire [63:0] _rdata_T_28_0 = rdata_REG ? rdata_mem_read_data_0 : rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:8]
  wire [31:0] rdata_lo_2 = {_rdata_T_28_0[31:24],_rdata_T_28_0[23:16],_rdata_T_28_0[15:8],_rdata_T_28_0[7:0]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] rdata_hi_2 = {_rdata_T_28_0[63:56],_rdata_T_28_0[55:48],_rdata_T_28_0[47:40],_rdata_T_28_0[39:32]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] _GEN_28 = reset ? 32'h0 : _GEN_7; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  DifftestMem1P rdata_mem ( // @[difftest/src/main/scala/common/Mem.scala 322:36]
    .clock(rdata_mem_clock),
    .reset(rdata_mem_reset),
    .read_valid(rdata_mem_read_valid),
    .read_index(rdata_mem_read_index),
    .read_data_0(rdata_mem_read_data_0),
    .write_valid(rdata_mem_write_valid),
    .write_index(rdata_mem_write_index),
    .write_data_0(rdata_mem_write_data_0),
    .write_mask_0(rdata_mem_write_mask_0)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {rdata_hi_2,rdata_lo_2}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  assign io_in_r_bits_last = c_value == _GEN_0; // @[src/main/scala/device/AXI4Slave.scala 47:36]
  assign rdata_mem_clock = clock;
  assign rdata_mem_reset = reset;
  assign rdata_mem_read_valid = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  assign rdata_mem_read_index = {{28'd0}, rIdx}; // @[difftest/src/main/scala/common/Mem.scala 237:16]
  assign rdata_mem_write_valid = _T_18 & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 37:25]
  assign rdata_mem_write_index = {{35'd0}, wIdx};
  assign rdata_mem_write_data_0 = {rdata_hi,rdata_lo}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  assign rdata_mem_write_mask_0 = {rdata_hi_1,rdata_lo_1}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      c_value <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_in_r_valid) begin // @[src/main/scala/device/AXI4Slave.scala 52:28]
      if (io_in_r_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 54:33]
        c_value <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 54:43]
      end else begin
        c_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    readBeatCnt <= _GEN_28[7:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= 8'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= io_in_ar_bits_len; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= io_in_ar_bits_burst; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= 39'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= wrapAddr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _len_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_11;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T_18) begin // @[src/main/scala/device/AXI4Slave.scala 82:28]
      if (io_in_w_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 84:33]
        writeBeatCnt <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 84:43]
      end else begin
        writeBeatCnt <= _value_T_7; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= 32'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_waddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= io_in_aw_bits_addr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_16;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_18;
    end
    rdata_REG <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    rdata_REG_1 <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    if (rdata_REG_1) begin // @[difftest/src/main/scala/common/Mem.scala 238:42]
      rdata_r_0 <= rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_len_T & _T_7 & ~reset & ~_T_14) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at AXI4Slave.scala:59 assert(axi4.ar.bits.len === 1.U || axi4.ar.bits.len === 3.U ||\n"
            ); // @[src/main/scala/device/AXI4Slave.scala 59:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_value = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  readBeatCnt = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  len_r = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  burst_r = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  raddr_r = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  ren_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_busy = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  writeBeatCnt = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  waddr_r = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  w_busy = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rdata_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rdata_REG_1 = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  rdata_r_0 = _RAND_14[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_len_T & _T_7 & ~reset) begin
      assert(_T_14); // @[src/main/scala/device/AXI4Slave.scala 59:17]
    end
  end
endmodule
module LatencyPipe(
  output        io_in_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [7:0]  io_in_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [1:0]  io_in_bits_burst, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_out_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [7:0]  io_out_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [1:0]  io_out_bits_burst // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_len = io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_burst = io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
endmodule
module AXI4Delayer(
  output        io_in_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_aw_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [2:0]  io_in_aw_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [1:0]  io_in_aw_bits_burst, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_ar_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [1:0]  io_out_ar_bits_burst, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
);
  wire  io_out_ar_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_ar_pipe_io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_ar_pipe_io_out_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_aw_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_aw_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_aw_pipe_io_in_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_aw_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_aw_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [1:0] io_out_aw_pipe_io_out_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  LatencyPipe io_out_ar_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .io_in_ready(io_out_ar_pipe_io_in_ready),
    .io_in_valid(io_out_ar_pipe_io_in_valid),
    .io_in_bits_addr(io_out_ar_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_ar_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_ar_pipe_io_in_bits_size),
    .io_in_bits_burst(io_out_ar_pipe_io_in_bits_burst),
    .io_out_ready(io_out_ar_pipe_io_out_ready),
    .io_out_valid(io_out_ar_pipe_io_out_valid),
    .io_out_bits_addr(io_out_ar_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_ar_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_ar_pipe_io_out_bits_size),
    .io_out_bits_burst(io_out_ar_pipe_io_out_bits_burst)
  );
  LatencyPipe io_out_aw_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .io_in_ready(io_out_aw_pipe_io_in_ready),
    .io_in_valid(io_out_aw_pipe_io_in_valid),
    .io_in_bits_addr(io_out_aw_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_aw_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_aw_pipe_io_in_bits_size),
    .io_in_bits_burst(io_out_aw_pipe_io_in_bits_burst),
    .io_out_ready(io_out_aw_pipe_io_out_ready),
    .io_out_valid(io_out_aw_pipe_io_out_valid),
    .io_out_bits_addr(io_out_aw_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_aw_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_aw_pipe_io_out_bits_size),
    .io_out_bits_burst(io_out_aw_pipe_io_out_bits_burst)
  );
  assign io_in_aw_ready = io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_w_ready = io_out_w_ready; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_in_b_valid = io_out_b_valid; // @[src/main/scala/bus/axi4/Delayer.scala 18:13]
  assign io_in_ar_ready = io_out_ar_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_r_valid = io_out_r_valid; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_data = io_out_r_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_last = io_out_r_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_out_aw_valid = io_out_aw_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_aw_bits_addr = io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_w_valid = io_in_w_valid; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_data = io_in_w_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_strb = io_in_w_bits_strb; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_last = io_in_w_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_ar_valid = io_out_ar_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_addr = io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_len = io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_size = io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_burst = io_out_ar_pipe_io_out_bits_burst; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_pipe_io_in_valid = io_in_ar_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_addr = io_in_ar_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_len = io_in_ar_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_size = io_in_ar_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_burst = 2'h2; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_out_ready = 1'h1; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_aw_pipe_io_in_valid = io_in_aw_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_addr = io_in_aw_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_len = io_in_aw_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_size = io_in_aw_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_burst = io_in_aw_bits_burst; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_out_ready = io_out_aw_ready; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
endmodule
module SimpleBusCrossbar1toN_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_3_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_3_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_4_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_4_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_4_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_4_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_4_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h40600010; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h50000000 & io_in_req_bits_addr < 32'h50400000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40001000 & io_in_req_bits_addr < 32'h40001008; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_3 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h40001000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_4 = io_in_req_bits_addr >= 32'h40002000 & io_in_req_bits_addr < 32'h40003000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [4:0] _outSelVec_enc_T = outMatchVec_4 ? 5'h10 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_1 = outMatchVec_3 ? 5'h8 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_2 = outMatchVec_2 ? 5'h4 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_3 = outMatchVec_1 ? 5'h2 : _outSelVec_enc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] outSelVec_enc = outMatchVec_0 ? 5'h1 : _outSelVec_enc_T_3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_3 = outSelVec_enc[3]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_4 = outSelVec_enc[4]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [4:0] _reqInvalidAddr_T = {outSelVec_4,outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire  _T_7 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_7 = _T_7 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  _io_in_req_ready_T_8 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready | outSelVec_3 & io_out_3_req_ready | outSelVec_4 & io_out_4_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_8 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid | outSelRespVec_3 & io_out_3_resp_valid | outSelRespVec_4 &
    io_out_4_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = outSelRespVec_3 ? io_out_3_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_4 = outSelRespVec_4 ? io_out_4_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_5 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_6 = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_7 = _io_in_resp_bits_T_6 | _io_in_resp_bits_T_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_9 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_10 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_11 = outSelRespVec_2 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_12 = outSelRespVec_3 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_13 = outSelRespVec_4 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_14 = _io_in_resp_bits_T_9 | _io_in_resp_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_15 = _io_in_resp_bits_T_14 | _io_in_resp_bits_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_16 = _io_in_resp_bits_T_15 | _io_in_resp_bits_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_req_ready = _io_in_req_ready_T_8 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_8 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_16 | _io_in_resp_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_7 | _io_in_resp_bits_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_3_req_valid = outSelVec_3 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_3_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_resp_ready = outSelRespVec_3 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_4_req_valid = outSelVec_4 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_4_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_resp_ready = outSelRespVec_4 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_7;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= outSelVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= outSelVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  outSelRespVec_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  outSelRespVec_4 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
  end
endmodule
module AXI4UART(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_out_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_out_ch, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_in_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_extra_in_ch // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] txfifo; // @[src/main/scala/device/AXI4UART.scala 29:19]
  reg [31:0] stat; // @[src/main/scala/device/AXI4UART.scala 30:21]
  reg [31:0] ctrl; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire  _io_extra_out_valid_T_1 = io_in_aw_bits_addr[3:0] == 4'h4; // @[src/main/scala/device/AXI4UART.scala 33:41]
  wire [7:0] _T_5 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4UART.scala 45:79]
  wire [7:0] _T_14 = _T_5[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_15 = _T_5[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_16 = _T_5[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_17 = _T_5[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_18 = _T_5[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_19 = _T_5[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_20 = _T_5[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_21 = _T_5[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_22 = {_T_21,_T_20,_T_19,_T_18,_T_17,_T_16,_T_15,_T_14}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 4'hc == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [7:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T ? io_extra_in_ch : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_1 ? txfifo : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_2 ? stat : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_3 ? ctrl : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_11 = {{24'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_8 = _GEN_11 | _io_in_r_bits_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_8 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_9 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _txfifo_T = io_in_w_bits_data[31:0] & _T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _txfifo_T_1 = ~_T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _txfifo_T_2 = txfifo & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _txfifo_T_3 = _txfifo_T | _txfifo_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _stat_T_2 = stat & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _stat_T_3 = _txfifo_T | _stat_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _ctrl_T_2 = ctrl & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _ctrl_T_3 = _txfifo_T | _ctrl_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_10}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_out_valid = io_in_aw_bits_addr[3:0] == 4'h4 & _io_in_b_valid_T; // @[src/main/scala/device/AXI4UART.scala 33:49]
  assign io_extra_out_ch = io_in_w_bits_data[7:0]; // @[src/main/scala/device/AXI4UART.scala 34:40]
  assign io_extra_in_valid = io_in_ar_bits_addr[3:0] == 4'h0 & _r_busy_T_1; // @[src/main/scala/device/AXI4UART.scala 35:48]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & _io_extra_out_valid_T_1) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      txfifo <= _txfifo_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 30:21]
      stat <= 32'h1; // @[src/main/scala/device/AXI4UART.scala 30:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      stat <= _stat_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 31:21]
      ctrl <= 32'h0; // @[src/main/scala/device/AXI4UART.scala 31:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'hc) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      ctrl <= _ctrl_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  txfifo = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stat = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_sync // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _io_in_r_bits_data_T_2 = _io_in_r_bits_data_T ? 32'h190012c : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_r_bits_data_T_3 = _io_in_r_bits_data_T_1 & _w_busy_T; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_8 = {{31'd0}, _io_in_r_bits_data_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T_2 | _GEN_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_sync = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4RAM_1(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] rdata_mem_0 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_1 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_2 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_3 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_4 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_5 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_6 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_7 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_r_valid ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = io_in_aw_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _wIdx_T_2 = {{1'd0}, _wIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [31:0] _rIdx_T = io_in_ar_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _rIdx_T_2 = {{1'd0}, _rIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [28:0] rIdx = _rIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'hea60; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire [63:0] _rdata_T_12 = {rdata_mem_7_rdata_MPORT_1_data,rdata_mem_6_rdata_MPORT_1_data,
    rdata_mem_5_rdata_MPORT_1_data,rdata_mem_4_rdata_MPORT_1_data,rdata_mem_3_rdata_MPORT_1_data,
    rdata_mem_2_rdata_MPORT_1_data,rdata_mem_1_rdata_MPORT_1_data,rdata_mem_0_rdata_MPORT_1_data}; // @[src/main/scala/device/AXI4RAM.scala 55:18]
  reg [63:0] rdata; // @[src/main/scala/device/AXI4RAM.scala 55:14]
  assign rdata_mem_0_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_0_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_1[7:0] :
    rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_data = io_in_w_bits_data[7:0];
  assign rdata_mem_0_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_0_rdata_MPORT_mask = io_in_w_bits_strb[0];
  assign rdata_mem_0_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_1_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_1_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_3[7:0] :
    rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_data = io_in_w_bits_data[15:8];
  assign rdata_mem_1_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_1_rdata_MPORT_mask = io_in_w_bits_strb[1];
  assign rdata_mem_1_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_2_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_2_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_5[7:0] :
    rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_data = io_in_w_bits_data[23:16];
  assign rdata_mem_2_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_2_rdata_MPORT_mask = io_in_w_bits_strb[2];
  assign rdata_mem_2_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_3_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_3_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_7[7:0] :
    rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_data = io_in_w_bits_data[31:24];
  assign rdata_mem_3_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_3_rdata_MPORT_mask = io_in_w_bits_strb[3];
  assign rdata_mem_3_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_4_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_4_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_9[7:0] :
    rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_data = io_in_w_bits_data[39:32];
  assign rdata_mem_4_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_4_rdata_MPORT_mask = io_in_w_bits_strb[4];
  assign rdata_mem_4_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_5_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_5_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_11[7:0] :
    rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_data = io_in_w_bits_data[47:40];
  assign rdata_mem_5_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_5_rdata_MPORT_mask = io_in_w_bits_strb[5];
  assign rdata_mem_5_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_6_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_6_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_13[7:0] :
    rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_data = io_in_w_bits_data[55:48];
  assign rdata_mem_6_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_6_rdata_MPORT_mask = io_in_w_bits_strb[6];
  assign rdata_mem_6_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_7_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_7_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_15[7:0] :
    rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_data = io_in_w_bits_data[63:56];
  assign rdata_mem_7_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_7_rdata_MPORT_mask = io_in_w_bits_strb[7];
  assign rdata_mem_7_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = rdata; // @[src/main/scala/device/AXI4RAM.scala 58:18]
  always @(posedge clock) begin
    if (rdata_mem_0_rdata_MPORT_en & rdata_mem_0_rdata_MPORT_mask) begin
      rdata_mem_0[rdata_mem_0_rdata_MPORT_addr] <= rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_1_rdata_MPORT_en & rdata_mem_1_rdata_MPORT_mask) begin
      rdata_mem_1[rdata_mem_1_rdata_MPORT_addr] <= rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_2_rdata_MPORT_en & rdata_mem_2_rdata_MPORT_mask) begin
      rdata_mem_2[rdata_mem_2_rdata_MPORT_addr] <= rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_3_rdata_MPORT_en & rdata_mem_3_rdata_MPORT_mask) begin
      rdata_mem_3[rdata_mem_3_rdata_MPORT_addr] <= rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_4_rdata_MPORT_en & rdata_mem_4_rdata_MPORT_mask) begin
      rdata_mem_4[rdata_mem_4_rdata_MPORT_addr] <= rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_5_rdata_MPORT_en & rdata_mem_5_rdata_MPORT_mask) begin
      rdata_mem_5[rdata_mem_5_rdata_MPORT_addr] <= rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_6_rdata_MPORT_en & rdata_mem_6_rdata_MPORT_mask) begin
      rdata_mem_6[rdata_mem_6_rdata_MPORT_addr] <= rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_7_rdata_MPORT_en & rdata_mem_7_rdata_MPORT_mask) begin
      rdata_mem_7[rdata_mem_7_rdata_MPORT_addr] <= rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (ren_REG) begin // @[src/main/scala/device/AXI4RAM.scala 55:14]
      rdata <= _rdata_T_12; // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ren_REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  rdata = _RAND_21[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_fb_aw_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [63:0] io_in_fb_w_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [7:0]  io_in_fb_w_bits_strb, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_ctrl_ar_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output [63:0] io_in_ctrl_r_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_vga_valid // @[src/main/scala/device/AXI4VGA.scala 117:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  fb_clock; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_reset; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fbHelper_clk; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_valid; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire [31:0] fbHelper_pixel; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_sync; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  _io_in_fb_r_valid_T = io_in_fb_ar_ready & io_in_fb_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _io_in_fb_r_valid_T_1 = io_in_fb_r_ready & io_in_fb_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _io_in_fb_r_valid_T_1 ? 1'h0 : io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _io_in_fb_r_valid_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [10:0] hCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = hCounter == 11'h41f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [10:0] _wrap_value_T_1 = hCounter + 11'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg [9:0] vCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap_1 = vCounter == 10'h273; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [9:0] _wrap_value_T_3 = vCounter + 10'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  hInRange = hCounter >= 11'ha8 & hCounter < 11'h3c8; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  vInRange = vCounter >= 10'h5 & vCounter < 10'h25d; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[src/main/scala/device/AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 152:31]
  wire  _nextPixel_T_2 = hCounter >= 11'ha7 & hCounter < 11'h3c7; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  nextPixel = _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
  wire  _fbPixelAddrV0_T_1 = nextPixel & ~vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  fbPixelAddrV0_wrap_wrap = fbPixelAddrV0 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV0_wrap_value_T_1 = fbPixelAddrV0 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _fbPixelAddrV1_T = nextPixel & vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  fbPixelAddrV1_wrap_wrap = fbPixelAddrV1 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV1_wrap_value_T_1 = fbPixelAddrV1 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [16:0] _fb_io_in_ar_bits_addr_T = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[src/main/scala/device/AXI4VGA.scala 161:35]
  wire [18:0] _fb_io_in_ar_bits_addr_T_1 = {_fb_io_in_ar_bits_addr_T,2'h0}; // @[src/main/scala/device/AXI4VGA.scala 161:31]
  reg  fb_io_in_ar_valid_REG; // @[src/main/scala/device/AXI4VGA.scala 162:31]
  wire  _data_T = fb_io_in_r_ready & fb_io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] data_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] _GEN_14 = _data_T ? fb_io_in_r_bits_data : data_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  VGACtrl ctrl ( // @[src/main/scala/device/AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_aw_ready(ctrl_io_in_aw_ready),
    .io_in_aw_valid(ctrl_io_in_aw_valid),
    .io_in_w_ready(ctrl_io_in_w_ready),
    .io_in_w_valid(ctrl_io_in_w_valid),
    .io_in_b_ready(ctrl_io_in_b_ready),
    .io_in_b_valid(ctrl_io_in_b_valid),
    .io_in_ar_ready(ctrl_io_in_ar_ready),
    .io_in_ar_valid(ctrl_io_in_ar_valid),
    .io_in_ar_bits_addr(ctrl_io_in_ar_bits_addr),
    .io_in_r_ready(ctrl_io_in_r_ready),
    .io_in_r_valid(ctrl_io_in_r_valid),
    .io_in_r_bits_data(ctrl_io_in_r_bits_data),
    .io_extra_sync(ctrl_io_extra_sync)
  );
  AXI4RAM_1 fb ( // @[src/main/scala/device/AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_aw_ready(fb_io_in_aw_ready),
    .io_in_aw_valid(fb_io_in_aw_valid),
    .io_in_aw_bits_addr(fb_io_in_aw_bits_addr),
    .io_in_w_ready(fb_io_in_w_ready),
    .io_in_w_valid(fb_io_in_w_valid),
    .io_in_w_bits_data(fb_io_in_w_bits_data),
    .io_in_w_bits_strb(fb_io_in_w_bits_strb),
    .io_in_b_ready(fb_io_in_b_ready),
    .io_in_b_valid(fb_io_in_b_valid),
    .io_in_ar_ready(fb_io_in_ar_ready),
    .io_in_ar_valid(fb_io_in_ar_valid),
    .io_in_ar_bits_addr(fb_io_in_ar_bits_addr),
    .io_in_r_ready(fb_io_in_r_ready),
    .io_in_r_valid(fb_io_in_r_valid),
    .io_in_r_bits_data(fb_io_in_r_bits_data)
  );
  FBHelper fbHelper ( // @[src/main/scala/device/AXI4VGA.scala 171:26]
    .clk(fbHelper_clk),
    .valid(fbHelper_valid),
    .pixel(fbHelper_pixel),
    .sync(fbHelper_sync)
  );
  assign io_in_fb_aw_ready = fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign io_in_fb_w_ready = fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign io_in_fb_b_valid = fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign io_in_fb_ar_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 133:21]
  assign io_in_fb_r_valid = io_in_fb_r_valid_r; // @[src/main/scala/device/AXI4VGA.scala 136:20]
  assign io_in_ctrl_aw_ready = ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_w_ready = ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_b_valid = ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_ar_ready = ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_valid = ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_bits_data = ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_vga_valid = hInRange & vInRange; // @[src/main/scala/device/AXI4VGA.scala 148:28]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_aw_valid = io_in_ctrl_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_w_valid = io_in_ctrl_w_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_b_ready = io_in_ctrl_b_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_valid = io_in_ctrl_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_bits_addr = io_in_ctrl_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_r_ready = io_in_ctrl_r_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_aw_valid = io_in_fb_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_aw_bits_addr = io_in_fb_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_w_valid = io_in_fb_w_valid; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_data = io_in_fb_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_strb = io_in_fb_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_b_ready = io_in_fb_b_ready; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign fb_io_in_ar_valid = fb_io_in_ar_valid_REG & hCounterIs2; // @[src/main/scala/device/AXI4VGA.scala 162:43]
  assign fb_io_in_ar_bits_addr = {{13'd0}, _fb_io_in_ar_bits_addr_T_1}; // @[src/main/scala/device/AXI4VGA.scala 161:25]
  assign fb_io_in_r_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 164:20]
  assign fbHelper_clk = clock; // @[src/main/scala/device/AXI4VGA.scala 172:21]
  assign fbHelper_valid = io_vga_valid; // @[src/main/scala/device/AXI4VGA.scala 173:23]
  assign fbHelper_pixel = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[src/main/scala/device/AXI4VGA.scala 167:23]
  assign fbHelper_sync = ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 175:22]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_fb_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_fb_r_valid_r <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
    end else begin
      hCounter <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (wrap_wrap_1) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        vCounter <= _wrap_value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV0_T_1) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV0_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV0 <= _fbPixelAddrV0_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV1_T) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV1_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV1 <= _fbPixelAddrV1_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    fb_io_in_ar_valid_REG <= _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_data_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= fb_io_in_r_bits_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_in_fb_r_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  fb_io_in_ar_valid_REG = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  data_r = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Flash(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _rdata_T = 11'h0 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 11'h1 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 11'h2 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [20:0] _rdata_T_3 = _rdata_T ? 21'h10029b : 21'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_4 = _rdata_T_1 ? 25'h1f29293 : 25'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [17:0] _rdata_T_5 = _rdata_T_2 ? 18'h28067 : 18'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_9 = {{4'd0}, _rdata_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_6 = _GEN_9 | _rdata_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_10 = {{7'd0}, _rdata_T_5}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_7 = _rdata_T_6 | _GEN_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = {{39'd0}, _rdata_T_7}; // @[src/main/scala/device/AXI4Flash.scala 37:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4Flash.scala 41:43]
    if (ren_REG) begin // @[src/main/scala/device/AXI4Flash.scala 41:30]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4DummySD(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  sdHelper_clk; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_ren; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_data; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_setAddr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_addr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] regs_0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_1; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_4; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_5; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_6; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_7; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_8; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_15; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_20; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [3:0] strb = io_in_aw_bits_addr[2] ? io_in_w_bits_strb[7:4] : io_in_w_bits_strb[3:0]; // @[src/main/scala/device/AXI4DummySD.scala 138:22]
  wire [7:0] _T_8 = strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_9 = strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_10 = strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_11 = strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [31:0] _T_12 = {_T_11,_T_10,_T_9,_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T = 13'h0 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 13'h38 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 13'h18 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 13'h34 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 13'h14 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_5 = 13'h1c == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_6 = 13'h50 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_7 = 13'h10 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_8 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_9 = 13'h20 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_10 = 13'h40 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_11 = _rdata_T ? regs_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_1 ? regs_15 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_13 = _rdata_T_2 ? regs_6 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdata_T_14 = _rdata_T_3 ? 8'h80 : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_15 = _rdata_T_4 ? regs_5 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_16 = _rdata_T_5 ? regs_7 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_17 = _rdata_T_6 ? regs_20 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_18 = _rdata_T_7 ? regs_4 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_19 = _rdata_T_8 ? regs_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_20 = _rdata_T_9 ? regs_8 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_21 = _rdata_T_10 ? sdHelper_data : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_22 = _rdata_T_11 | _rdata_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_23 = _rdata_T_22 | _rdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_40 = {{24'd0}, _rdata_T_14}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_24 = _rdata_T_23 | _GEN_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_25 = _rdata_T_24 | _rdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_26 = _rdata_T_25 | _rdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_27 = _rdata_T_26 | _rdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_28 = _rdata_T_27 | _rdata_T_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_29 = _rdata_T_28 | _rdata_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_30 = _rdata_T_29 | _rdata_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_31 = _rdata_T_30 | _rdata_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _regs_0_T = io_in_w_bits_data[31:0] & _T_12; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _regs_0_T_1 = ~_T_12; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _regs_0_T_2 = regs_0 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_0_T_3 = _regs_0_T | _regs_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [5:0] regs_0_cmd = _regs_0_T_3[5:0]; // @[src/main/scala/device/AXI4DummySD.scala 84:20]
  wire [31:0] _GEN_9 = 6'hd == regs_0_cmd ? 32'h0 : regs_4; // @[src/main/scala/device/AXI4DummySD.scala 85:18 102:22 72:43]
  wire [31:0] _GEN_10 = 6'hd == regs_0_cmd ? 32'h0 : regs_5; // @[src/main/scala/device/AXI4DummySD.scala 85:18 103:22 72:43]
  wire [31:0] _GEN_11 = 6'hd == regs_0_cmd ? 32'h0 : regs_6; // @[src/main/scala/device/AXI4DummySD.scala 85:18 104:22 72:43]
  wire [31:0] _GEN_12 = 6'hd == regs_0_cmd ? 32'h0 : regs_7; // @[src/main/scala/device/AXI4DummySD.scala 85:18 105:22 72:43]
  wire  _GEN_13 = 6'hd == regs_0_cmd ? 1'h0 : 6'h12 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire [31:0] _GEN_14 = 6'h9 == regs_0_cmd ? 32'h92404001 : _GEN_9; // @[src/main/scala/device/AXI4DummySD.scala 85:18 96:22]
  wire [31:0] _GEN_15 = 6'h9 == regs_0_cmd ? 32'hd24b97e3 : _GEN_10; // @[src/main/scala/device/AXI4DummySD.scala 85:18 97:22]
  wire [31:0] _GEN_16 = 6'h9 == regs_0_cmd ? 32'hf5f803f : _GEN_11; // @[src/main/scala/device/AXI4DummySD.scala 85:18 98:22]
  wire [31:0] _GEN_17 = 6'h9 == regs_0_cmd ? 32'h8c26012a : _GEN_12; // @[src/main/scala/device/AXI4DummySD.scala 85:18 99:22]
  wire  _GEN_18 = 6'h9 == regs_0_cmd ? 1'h0 : _GEN_13; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_23 = 6'h2 == regs_0_cmd ? 1'h0 : _GEN_18; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_28 = 6'h1 == regs_0_cmd ? 1'h0 : _GEN_23; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire [31:0] _regs_15_T_2 = regs_15 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_15_T_3 = _regs_0_T | _regs_15_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_20_T_2 = regs_20 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_20_T_3 = _regs_0_T | _regs_20_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_1_T_2 = regs_1 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_1_T_3 = _regs_0_T | _regs_1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_8_T_2 = regs_8 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_8_T_3 = _regs_0_T | _regs_8_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] rdata = {{32'd0}, _rdata_T_31}; // @[src/main/scala/device/AXI4DummySD.scala 139:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
  SDHelper sdHelper ( // @[src/main/scala/device/AXI4DummySD.scala 114:24]
    .clk(sdHelper_clk),
    .ren(sdHelper_ren),
    .data(sdHelper_data),
    .setAddr(sdHelper_setAddr),
    .addr(sdHelper_addr)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 143:18]
  assign sdHelper_clk = clock; // @[src/main/scala/device/AXI4DummySD.scala 115:19]
  assign sdHelper_ren = io_in_ar_bits_addr[12:0] == 13'h40 & _r_busy_T; // @[src/main/scala/device/AXI4DummySD.scala 116:51]
  assign sdHelper_setAddr = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0 & _GEN_28; // @[src/main/scala/utils/RegMap.scala 32:48 src/main/scala/device/AXI4DummySD.scala 81:25]
  assign sdHelper_addr = regs_1; // @[src/main/scala/device/AXI4DummySD.scala 118:20]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_0 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_0 <= _regs_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_1 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_1 <= _regs_1_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_4 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (6'h1 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h80ff8000; // @[src/main/scala/device/AXI4DummySD.scala 87:22]
      end else if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h1; // @[src/main/scala/device/AXI4DummySD.scala 90:22]
      end else begin
        regs_4 <= _GEN_14;
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 91:22]
        end else begin
          regs_5 <= _GEN_15;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 92:22]
        end else begin
          regs_6 <= _GEN_16;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_7 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_7 <= 32'h15000000; // @[src/main/scala/device/AXI4DummySD.scala 93:22]
        end else begin
          regs_7 <= _GEN_17;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_8 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h20) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_8 <= _regs_8_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_15 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h38) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_15 <= _regs_15_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_20 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h50) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_20 <= _regs_20_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4DummySD.scala 144:49]
    if (ren_REG) begin // @[src/main/scala/device/AXI4DummySD.scala 144:36]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regs_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_4 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_5 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_6 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_7 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_8 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_15 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_20 = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_15[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_rw_req_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_req_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [31:0] io_rw_req_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [3:0]  io_rw_req_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_rw_req_bits_wmask, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [63:0] io_rw_req_bits_wdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_resp_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_rw_resp_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [3:0]  io_rw_resp_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [63:0] io_rw_resp_bits_rdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_out_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_uart_out_ch, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_in_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_uart_in_ch // @[src/main/scala/sim/SimMMIO.scala 28:14]
);
  wire  xbar_clock; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_reset; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_in_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_in_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_0_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_0_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_0_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_1_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_1_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_1_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_2_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_2_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_2_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_3_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_3_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_3_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_4_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_4_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_4_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  uart_clock; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_reset; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_in_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  vga_clock; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_reset; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_fb_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_fb_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [7:0] vga_io_in_fb_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_ctrl_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_vga_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  flash_clock; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_reset; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [31:0] flash_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [63:0] flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  sd_clock; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_reset; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [7:0] sd_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  uart_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] uart_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_fb_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_ctrl_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_ctrl_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_ctrl_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] flash_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] flash_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] flash_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] sd_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  SimpleBusCrossbar1toN_1 xbar ( // @[src/main/scala/sim/SimMMIO.scala 45:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_req_ready(xbar_io_in_req_ready),
    .io_in_req_valid(xbar_io_in_req_valid),
    .io_in_req_bits_addr(xbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(xbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(xbar_io_in_req_bits_wdata),
    .io_in_resp_ready(xbar_io_in_resp_ready),
    .io_in_resp_valid(xbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(xbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(xbar_io_out_0_req_ready),
    .io_out_0_req_valid(xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(xbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(xbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(xbar_io_out_1_req_ready),
    .io_out_1_req_valid(xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(xbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(xbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(xbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(xbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(xbar_io_out_2_req_ready),
    .io_out_2_req_valid(xbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(xbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(xbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(xbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(xbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(xbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(xbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(xbar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(xbar_io_out_3_req_ready),
    .io_out_3_req_valid(xbar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(xbar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_cmd(xbar_io_out_3_req_bits_cmd),
    .io_out_3_req_bits_wmask(xbar_io_out_3_req_bits_wmask),
    .io_out_3_req_bits_wdata(xbar_io_out_3_req_bits_wdata),
    .io_out_3_resp_ready(xbar_io_out_3_resp_ready),
    .io_out_3_resp_valid(xbar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(xbar_io_out_3_resp_bits_rdata),
    .io_out_4_req_ready(xbar_io_out_4_req_ready),
    .io_out_4_req_valid(xbar_io_out_4_req_valid),
    .io_out_4_req_bits_addr(xbar_io_out_4_req_bits_addr),
    .io_out_4_req_bits_cmd(xbar_io_out_4_req_bits_cmd),
    .io_out_4_req_bits_wmask(xbar_io_out_4_req_bits_wmask),
    .io_out_4_req_bits_wdata(xbar_io_out_4_req_bits_wdata),
    .io_out_4_resp_ready(xbar_io_out_4_resp_ready),
    .io_out_4_resp_valid(xbar_io_out_4_resp_valid),
    .io_out_4_resp_bits_rdata(xbar_io_out_4_resp_bits_rdata)
  );
  AXI4UART uart ( // @[src/main/scala/sim/SimMMIO.scala 48:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in_aw_ready(uart_io_in_aw_ready),
    .io_in_aw_valid(uart_io_in_aw_valid),
    .io_in_aw_bits_addr(uart_io_in_aw_bits_addr),
    .io_in_w_ready(uart_io_in_w_ready),
    .io_in_w_valid(uart_io_in_w_valid),
    .io_in_w_bits_data(uart_io_in_w_bits_data),
    .io_in_w_bits_strb(uart_io_in_w_bits_strb),
    .io_in_b_ready(uart_io_in_b_ready),
    .io_in_b_valid(uart_io_in_b_valid),
    .io_in_ar_ready(uart_io_in_ar_ready),
    .io_in_ar_valid(uart_io_in_ar_valid),
    .io_in_ar_bits_addr(uart_io_in_ar_bits_addr),
    .io_in_r_ready(uart_io_in_r_ready),
    .io_in_r_valid(uart_io_in_r_valid),
    .io_in_r_bits_data(uart_io_in_r_bits_data),
    .io_extra_out_valid(uart_io_extra_out_valid),
    .io_extra_out_ch(uart_io_extra_out_ch),
    .io_extra_in_valid(uart_io_extra_in_valid),
    .io_extra_in_ch(uart_io_extra_in_ch)
  );
  AXI4VGA vga ( // @[src/main/scala/sim/SimMMIO.scala 49:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_aw_ready(vga_io_in_fb_aw_ready),
    .io_in_fb_aw_valid(vga_io_in_fb_aw_valid),
    .io_in_fb_aw_bits_addr(vga_io_in_fb_aw_bits_addr),
    .io_in_fb_w_ready(vga_io_in_fb_w_ready),
    .io_in_fb_w_valid(vga_io_in_fb_w_valid),
    .io_in_fb_w_bits_data(vga_io_in_fb_w_bits_data),
    .io_in_fb_w_bits_strb(vga_io_in_fb_w_bits_strb),
    .io_in_fb_b_ready(vga_io_in_fb_b_ready),
    .io_in_fb_b_valid(vga_io_in_fb_b_valid),
    .io_in_fb_ar_ready(vga_io_in_fb_ar_ready),
    .io_in_fb_ar_valid(vga_io_in_fb_ar_valid),
    .io_in_fb_r_ready(vga_io_in_fb_r_ready),
    .io_in_fb_r_valid(vga_io_in_fb_r_valid),
    .io_in_ctrl_aw_ready(vga_io_in_ctrl_aw_ready),
    .io_in_ctrl_aw_valid(vga_io_in_ctrl_aw_valid),
    .io_in_ctrl_w_ready(vga_io_in_ctrl_w_ready),
    .io_in_ctrl_w_valid(vga_io_in_ctrl_w_valid),
    .io_in_ctrl_b_ready(vga_io_in_ctrl_b_ready),
    .io_in_ctrl_b_valid(vga_io_in_ctrl_b_valid),
    .io_in_ctrl_ar_ready(vga_io_in_ctrl_ar_ready),
    .io_in_ctrl_ar_valid(vga_io_in_ctrl_ar_valid),
    .io_in_ctrl_ar_bits_addr(vga_io_in_ctrl_ar_bits_addr),
    .io_in_ctrl_r_ready(vga_io_in_ctrl_r_ready),
    .io_in_ctrl_r_valid(vga_io_in_ctrl_r_valid),
    .io_in_ctrl_r_bits_data(vga_io_in_ctrl_r_bits_data),
    .io_vga_valid(vga_io_vga_valid)
  );
  AXI4Flash flash ( // @[src/main/scala/sim/SimMMIO.scala 50:21]
    .clock(flash_clock),
    .reset(flash_reset),
    .io_in_aw_ready(flash_io_in_aw_ready),
    .io_in_aw_valid(flash_io_in_aw_valid),
    .io_in_w_ready(flash_io_in_w_ready),
    .io_in_w_valid(flash_io_in_w_valid),
    .io_in_b_ready(flash_io_in_b_ready),
    .io_in_b_valid(flash_io_in_b_valid),
    .io_in_ar_ready(flash_io_in_ar_ready),
    .io_in_ar_valid(flash_io_in_ar_valid),
    .io_in_ar_bits_addr(flash_io_in_ar_bits_addr),
    .io_in_r_ready(flash_io_in_r_ready),
    .io_in_r_valid(flash_io_in_r_valid),
    .io_in_r_bits_data(flash_io_in_r_bits_data)
  );
  AXI4DummySD sd ( // @[src/main/scala/sim/SimMMIO.scala 51:18]
    .clock(sd_clock),
    .reset(sd_reset),
    .io_in_aw_ready(sd_io_in_aw_ready),
    .io_in_aw_valid(sd_io_in_aw_valid),
    .io_in_aw_bits_addr(sd_io_in_aw_bits_addr),
    .io_in_w_ready(sd_io_in_w_ready),
    .io_in_w_valid(sd_io_in_w_valid),
    .io_in_w_bits_data(sd_io_in_w_bits_data),
    .io_in_w_bits_strb(sd_io_in_w_bits_strb),
    .io_in_b_ready(sd_io_in_b_ready),
    .io_in_b_valid(sd_io_in_b_valid),
    .io_in_ar_ready(sd_io_in_ar_ready),
    .io_in_ar_valid(sd_io_in_ar_valid),
    .io_in_ar_bits_addr(sd_io_in_ar_bits_addr),
    .io_in_r_ready(sd_io_in_r_ready),
    .io_in_r_valid(sd_io_in_r_valid),
    .io_in_r_bits_data(sd_io_in_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 uart_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(uart_io_in_bridge_clock),
    .reset(uart_io_in_bridge_reset),
    .io_in_req_ready(uart_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(uart_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(uart_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(uart_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(uart_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(uart_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(uart_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(uart_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(uart_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(uart_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(uart_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(uart_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(uart_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(uart_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(uart_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(uart_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(uart_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(uart_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(uart_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(uart_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(uart_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(uart_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(uart_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(uart_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 vga_io_in_fb_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_fb_bridge_clock),
    .reset(vga_io_in_fb_bridge_reset),
    .io_in_req_ready(vga_io_in_fb_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_fb_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_fb_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_fb_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(vga_io_in_fb_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(vga_io_in_fb_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(vga_io_in_fb_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_fb_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(vga_io_in_fb_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(vga_io_in_fb_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_fb_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(vga_io_in_fb_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(vga_io_in_fb_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_fb_bridge_io_out_w_valid),
    .io_out_w_bits_data(vga_io_in_fb_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(vga_io_in_fb_bridge_io_out_w_bits_strb),
    .io_out_b_ready(vga_io_in_fb_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_fb_bridge_io_out_b_valid),
    .io_out_ar_ready(vga_io_in_fb_bridge_io_out_ar_ready),
    .io_out_ar_valid(vga_io_in_fb_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_fb_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_fb_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_fb_bridge_io_out_r_valid),
    .io_out_r_bits_data(vga_io_in_fb_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 vga_io_in_ctrl_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_ctrl_bridge_clock),
    .reset(vga_io_in_ctrl_bridge_reset),
    .io_in_req_ready(vga_io_in_ctrl_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_ctrl_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_ctrl_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_ctrl_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(vga_io_in_ctrl_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(vga_io_in_ctrl_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(vga_io_in_ctrl_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_ctrl_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(vga_io_in_ctrl_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(vga_io_in_ctrl_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_ctrl_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(vga_io_in_ctrl_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(vga_io_in_ctrl_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_ctrl_bridge_io_out_w_valid),
    .io_out_w_bits_data(vga_io_in_ctrl_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(vga_io_in_ctrl_bridge_io_out_w_bits_strb),
    .io_out_b_ready(vga_io_in_ctrl_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_ctrl_bridge_io_out_b_valid),
    .io_out_ar_ready(vga_io_in_ctrl_bridge_io_out_ar_ready),
    .io_out_ar_valid(vga_io_in_ctrl_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_ctrl_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_ctrl_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_ctrl_bridge_io_out_r_valid),
    .io_out_r_bits_data(vga_io_in_ctrl_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 flash_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(flash_io_in_bridge_clock),
    .reset(flash_io_in_bridge_reset),
    .io_in_req_ready(flash_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(flash_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(flash_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(flash_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(flash_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(flash_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(flash_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(flash_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(flash_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(flash_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(flash_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(flash_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(flash_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(flash_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(flash_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(flash_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(flash_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(flash_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(flash_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(flash_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(flash_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(flash_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(flash_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(flash_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 sd_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(sd_io_in_bridge_clock),
    .reset(sd_io_in_bridge_reset),
    .io_in_req_ready(sd_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(sd_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(sd_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(sd_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(sd_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(sd_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(sd_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(sd_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(sd_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(sd_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(sd_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(sd_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(sd_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(sd_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(sd_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(sd_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(sd_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(sd_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(sd_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(sd_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(sd_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(sd_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(sd_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(sd_io_in_bridge_io_out_r_bits_data)
  );
  assign io_rw_req_ready = xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_valid = xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_cmd = xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_rdata = xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_uart_out_valid = uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_out_ch = uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_in_valid = uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_req_valid = io_rw_req_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_addr = io_rw_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_cmd = io_rw_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wmask = io_rw_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wdata = io_rw_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_resp_ready = io_rw_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_out_0_req_ready = uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_valid = uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_bits_rdata = uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_req_ready = vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_valid = vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_bits_rdata = vga_io_in_fb_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_req_ready = vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_valid = vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_bits_rdata = vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_req_ready = flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_valid = flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_bits_rdata = flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_req_ready = sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_valid = sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_bits_rdata = sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in_aw_valid = uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_aw_bits_addr = uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_valid = uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_data = uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_strb = uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_b_ready = uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_valid = uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_bits_addr = uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_r_ready = uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_extra_in_ch = io_uart_in_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_aw_valid = vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_aw_bits_addr = vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_valid = vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_data = vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_strb = vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_b_ready = vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_ar_valid = vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_r_ready = vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_aw_valid = vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_w_valid = vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_b_ready = vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_valid = vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_bits_addr = vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_r_ready = vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_clock = clock;
  assign flash_reset = reset;
  assign flash_io_in_aw_valid = flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_w_valid = flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_b_ready = flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_valid = flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_bits_addr = flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_r_ready = flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_clock = clock;
  assign sd_reset = reset;
  assign sd_io_in_aw_valid = sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_aw_bits_addr = sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_valid = sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_data = sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_strb = sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_b_ready = sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_valid = sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_bits_addr = sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_r_ready = sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign uart_io_in_bridge_clock = clock;
  assign uart_io_in_bridge_reset = reset;
  assign uart_io_in_bridge_io_in_req_valid = xbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_addr = xbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_resp_ready = xbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_out_aw_ready = uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_w_ready = uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_b_valid = uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_ar_ready = uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_valid = uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_bits_data = uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign vga_io_in_fb_bridge_clock = clock;
  assign vga_io_in_fb_bridge_reset = reset;
  assign vga_io_in_fb_bridge_io_in_req_valid = xbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_addr = xbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_cmd = xbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wmask = xbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wdata = xbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_resp_ready = xbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_out_aw_ready = vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_w_ready = vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_b_valid = vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_ar_ready = 1'h1; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_r_valid = vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_r_bits_data = 64'h0; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_bridge_clock = clock;
  assign vga_io_in_ctrl_bridge_reset = reset;
  assign vga_io_in_ctrl_bridge_io_in_req_valid = xbar_io_out_2_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_addr = xbar_io_out_2_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_cmd = xbar_io_out_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_wmask = xbar_io_out_2_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_wdata = xbar_io_out_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_resp_ready = xbar_io_out_2_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_out_aw_ready = vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_w_ready = vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_b_valid = vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_ar_ready = vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_valid = vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_bits_data = vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_io_in_bridge_clock = clock;
  assign flash_io_in_bridge_reset = reset;
  assign flash_io_in_bridge_io_in_req_valid = xbar_io_out_3_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_addr = xbar_io_out_3_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_3_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_3_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_resp_ready = xbar_io_out_3_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_out_aw_ready = flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_w_ready = flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_b_valid = flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_ar_ready = flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_valid = flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_bits_data = flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_io_in_bridge_clock = clock;
  assign sd_io_in_bridge_reset = reset;
  assign sd_io_in_bridge_io_in_req_valid = xbar_io_out_4_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_addr = xbar_io_out_4_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_4_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_4_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_4_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_resp_ready = xbar_io_out_4_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_out_aw_ready = sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_w_ready = sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_b_valid = sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_ar_ready = sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_valid = sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_bits_data = sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
endmodule
module SimTop(
  input         clock,
  input         reset,
  output [63:0] difftest_exit, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [63:0] difftest_step, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_clean, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_dump, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_begin, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_end, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_level, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_out_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [7:0]  difftest_uart_out_ch, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_in_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [7:0]  difftest_uart_in_ch // @[difftest/src/main/scala/Difftest.scala 496:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  soc_clock; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_reset; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [2:0] soc_io_mem_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [1:0] soc_io_mem_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_b_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [2:0] soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  mem_clock; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_reset; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [2:0] mem_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [1:0] mem_io_in_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_in_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [1:0] memdelay_io_in_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [1:0] memdelay_io_out_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  mmio_clock; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_reset; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [31:0] mmio_io_rw_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_rw_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  reg [63:0] difftest_timer; // @[difftest/src/main/scala/Difftest.scala 501:24]
  wire [63:0] _difftest_timer_T_1 = difftest_timer + 64'h1; // @[difftest/src/main/scala/Difftest.scala 502:20]
  wire  difftest_log_enable = difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end; // @[difftest/src/main/scala/Difftest.scala 650:26]
  NutShell soc ( // @[src/main/scala/sim/NutShellSim.scala 34:19]
    .clock(soc_clock),
    .reset(soc_reset),
    .io_mem_aw_ready(soc_io_mem_aw_ready),
    .io_mem_aw_valid(soc_io_mem_aw_valid),
    .io_mem_aw_bits_addr(soc_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(soc_io_mem_aw_bits_len),
    .io_mem_aw_bits_size(soc_io_mem_aw_bits_size),
    .io_mem_aw_bits_burst(soc_io_mem_aw_bits_burst),
    .io_mem_w_ready(soc_io_mem_w_ready),
    .io_mem_w_valid(soc_io_mem_w_valid),
    .io_mem_w_bits_data(soc_io_mem_w_bits_data),
    .io_mem_w_bits_strb(soc_io_mem_w_bits_strb),
    .io_mem_w_bits_last(soc_io_mem_w_bits_last),
    .io_mem_b_valid(soc_io_mem_b_valid),
    .io_mem_ar_ready(soc_io_mem_ar_ready),
    .io_mem_ar_valid(soc_io_mem_ar_valid),
    .io_mem_ar_bits_addr(soc_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(soc_io_mem_ar_bits_len),
    .io_mem_ar_bits_size(soc_io_mem_ar_bits_size),
    .io_mem_r_valid(soc_io_mem_r_valid),
    .io_mem_r_bits_data(soc_io_mem_r_bits_data),
    .io_mem_r_bits_last(soc_io_mem_r_bits_last),
    .io_mmio_req_ready(soc_io_mmio_req_ready),
    .io_mmio_req_valid(soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr(soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(soc_io_mmio_resp_ready),
    .io_mmio_resp_valid(soc_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(soc_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(soc_io_mmio_resp_bits_rdata)
  );
  AXI4RAM mem ( // @[src/main/scala/sim/NutShellSim.scala 35:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_aw_ready(mem_io_in_aw_ready),
    .io_in_aw_valid(mem_io_in_aw_valid),
    .io_in_aw_bits_addr(mem_io_in_aw_bits_addr),
    .io_in_w_ready(mem_io_in_w_ready),
    .io_in_w_valid(mem_io_in_w_valid),
    .io_in_w_bits_data(mem_io_in_w_bits_data),
    .io_in_w_bits_strb(mem_io_in_w_bits_strb),
    .io_in_w_bits_last(mem_io_in_w_bits_last),
    .io_in_b_valid(mem_io_in_b_valid),
    .io_in_ar_ready(mem_io_in_ar_ready),
    .io_in_ar_valid(mem_io_in_ar_valid),
    .io_in_ar_bits_addr(mem_io_in_ar_bits_addr),
    .io_in_ar_bits_len(mem_io_in_ar_bits_len),
    .io_in_ar_bits_size(mem_io_in_ar_bits_size),
    .io_in_ar_bits_burst(mem_io_in_ar_bits_burst),
    .io_in_r_valid(mem_io_in_r_valid),
    .io_in_r_bits_data(mem_io_in_r_bits_data),
    .io_in_r_bits_last(mem_io_in_r_bits_last)
  );
  AXI4Delayer memdelay ( // @[src/main/scala/sim/NutShellSim.scala 38:24]
    .io_in_aw_ready(memdelay_io_in_aw_ready),
    .io_in_aw_valid(memdelay_io_in_aw_valid),
    .io_in_aw_bits_addr(memdelay_io_in_aw_bits_addr),
    .io_in_aw_bits_len(memdelay_io_in_aw_bits_len),
    .io_in_aw_bits_size(memdelay_io_in_aw_bits_size),
    .io_in_aw_bits_burst(memdelay_io_in_aw_bits_burst),
    .io_in_w_ready(memdelay_io_in_w_ready),
    .io_in_w_valid(memdelay_io_in_w_valid),
    .io_in_w_bits_data(memdelay_io_in_w_bits_data),
    .io_in_w_bits_strb(memdelay_io_in_w_bits_strb),
    .io_in_w_bits_last(memdelay_io_in_w_bits_last),
    .io_in_b_valid(memdelay_io_in_b_valid),
    .io_in_ar_ready(memdelay_io_in_ar_ready),
    .io_in_ar_valid(memdelay_io_in_ar_valid),
    .io_in_ar_bits_addr(memdelay_io_in_ar_bits_addr),
    .io_in_ar_bits_len(memdelay_io_in_ar_bits_len),
    .io_in_ar_bits_size(memdelay_io_in_ar_bits_size),
    .io_in_r_valid(memdelay_io_in_r_valid),
    .io_in_r_bits_data(memdelay_io_in_r_bits_data),
    .io_in_r_bits_last(memdelay_io_in_r_bits_last),
    .io_out_aw_ready(memdelay_io_out_aw_ready),
    .io_out_aw_valid(memdelay_io_out_aw_valid),
    .io_out_aw_bits_addr(memdelay_io_out_aw_bits_addr),
    .io_out_w_ready(memdelay_io_out_w_ready),
    .io_out_w_valid(memdelay_io_out_w_valid),
    .io_out_w_bits_data(memdelay_io_out_w_bits_data),
    .io_out_w_bits_strb(memdelay_io_out_w_bits_strb),
    .io_out_w_bits_last(memdelay_io_out_w_bits_last),
    .io_out_b_valid(memdelay_io_out_b_valid),
    .io_out_ar_valid(memdelay_io_out_ar_valid),
    .io_out_ar_bits_addr(memdelay_io_out_ar_bits_addr),
    .io_out_ar_bits_len(memdelay_io_out_ar_bits_len),
    .io_out_ar_bits_size(memdelay_io_out_ar_bits_size),
    .io_out_ar_bits_burst(memdelay_io_out_ar_bits_burst),
    .io_out_r_valid(memdelay_io_out_r_valid),
    .io_out_r_bits_data(memdelay_io_out_r_bits_data),
    .io_out_r_bits_last(memdelay_io_out_r_bits_last)
  );
  SimMMIO mmio ( // @[src/main/scala/sim/NutShellSim.scala 39:20]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_rw_req_ready(mmio_io_rw_req_ready),
    .io_rw_req_valid(mmio_io_rw_req_valid),
    .io_rw_req_bits_addr(mmio_io_rw_req_bits_addr),
    .io_rw_req_bits_cmd(mmio_io_rw_req_bits_cmd),
    .io_rw_req_bits_wmask(mmio_io_rw_req_bits_wmask),
    .io_rw_req_bits_wdata(mmio_io_rw_req_bits_wdata),
    .io_rw_resp_ready(mmio_io_rw_resp_ready),
    .io_rw_resp_valid(mmio_io_rw_resp_valid),
    .io_rw_resp_bits_cmd(mmio_io_rw_resp_bits_cmd),
    .io_rw_resp_bits_rdata(mmio_io_rw_resp_bits_rdata),
    .io_uart_out_valid(mmio_io_uart_out_valid),
    .io_uart_out_ch(mmio_io_uart_out_ch),
    .io_uart_in_valid(mmio_io_uart_in_valid),
    .io_uart_in_ch(mmio_io_uart_in_ch)
  );
  assign difftest_exit = 64'h0; // @[difftest/src/main/scala/Difftest.scala 498:19]
  assign difftest_step = 64'h1; // @[difftest/src/main/scala/Difftest.scala 499:19]
  assign difftest_uart_out_valid = mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_out_ch = mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_in_valid = mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign soc_clock = clock;
  assign soc_reset = reset;
  assign soc_io_mem_aw_ready = memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_w_ready = memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_b_valid = memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_ar_ready = memdelay_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_valid = memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_data = memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_last = memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mmio_req_ready = mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_valid = mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_cmd = mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_rdata = mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_aw_valid = memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_aw_bits_addr = memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_valid = memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_data = memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_strb = memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_last = memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_valid = memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_addr = memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_len = memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_size = memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_burst = memdelay_io_out_ar_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_in_aw_valid = soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_addr = soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_len = soc_io_mem_aw_bits_len; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_size = soc_io_mem_aw_bits_size; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_burst = soc_io_mem_aw_bits_burst; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_valid = soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_data = soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_strb = soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_last = soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_valid = soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_addr = soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_len = soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_size = soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_out_aw_ready = mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_w_ready = mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_b_valid = mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_valid = mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_data = mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_last = mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_rw_req_valid = soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_addr = soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_cmd = soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wmask = soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wdata = soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_resp_ready = soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_uart_in_ch = difftest_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/Difftest.scala 501:24]
      difftest_timer <= 64'h0; // @[difftest/src/main/scala/Difftest.scala 501:24]
    end else begin
      difftest_timer <= _difftest_timer_T_1; // @[difftest/src/main/scala/Difftest.scala 502:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(difftest_logCtrl_begin <= difftest_logCtrl_end)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutShellSim.scala:57 assert(log_begin <= log_end)\n"); // @[src/main/scala/sim/NutShellSim.scala 57:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_timer = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(difftest_logCtrl_begin <= difftest_logCtrl_end); // @[src/main/scala/sim/NutShellSim.scala 57:9]
    end
  end
endmodule
module array_0(
  input  [8:0]  R0_addr,
  input         R0_en,
  input         R0_clk,
  output [73:0] R0_data,
  input  [8:0]  W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [73:0] W0_data
);
  wire [8:0] array_0_ext_R0_addr;
  wire  array_0_ext_R0_en;
  wire  array_0_ext_R0_clk;
  wire [73:0] array_0_ext_R0_data;
  wire [8:0] array_0_ext_W0_addr;
  wire  array_0_ext_W0_en;
  wire  array_0_ext_W0_clk;
  wire [73:0] array_0_ext_W0_data;
  array_0_ext array_0_ext (
    .R0_addr(array_0_ext_R0_addr),
    .R0_en(array_0_ext_R0_en),
    .R0_clk(array_0_ext_R0_clk),
    .R0_data(array_0_ext_R0_data),
    .W0_addr(array_0_ext_W0_addr),
    .W0_en(array_0_ext_W0_en),
    .W0_clk(array_0_ext_W0_clk),
    .W0_data(array_0_ext_W0_data)
  );
  assign array_0_ext_R0_clk = R0_clk;
  assign array_0_ext_R0_en = R0_en;
  assign array_0_ext_R0_addr = R0_addr;
  assign R0_data = array_0_ext_R0_data;
  assign array_0_ext_W0_clk = W0_clk;
  assign array_0_ext_W0_en = W0_en;
  assign array_0_ext_W0_addr = W0_addr;
  assign array_0_ext_W0_data = W0_data;
endmodule
