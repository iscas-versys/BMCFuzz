
/*verilator tracing_off*/
module GEN_w129_toggle(
  input clock,
  input reset,
  input [129 - 1: 0] valid
);
  parameter COVER_TOTAL = 11747;
  parameter COVER_INDEX;
`ifndef SYNTHESIS
  import "DPI-C" function void v_cover_toggle (
    longint cover_index
  );
  always @(posedge clock) begin
    if (!reset) begin
            if (valid[0]) begin
        v_cover_toggle(COVER_INDEX + 0);
      end
      if (valid[1]) begin
        v_cover_toggle(COVER_INDEX + 1);
      end
      if (valid[2]) begin
        v_cover_toggle(COVER_INDEX + 2);
      end
      if (valid[3]) begin
        v_cover_toggle(COVER_INDEX + 3);
      end
      if (valid[4]) begin
        v_cover_toggle(COVER_INDEX + 4);
      end
      if (valid[5]) begin
        v_cover_toggle(COVER_INDEX + 5);
      end
      if (valid[6]) begin
        v_cover_toggle(COVER_INDEX + 6);
      end
      if (valid[7]) begin
        v_cover_toggle(COVER_INDEX + 7);
      end
      if (valid[8]) begin
        v_cover_toggle(COVER_INDEX + 8);
      end
      if (valid[9]) begin
        v_cover_toggle(COVER_INDEX + 9);
      end
      if (valid[10]) begin
        v_cover_toggle(COVER_INDEX + 10);
      end
      if (valid[11]) begin
        v_cover_toggle(COVER_INDEX + 11);
      end
      if (valid[12]) begin
        v_cover_toggle(COVER_INDEX + 12);
      end
      if (valid[13]) begin
        v_cover_toggle(COVER_INDEX + 13);
      end
      if (valid[14]) begin
        v_cover_toggle(COVER_INDEX + 14);
      end
      if (valid[15]) begin
        v_cover_toggle(COVER_INDEX + 15);
      end
      if (valid[16]) begin
        v_cover_toggle(COVER_INDEX + 16);
      end
      if (valid[17]) begin
        v_cover_toggle(COVER_INDEX + 17);
      end
      if (valid[18]) begin
        v_cover_toggle(COVER_INDEX + 18);
      end
      if (valid[19]) begin
        v_cover_toggle(COVER_INDEX + 19);
      end
      if (valid[20]) begin
        v_cover_toggle(COVER_INDEX + 20);
      end
      if (valid[21]) begin
        v_cover_toggle(COVER_INDEX + 21);
      end
      if (valid[22]) begin
        v_cover_toggle(COVER_INDEX + 22);
      end
      if (valid[23]) begin
        v_cover_toggle(COVER_INDEX + 23);
      end
      if (valid[24]) begin
        v_cover_toggle(COVER_INDEX + 24);
      end
      if (valid[25]) begin
        v_cover_toggle(COVER_INDEX + 25);
      end
      if (valid[26]) begin
        v_cover_toggle(COVER_INDEX + 26);
      end
      if (valid[27]) begin
        v_cover_toggle(COVER_INDEX + 27);
      end
      if (valid[28]) begin
        v_cover_toggle(COVER_INDEX + 28);
      end
      if (valid[29]) begin
        v_cover_toggle(COVER_INDEX + 29);
      end
      if (valid[30]) begin
        v_cover_toggle(COVER_INDEX + 30);
      end
      if (valid[31]) begin
        v_cover_toggle(COVER_INDEX + 31);
      end
      if (valid[32]) begin
        v_cover_toggle(COVER_INDEX + 32);
      end
      if (valid[33]) begin
        v_cover_toggle(COVER_INDEX + 33);
      end
      if (valid[34]) begin
        v_cover_toggle(COVER_INDEX + 34);
      end
      if (valid[35]) begin
        v_cover_toggle(COVER_INDEX + 35);
      end
      if (valid[36]) begin
        v_cover_toggle(COVER_INDEX + 36);
      end
      if (valid[37]) begin
        v_cover_toggle(COVER_INDEX + 37);
      end
      if (valid[38]) begin
        v_cover_toggle(COVER_INDEX + 38);
      end
      if (valid[39]) begin
        v_cover_toggle(COVER_INDEX + 39);
      end
      if (valid[40]) begin
        v_cover_toggle(COVER_INDEX + 40);
      end
      if (valid[41]) begin
        v_cover_toggle(COVER_INDEX + 41);
      end
      if (valid[42]) begin
        v_cover_toggle(COVER_INDEX + 42);
      end
      if (valid[43]) begin
        v_cover_toggle(COVER_INDEX + 43);
      end
      if (valid[44]) begin
        v_cover_toggle(COVER_INDEX + 44);
      end
      if (valid[45]) begin
        v_cover_toggle(COVER_INDEX + 45);
      end
      if (valid[46]) begin
        v_cover_toggle(COVER_INDEX + 46);
      end
      if (valid[47]) begin
        v_cover_toggle(COVER_INDEX + 47);
      end
      if (valid[48]) begin
        v_cover_toggle(COVER_INDEX + 48);
      end
      if (valid[49]) begin
        v_cover_toggle(COVER_INDEX + 49);
      end
      if (valid[50]) begin
        v_cover_toggle(COVER_INDEX + 50);
      end
      if (valid[51]) begin
        v_cover_toggle(COVER_INDEX + 51);
      end
      if (valid[52]) begin
        v_cover_toggle(COVER_INDEX + 52);
      end
      if (valid[53]) begin
        v_cover_toggle(COVER_INDEX + 53);
      end
      if (valid[54]) begin
        v_cover_toggle(COVER_INDEX + 54);
      end
      if (valid[55]) begin
        v_cover_toggle(COVER_INDEX + 55);
      end
      if (valid[56]) begin
        v_cover_toggle(COVER_INDEX + 56);
      end
      if (valid[57]) begin
        v_cover_toggle(COVER_INDEX + 57);
      end
      if (valid[58]) begin
        v_cover_toggle(COVER_INDEX + 58);
      end
      if (valid[59]) begin
        v_cover_toggle(COVER_INDEX + 59);
      end
      if (valid[60]) begin
        v_cover_toggle(COVER_INDEX + 60);
      end
      if (valid[61]) begin
        v_cover_toggle(COVER_INDEX + 61);
      end
      if (valid[62]) begin
        v_cover_toggle(COVER_INDEX + 62);
      end
      if (valid[63]) begin
        v_cover_toggle(COVER_INDEX + 63);
      end
      if (valid[64]) begin
        v_cover_toggle(COVER_INDEX + 64);
      end
      if (valid[65]) begin
        v_cover_toggle(COVER_INDEX + 65);
      end
      if (valid[66]) begin
        v_cover_toggle(COVER_INDEX + 66);
      end
      if (valid[67]) begin
        v_cover_toggle(COVER_INDEX + 67);
      end
      if (valid[68]) begin
        v_cover_toggle(COVER_INDEX + 68);
      end
      if (valid[69]) begin
        v_cover_toggle(COVER_INDEX + 69);
      end
      if (valid[70]) begin
        v_cover_toggle(COVER_INDEX + 70);
      end
      if (valid[71]) begin
        v_cover_toggle(COVER_INDEX + 71);
      end
      if (valid[72]) begin
        v_cover_toggle(COVER_INDEX + 72);
      end
      if (valid[73]) begin
        v_cover_toggle(COVER_INDEX + 73);
      end
      if (valid[74]) begin
        v_cover_toggle(COVER_INDEX + 74);
      end
      if (valid[75]) begin
        v_cover_toggle(COVER_INDEX + 75);
      end
      if (valid[76]) begin
        v_cover_toggle(COVER_INDEX + 76);
      end
      if (valid[77]) begin
        v_cover_toggle(COVER_INDEX + 77);
      end
      if (valid[78]) begin
        v_cover_toggle(COVER_INDEX + 78);
      end
      if (valid[79]) begin
        v_cover_toggle(COVER_INDEX + 79);
      end
      if (valid[80]) begin
        v_cover_toggle(COVER_INDEX + 80);
      end
      if (valid[81]) begin
        v_cover_toggle(COVER_INDEX + 81);
      end
      if (valid[82]) begin
        v_cover_toggle(COVER_INDEX + 82);
      end
      if (valid[83]) begin
        v_cover_toggle(COVER_INDEX + 83);
      end
      if (valid[84]) begin
        v_cover_toggle(COVER_INDEX + 84);
      end
      if (valid[85]) begin
        v_cover_toggle(COVER_INDEX + 85);
      end
      if (valid[86]) begin
        v_cover_toggle(COVER_INDEX + 86);
      end
      if (valid[87]) begin
        v_cover_toggle(COVER_INDEX + 87);
      end
      if (valid[88]) begin
        v_cover_toggle(COVER_INDEX + 88);
      end
      if (valid[89]) begin
        v_cover_toggle(COVER_INDEX + 89);
      end
      if (valid[90]) begin
        v_cover_toggle(COVER_INDEX + 90);
      end
      if (valid[91]) begin
        v_cover_toggle(COVER_INDEX + 91);
      end
      if (valid[92]) begin
        v_cover_toggle(COVER_INDEX + 92);
      end
      if (valid[93]) begin
        v_cover_toggle(COVER_INDEX + 93);
      end
      if (valid[94]) begin
        v_cover_toggle(COVER_INDEX + 94);
      end
      if (valid[95]) begin
        v_cover_toggle(COVER_INDEX + 95);
      end
      if (valid[96]) begin
        v_cover_toggle(COVER_INDEX + 96);
      end
      if (valid[97]) begin
        v_cover_toggle(COVER_INDEX + 97);
      end
      if (valid[98]) begin
        v_cover_toggle(COVER_INDEX + 98);
      end
      if (valid[99]) begin
        v_cover_toggle(COVER_INDEX + 99);
      end
      if (valid[100]) begin
        v_cover_toggle(COVER_INDEX + 100);
      end
      if (valid[101]) begin
        v_cover_toggle(COVER_INDEX + 101);
      end
      if (valid[102]) begin
        v_cover_toggle(COVER_INDEX + 102);
      end
      if (valid[103]) begin
        v_cover_toggle(COVER_INDEX + 103);
      end
      if (valid[104]) begin
        v_cover_toggle(COVER_INDEX + 104);
      end
      if (valid[105]) begin
        v_cover_toggle(COVER_INDEX + 105);
      end
      if (valid[106]) begin
        v_cover_toggle(COVER_INDEX + 106);
      end
      if (valid[107]) begin
        v_cover_toggle(COVER_INDEX + 107);
      end
      if (valid[108]) begin
        v_cover_toggle(COVER_INDEX + 108);
      end
      if (valid[109]) begin
        v_cover_toggle(COVER_INDEX + 109);
      end
      if (valid[110]) begin
        v_cover_toggle(COVER_INDEX + 110);
      end
      if (valid[111]) begin
        v_cover_toggle(COVER_INDEX + 111);
      end
      if (valid[112]) begin
        v_cover_toggle(COVER_INDEX + 112);
      end
      if (valid[113]) begin
        v_cover_toggle(COVER_INDEX + 113);
      end
      if (valid[114]) begin
        v_cover_toggle(COVER_INDEX + 114);
      end
      if (valid[115]) begin
        v_cover_toggle(COVER_INDEX + 115);
      end
      if (valid[116]) begin
        v_cover_toggle(COVER_INDEX + 116);
      end
      if (valid[117]) begin
        v_cover_toggle(COVER_INDEX + 117);
      end
      if (valid[118]) begin
        v_cover_toggle(COVER_INDEX + 118);
      end
      if (valid[119]) begin
        v_cover_toggle(COVER_INDEX + 119);
      end
      if (valid[120]) begin
        v_cover_toggle(COVER_INDEX + 120);
      end
      if (valid[121]) begin
        v_cover_toggle(COVER_INDEX + 121);
      end
      if (valid[122]) begin
        v_cover_toggle(COVER_INDEX + 122);
      end
      if (valid[123]) begin
        v_cover_toggle(COVER_INDEX + 123);
      end
      if (valid[124]) begin
        v_cover_toggle(COVER_INDEX + 124);
      end
      if (valid[125]) begin
        v_cover_toggle(COVER_INDEX + 125);
      end
      if (valid[126]) begin
        v_cover_toggle(COVER_INDEX + 126);
      end
      if (valid[127]) begin
        v_cover_toggle(COVER_INDEX + 127);
      end
      if (valid[128]) begin
        v_cover_toggle(COVER_INDEX + 128);
      end
    end
  end
`endif
endmodule
